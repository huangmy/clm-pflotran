netcdf ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-12-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-12-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "fractional area burned" ;
		FAREA_BURNED:units = "proportion/sec" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 08/21/14 13:06:43" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:natpft_not_vegetated = 1 ;
		:natpft_needleleaf_evergreen_temperate_tree = 2 ;
		:natpft_needleleaf_evergreen_boreal_tree = 3 ;
		:natpft_needleleaf_deciduous_boreal_tree = 4 ;
		:natpft_broadleaf_evergreen_tropical_tree = 5 ;
		:natpft_broadleaf_evergreen_temperate_tree = 6 ;
		:natpft_broadleaf_deciduous_tropical_tree = 7 ;
		:natpft_broadleaf_deciduous_temperate_tree = 8 ;
		:natpft_broadleaf_deciduous_boreal_tree = 9 ;
		:natpft_broadleaf_evergreen_shrub = 10 ;
		:natpft_broadleaf_deciduous_temperate_shrub = 11 ;
		:natpft_broadleaf_deciduous_boreal_shrub = 12 ;
		:natpft_c3_arctic_grass = 13 ;
		:natpft_c3_non-arctic_grass = 14 ;
		:natpft_c4_grass = 15 ;
		:natpft_c3_crop = 16 ;
		:natpft_c3_irrigated = 17 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-12-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 11202 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "08/21/14" ;

 time_written =
  "13:06:43" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  5.044949e-14, 5.058576e-14, 5.055929e-14, 5.066909e-14, 5.060821e-14, 
    5.068008e-14, 5.047715e-14, 5.059115e-14, 5.051839e-14, 5.046179e-14, 
    5.088186e-14, 5.067399e-14, 5.109757e-14, 5.096525e-14, 5.129742e-14, 
    5.107696e-14, 5.134183e-14, 5.129111e-14, 5.144381e-14, 5.140008e-14, 
    5.159509e-14, 5.146398e-14, 5.169611e-14, 5.156382e-14, 5.158451e-14, 
    5.145965e-14, 5.071589e-14, 5.085598e-14, 5.070758e-14, 5.072757e-14, 
    5.07186e-14, 5.060945e-14, 5.055439e-14, 5.04391e-14, 5.046004e-14, 
    5.054473e-14, 5.073656e-14, 5.06715e-14, 5.083547e-14, 5.083177e-14, 
    5.101405e-14, 5.093189e-14, 5.123788e-14, 5.1151e-14, 5.140191e-14, 
    5.133885e-14, 5.139894e-14, 5.138073e-14, 5.139918e-14, 5.130669e-14, 
    5.134632e-14, 5.126492e-14, 5.094728e-14, 5.10407e-14, 5.076183e-14, 
    5.059379e-14, 5.048214e-14, 5.040283e-14, 5.041405e-14, 5.043541e-14, 
    5.054522e-14, 5.064841e-14, 5.072698e-14, 5.07795e-14, 5.083124e-14, 
    5.09876e-14, 5.107037e-14, 5.125542e-14, 5.122208e-14, 5.127858e-14, 
    5.133258e-14, 5.142314e-14, 5.140825e-14, 5.144812e-14, 5.127711e-14, 
    5.139078e-14, 5.120307e-14, 5.125444e-14, 5.084517e-14, 5.068906e-14, 
    5.062253e-14, 5.056437e-14, 5.042267e-14, 5.052053e-14, 5.048196e-14, 
    5.057374e-14, 5.063201e-14, 5.06032e-14, 5.078094e-14, 5.071186e-14, 
    5.107527e-14, 5.091887e-14, 5.132628e-14, 5.122893e-14, 5.134961e-14, 
    5.128805e-14, 5.13935e-14, 5.12986e-14, 5.146297e-14, 5.149871e-14, 
    5.147428e-14, 5.156814e-14, 5.129333e-14, 5.139893e-14, 5.060239e-14, 
    5.060708e-14, 5.062899e-14, 5.053268e-14, 5.05268e-14, 5.043851e-14, 
    5.051708e-14, 5.055051e-14, 5.06354e-14, 5.068555e-14, 5.073322e-14, 
    5.083796e-14, 5.095482e-14, 5.111807e-14, 5.123524e-14, 5.131371e-14, 
    5.126561e-14, 5.130807e-14, 5.126059e-14, 5.123834e-14, 5.148531e-14, 
    5.134668e-14, 5.155464e-14, 5.154315e-14, 5.144906e-14, 5.154445e-14, 
    5.061038e-14, 5.058334e-14, 5.048937e-14, 5.056292e-14, 5.04289e-14, 
    5.050392e-14, 5.054702e-14, 5.071328e-14, 5.074981e-14, 5.078363e-14, 
    5.085044e-14, 5.09361e-14, 5.108622e-14, 5.121671e-14, 5.133573e-14, 
    5.132702e-14, 5.133008e-14, 5.135664e-14, 5.129082e-14, 5.136744e-14, 
    5.138028e-14, 5.134668e-14, 5.154161e-14, 5.148596e-14, 5.154291e-14, 
    5.150668e-14, 5.059214e-14, 5.063764e-14, 5.061305e-14, 5.065928e-14, 
    5.06267e-14, 5.077144e-14, 5.08148e-14, 5.101754e-14, 5.093441e-14, 
    5.106672e-14, 5.094787e-14, 5.096893e-14, 5.107098e-14, 5.09543e-14, 
    5.120949e-14, 5.103649e-14, 5.135767e-14, 5.118507e-14, 5.136848e-14, 
    5.133521e-14, 5.139029e-14, 5.143959e-14, 5.15016e-14, 5.161589e-14, 
    5.158944e-14, 5.168497e-14, 5.070545e-14, 5.07644e-14, 5.075924e-14, 
    5.082092e-14, 5.086651e-14, 5.09653e-14, 5.112355e-14, 5.106407e-14, 
    5.117327e-14, 5.119517e-14, 5.102928e-14, 5.113113e-14, 5.080386e-14, 
    5.085677e-14, 5.082528e-14, 5.071009e-14, 5.107774e-14, 5.088918e-14, 
    5.123717e-14, 5.11352e-14, 5.143256e-14, 5.128474e-14, 5.157487e-14, 
    5.169861e-14, 5.181506e-14, 5.195085e-14, 5.079659e-14, 5.075655e-14, 
    5.082826e-14, 5.092736e-14, 5.101932e-14, 5.114141e-14, 5.115391e-14, 
    5.117676e-14, 5.123596e-14, 5.12857e-14, 5.118396e-14, 5.129817e-14, 
    5.086898e-14, 5.109411e-14, 5.074138e-14, 5.084767e-14, 5.092153e-14, 
    5.088916e-14, 5.105728e-14, 5.109686e-14, 5.125756e-14, 5.117453e-14, 
    5.166806e-14, 5.144996e-14, 5.205423e-14, 5.188567e-14, 5.074255e-14, 
    5.079646e-14, 5.09839e-14, 5.089475e-14, 5.114957e-14, 5.12122e-14, 
    5.126311e-14, 5.132812e-14, 5.133515e-14, 5.137365e-14, 5.131056e-14, 
    5.137117e-14, 5.114167e-14, 5.124429e-14, 5.096252e-14, 5.103114e-14, 
    5.099959e-14, 5.096494e-14, 5.107183e-14, 5.118556e-14, 5.118803e-14, 
    5.122447e-14, 5.132701e-14, 5.115061e-14, 5.16961e-14, 5.135945e-14, 
    5.085523e-14, 5.095891e-14, 5.097376e-14, 5.093361e-14, 5.120592e-14, 
    5.110732e-14, 5.137272e-14, 5.130106e-14, 5.141846e-14, 5.136013e-14, 
    5.135155e-14, 5.12766e-14, 5.122989e-14, 5.111183e-14, 5.10157e-14, 
    5.093944e-14, 5.095718e-14, 5.104094e-14, 5.119252e-14, 5.133577e-14, 
    5.13044e-14, 5.140955e-14, 5.113111e-14, 5.124792e-14, 5.120278e-14, 
    5.132047e-14, 5.106248e-14, 5.128208e-14, 5.100627e-14, 5.103049e-14, 
    5.110536e-14, 5.125581e-14, 5.128914e-14, 5.132463e-14, 5.130274e-14, 
    5.119638e-14, 5.117896e-14, 5.110355e-14, 5.10827e-14, 5.102522e-14, 
    5.097758e-14, 5.102109e-14, 5.106677e-14, 5.119644e-14, 5.131315e-14, 
    5.144028e-14, 5.147139e-14, 5.161961e-14, 5.149891e-14, 5.169796e-14, 
    5.152867e-14, 5.182161e-14, 5.129486e-14, 5.152377e-14, 5.110878e-14, 
    5.115357e-14, 5.123449e-14, 5.141997e-14, 5.131992e-14, 5.143694e-14, 
    5.117828e-14, 5.104381e-14, 5.100904e-14, 5.094406e-14, 5.101053e-14, 
    5.100512e-14, 5.106868e-14, 5.104827e-14, 5.120074e-14, 5.111886e-14, 
    5.135132e-14, 5.143602e-14, 5.167495e-14, 5.182114e-14, 5.196983e-14, 
    5.203539e-14, 5.205534e-14, 5.206367e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -7.121268e-15, -7.110204e-15, -7.112354e-15, -7.10344e-15, -7.108385e-15, 
    -7.102549e-15, -7.119026e-15, -7.109763e-15, -7.115676e-15, 
    -7.120274e-15, -7.086174e-15, -7.103043e-15, -7.068723e-15, -7.07944e-15, 
    -7.052563e-15, -7.070387e-15, -7.048977e-15, -7.053081e-15, 
    -7.040748e-15, -7.044279e-15, -7.028524e-15, -7.03912e-15, -7.020384e-15, 
    -7.031056e-15, -7.029383e-15, -7.039469e-15, -7.099649e-15, -7.08827e-15, 
    -7.100323e-15, -7.098699e-15, -7.099429e-15, -7.108281e-15, 
    -7.112745e-15, -7.122118e-15, -7.120416e-15, -7.113533e-15, 
    -7.097969e-15, -7.103251e-15, -7.089958e-15, -7.090257e-15, -7.07549e-15, 
    -7.082144e-15, -7.057384e-15, -7.064411e-15, -7.044132e-15, 
    -7.049224e-15, -7.04437e-15, -7.045842e-15, -7.044351e-15, -7.051822e-15, 
    -7.048619e-15, -7.055199e-15, -7.080896e-15, -7.07333e-15, -7.095922e-15, 
    -7.109542e-15, -7.118618e-15, -7.125063e-15, -7.124152e-15, 
    -7.122414e-15, -7.113494e-15, -7.105124e-15, -7.098752e-15, 
    -7.094493e-15, -7.090301e-15, -7.077616e-15, -7.070924e-15, 
    -7.055961e-15, -7.058663e-15, -7.05409e-15, -7.049731e-15, -7.042415e-15, 
    -7.043619e-15, -7.040397e-15, -7.054214e-15, -7.045026e-15, 
    -7.060201e-15, -7.056046e-15, -7.089145e-15, -7.101826e-15, 
    -7.107211e-15, -7.11194e-15, -7.123451e-15, -7.115499e-15, -7.118632e-15, 
    -7.111184e-15, -7.106455e-15, -7.108793e-15, -7.094377e-15, 
    -7.099977e-15, -7.070528e-15, -7.083194e-15, -7.05024e-15, -7.058109e-15, 
    -7.048356e-15, -7.053331e-15, -7.044807e-15, -7.052478e-15, -7.0392e-15, 
    -7.036311e-15, -7.038284e-15, -7.030712e-15, -7.052903e-15, 
    -7.044369e-15, -7.108859e-15, -7.108477e-15, -7.1067e-15, -7.114512e-15, 
    -7.114991e-15, -7.122164e-15, -7.115782e-15, -7.113066e-15, 
    -7.106182e-15, -7.102111e-15, -7.098245e-15, -7.089753e-15, 
    -7.080282e-15, -7.067069e-15, -7.057598e-15, -7.051257e-15, 
    -7.055146e-15, -7.051713e-15, -7.05555e-15, -7.05735e-15, -7.037392e-15, 
    -7.048588e-15, -7.031801e-15, -7.032729e-15, -7.04032e-15, -7.032624e-15, 
    -7.108209e-15, -7.110405e-15, -7.118032e-15, -7.112063e-15, 
    -7.122946e-15, -7.11685e-15, -7.113345e-15, -7.099856e-15, -7.096901e-15, 
    -7.094156e-15, -7.088744e-15, -7.081803e-15, -7.069647e-15, 
    -7.059093e-15, -7.049478e-15, -7.050183e-15, -7.049934e-15, 
    -7.047787e-15, -7.053106e-15, -7.046915e-15, -7.045875e-15, 
    -7.048592e-15, -7.032853e-15, -7.037345e-15, -7.032749e-15, 
    -7.035673e-15, -7.109692e-15, -7.105998e-15, -7.107993e-15, 
    -7.104241e-15, -7.106883e-15, -7.095139e-15, -7.091622e-15, 
    -7.075201e-15, -7.081939e-15, -7.071223e-15, -7.08085e-15, -7.079143e-15, 
    -7.070868e-15, -7.080331e-15, -7.059671e-15, -7.073664e-15, 
    -7.047704e-15, -7.06164e-15, -7.046831e-15, -7.04952e-15, -7.04507e-15, 
    -7.041087e-15, -7.036082e-15, -7.026855e-15, -7.028991e-15, 
    -7.021286e-15, -7.100497e-15, -7.095713e-15, -7.096137e-15, 
    -7.091136e-15, -7.087439e-15, -7.07944e-15, -7.066629e-15, -7.071444e-15, 
    -7.062611e-15, -7.060838e-15, -7.074261e-15, -7.066013e-15, 
    -7.092515e-15, -7.088222e-15, -7.09078e-15, -7.100118e-15, -7.07033e-15, 
    -7.085596e-15, -7.057441e-15, -7.065688e-15, -7.041654e-15, 
    -7.053591e-15, -7.030166e-15, -7.020175e-15, -7.010803e-15, 
    -6.999854e-15, -7.093106e-15, -7.096355e-15, -7.090542e-15, 
    -7.082504e-15, -7.075064e-15, -7.065184e-15, -7.064176e-15, 
    -7.062326e-15, -7.057542e-15, -7.05352e-15, -7.061738e-15, -7.052513e-15, 
    -7.08722e-15, -7.069008e-15, -7.097581e-15, -7.088958e-15, -7.082979e-15, 
    -7.085604e-15, -7.071995e-15, -7.068791e-15, -7.05579e-15, -7.062509e-15, 
    -7.022636e-15, -7.040241e-15, -6.991543e-15, -7.005106e-15, -7.09749e-15, 
    -7.093119e-15, -7.077928e-15, -7.085152e-15, -7.064527e-15, -7.05946e-15, 
    -7.055347e-15, -7.050089e-15, -7.049524e-15, -7.046412e-15, 
    -7.051512e-15, -7.046614e-15, -7.065163e-15, -7.056867e-15, 
    -7.079667e-15, -7.074107e-15, -7.076665e-15, -7.07947e-15, -7.070817e-15, 
    -7.061608e-15, -7.061416e-15, -7.058466e-15, -7.050151e-15, 
    -7.064443e-15, -7.020359e-15, -7.047534e-15, -7.088356e-15, 
    -7.079947e-15, -7.078753e-15, -7.082007e-15, -7.059968e-15, 
    -7.067943e-15, -7.046488e-15, -7.052279e-15, -7.042795e-15, 
    -7.047506e-15, -7.048198e-15, -7.054256e-15, -7.05803e-15, -7.067576e-15, 
    -7.075356e-15, -7.081536e-15, -7.080099e-15, -7.073313e-15, 
    -7.061047e-15, -7.049471e-15, -7.052004e-15, -7.043515e-15, -7.06602e-15, 
    -7.05657e-15, -7.060218e-15, -7.05071e-15, -7.071571e-15, -7.053787e-15, 
    -7.076124e-15, -7.074163e-15, -7.068101e-15, -7.055926e-15, 
    -7.053243e-15, -7.050371e-15, -7.052144e-15, -7.060737e-15, 
    -7.062148e-15, -7.06825e-15, -7.069933e-15, -7.07459e-15, -7.078446e-15, 
    -7.074922e-15, -7.071222e-15, -7.060735e-15, -7.051298e-15, 
    -7.041029e-15, -7.038521e-15, -7.02654e-15, -7.036284e-15, -7.020207e-15, 
    -7.033862e-15, -7.010251e-15, -7.052765e-15, -7.034274e-15, 
    -7.067827e-15, -7.064204e-15, -7.057652e-15, -7.042662e-15, 
    -7.050754e-15, -7.041294e-15, -7.062203e-15, -7.073076e-15, 
    -7.075899e-15, -7.081159e-15, -7.075779e-15, -7.076216e-15, 
    -7.071072e-15, -7.072725e-15, -7.060387e-15, -7.067011e-15, 
    -7.048215e-15, -7.04137e-15, -7.022091e-15, -7.010303e-15, -6.998338e-15, 
    -6.993062e-15, -6.991457e-15, -6.990787e-15 ;

 CH4_SURF_DIFF_UNSAT =
  1.551417e-14, 1.509146e-14, 1.517365e-14, 1.483266e-14, 1.502184e-14, 
    1.479854e-14, 1.54285e-14, 1.507466e-14, 1.530056e-14, 1.547615e-14, 
    1.417076e-14, 1.481746e-14, 1.349908e-14, 1.39116e-14, 1.287525e-14, 
    1.356324e-14, 1.27365e-14, 1.289516e-14, 1.241773e-14, 1.255452e-14, 
    1.19436e-14, 1.235459e-14, 1.162692e-14, 1.204179e-14, 1.197688e-14, 
    1.236814e-14, 1.468737e-14, 1.425126e-14, 1.47132e-14, 1.465102e-14, 
    1.467893e-14, 1.501791e-14, 1.51887e-14, 1.554651e-14, 1.548156e-14, 
    1.521878e-14, 1.462305e-14, 1.482532e-14, 1.431564e-14, 1.432716e-14, 
    1.37596e-14, 1.401551e-14, 1.306143e-14, 1.333265e-14, 1.254881e-14, 
    1.274596e-14, 1.255806e-14, 1.261505e-14, 1.255732e-14, 1.284646e-14, 
    1.272258e-14, 1.297701e-14, 1.396757e-14, 1.367648e-14, 1.454455e-14, 
    1.506631e-14, 1.541297e-14, 1.56589e-14, 1.562414e-14, 1.555785e-14, 
    1.521724e-14, 1.489702e-14, 1.465296e-14, 1.448969e-14, 1.432881e-14, 
    1.384165e-14, 1.358389e-14, 1.300655e-14, 1.31108e-14, 1.293422e-14, 
    1.276558e-14, 1.248234e-14, 1.252897e-14, 1.240416e-14, 1.293891e-14, 
    1.258351e-14, 1.317017e-14, 1.300973e-14, 1.428488e-14, 1.477076e-14, 
    1.49771e-14, 1.515785e-14, 1.55974e-14, 1.529385e-14, 1.541351e-14, 
    1.512886e-14, 1.494796e-14, 1.503744e-14, 1.448522e-14, 1.469991e-14, 
    1.356861e-14, 1.405596e-14, 1.278525e-14, 1.308941e-14, 1.271234e-14, 
    1.290477e-14, 1.257503e-14, 1.28718e-14, 1.235772e-14, 1.224574e-14, 
    1.232226e-14, 1.202837e-14, 1.288824e-14, 1.255804e-14, 1.503994e-14, 
    1.502534e-14, 1.495737e-14, 1.525615e-14, 1.527444e-14, 1.554828e-14, 
    1.530464e-14, 1.520086e-14, 1.493749e-14, 1.478166e-14, 1.463354e-14, 
    1.430784e-14, 1.394402e-14, 1.343525e-14, 1.306969e-14, 1.282459e-14, 
    1.29749e-14, 1.28422e-14, 1.299054e-14, 1.306007e-14, 1.228769e-14, 
    1.272141e-14, 1.207064e-14, 1.210666e-14, 1.240118e-14, 1.210261e-14, 
    1.50151e-14, 1.509908e-14, 1.539058e-14, 1.516246e-14, 1.55781e-14, 
    1.534543e-14, 1.521162e-14, 1.469538e-14, 1.4582e-14, 1.44768e-14, 
    1.426906e-14, 1.400241e-14, 1.353457e-14, 1.312747e-14, 1.275577e-14, 
    1.278301e-14, 1.277342e-14, 1.269036e-14, 1.289608e-14, 1.265658e-14, 
    1.261637e-14, 1.272149e-14, 1.211149e-14, 1.228578e-14, 1.210743e-14, 
    1.222092e-14, 1.507179e-14, 1.493049e-14, 1.500684e-14, 1.486325e-14, 
    1.496439e-14, 1.451458e-14, 1.43797e-14, 1.374857e-14, 1.400765e-14, 
    1.359535e-14, 1.396579e-14, 1.390014e-14, 1.358182e-14, 1.394578e-14, 
    1.314988e-14, 1.368944e-14, 1.268713e-14, 1.322599e-14, 1.265335e-14, 
    1.275738e-14, 1.258516e-14, 1.243088e-14, 1.22368e-14, 1.187859e-14, 
    1.196155e-14, 1.166197e-14, 1.471984e-14, 1.453653e-14, 1.455271e-14, 
    1.436089e-14, 1.421901e-14, 1.391152e-14, 1.341823e-14, 1.360375e-14, 
    1.326319e-14, 1.31948e-14, 1.371221e-14, 1.339451e-14, 1.441387e-14, 
    1.424917e-14, 1.434726e-14, 1.470536e-14, 1.356095e-14, 1.41483e-14, 
    1.306364e-14, 1.338192e-14, 1.245287e-14, 1.291493e-14, 1.200721e-14, 
    1.161893e-14, 1.125358e-14, 1.08263e-14, 1.443652e-14, 1.456108e-14, 
    1.433808e-14, 1.402947e-14, 1.37432e-14, 1.33625e-14, 1.332357e-14, 
    1.325223e-14, 1.306748e-14, 1.29121e-14, 1.322964e-14, 1.287315e-14, 
    1.42109e-14, 1.350998e-14, 1.460814e-14, 1.427745e-14, 1.404768e-14, 
    1.414851e-14, 1.362496e-14, 1.350154e-14, 1.299991e-14, 1.325926e-14, 
    1.171474e-14, 1.239824e-14, 1.050101e-14, 1.103142e-14, 1.460459e-14, 
    1.443697e-14, 1.385347e-14, 1.413112e-14, 1.33371e-14, 1.31416e-14, 
    1.298269e-14, 1.277946e-14, 1.275754e-14, 1.263713e-14, 1.283444e-14, 
    1.264493e-14, 1.336169e-14, 1.304144e-14, 1.392021e-14, 1.370633e-14, 
    1.380474e-14, 1.391265e-14, 1.357958e-14, 1.322463e-14, 1.32171e-14, 
    1.310326e-14, 1.278232e-14, 1.333389e-14, 1.162639e-14, 1.268099e-14, 
    1.425418e-14, 1.393119e-14, 1.388512e-14, 1.401023e-14, 1.31612e-14, 
    1.346886e-14, 1.264007e-14, 1.286412e-14, 1.249702e-14, 1.267944e-14, 
    1.270628e-14, 1.294055e-14, 1.308638e-14, 1.345475e-14, 1.375444e-14, 
    1.399209e-14, 1.393684e-14, 1.367578e-14, 1.320293e-14, 1.275553e-14, 
    1.285354e-14, 1.252492e-14, 1.339468e-14, 1.303001e-14, 1.317094e-14, 
    1.280343e-14, 1.360867e-14, 1.292281e-14, 1.378392e-14, 1.370845e-14, 
    1.347497e-14, 1.300523e-14, 1.290137e-14, 1.279036e-14, 1.285887e-14, 
    1.319094e-14, 1.324536e-14, 1.348066e-14, 1.354559e-14, 1.372488e-14, 
    1.387328e-14, 1.373768e-14, 1.359526e-14, 1.319082e-14, 1.282623e-14, 
    1.242867e-14, 1.233139e-14, 1.186659e-14, 1.224489e-14, 1.16205e-14, 
    1.215124e-14, 1.123245e-14, 1.288314e-14, 1.216696e-14, 1.346436e-14, 
    1.332465e-14, 1.307187e-14, 1.249205e-14, 1.280516e-14, 1.243901e-14, 
    1.324749e-14, 1.366674e-14, 1.377527e-14, 1.397764e-14, 1.377065e-14, 
    1.378748e-14, 1.35894e-14, 1.365306e-14, 1.317739e-14, 1.343291e-14, 
    1.270693e-14, 1.244192e-14, 1.169335e-14, 1.123424e-14, 1.076686e-14, 
    1.056043e-14, 1.04976e-14, 1.047133e-14 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 
    1.93195e-23, 1.931952e-23, 1.931949e-23, 1.93195e-23, 1.931947e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931945e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931945e-23, 
    1.931946e-23, 1.931951e-23, 1.93195e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931951e-23, 1.931952e-23, 1.93195e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.93195e-23, 1.931949e-23, 1.931951e-23, 
    1.931952e-23, 1.931953e-23, 1.931954e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 1.93195e-23, 
    1.931949e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931947e-23, 1.93195e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 
    1.931949e-23, 1.93195e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931947e-23, 1.931946e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931945e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931953e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931946e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931951e-23, 1.931951e-23, 1.931949e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.93195e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931948e-23, 1.931951e-23, 
    1.93195e-23, 1.931951e-23, 1.931951e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 
    1.931944e-23, 1.931943e-23, 1.931942e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.93195e-23, 1.931949e-23, 1.931951e-23, 1.93195e-23, 1.93195e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 
    1.931944e-23, 1.931946e-23, 1.931942e-23, 1.931943e-23, 1.931951e-23, 
    1.931951e-23, 1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931948e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931944e-23, 1.931947e-23, 
    1.93195e-23, 1.93195e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931947e-23, 1.931949e-23, 1.931947e-23, 1.931949e-23, 1.931949e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931946e-23, 1.931946e-23, 1.931945e-23, 1.931946e-23, 1.931944e-23, 
    1.931945e-23, 1.931943e-23, 1.931947e-23, 1.931946e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 
    1.931948e-23, 1.931949e-23, 1.931949e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931946e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975388e-24, 1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 
    1.975386e-24, 1.975388e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975384e-24, 1.975386e-24, 1.975381e-24, 1.975383e-24, 1.975379e-24, 
    1.975382e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975376e-24, 1.975378e-24, 1.975375e-24, 1.975377e-24, 1.975377e-24, 
    1.975378e-24, 1.975385e-24, 1.975384e-24, 1.975385e-24, 1.975385e-24, 
    1.975385e-24, 1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975385e-24, 1.975386e-24, 1.975384e-24, 1.975384e-24, 
    1.975382e-24, 1.975383e-24, 1.97538e-24, 1.975381e-24, 1.975378e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 1.975385e-24, 
    1.975387e-24, 1.975388e-24, 1.975388e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 1.975384e-24, 
    1.975383e-24, 1.975382e-24, 1.97538e-24, 1.97538e-24, 1.97538e-24, 
    1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 1.97538e-24, 
    1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975384e-24, 1.975386e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 
    1.975382e-24, 1.975383e-24, 1.975379e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975377e-24, 
    1.975378e-24, 1.975377e-24, 1.975379e-24, 1.975379e-24, 1.975386e-24, 
    1.975386e-24, 1.975386e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 1.975379e-24, 
    1.97538e-24, 1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975378e-24, 
    1.975379e-24, 1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975385e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975377e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975386e-24, 
    1.975386e-24, 1.975385e-24, 1.975384e-24, 1.975382e-24, 1.975383e-24, 
    1.975382e-24, 1.975383e-24, 1.975383e-24, 1.975382e-24, 1.975383e-24, 
    1.97538e-24, 1.975382e-24, 1.975379e-24, 1.975381e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975377e-24, 1.975376e-24, 
    1.975377e-24, 1.975376e-24, 1.975385e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975384e-24, 1.975383e-24, 1.975381e-24, 1.975382e-24, 
    1.975381e-24, 1.97538e-24, 1.975382e-24, 1.975381e-24, 1.975384e-24, 
    1.975384e-24, 1.975384e-24, 1.975385e-24, 1.975382e-24, 1.975384e-24, 
    1.97538e-24, 1.975381e-24, 1.975378e-24, 1.975379e-24, 1.975377e-24, 
    1.975375e-24, 1.975374e-24, 1.975373e-24, 1.975384e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.975379e-24, 1.975381e-24, 1.975379e-24, 
    1.975384e-24, 1.975381e-24, 1.975385e-24, 1.975384e-24, 1.975383e-24, 
    1.975384e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.975376e-24, 1.975378e-24, 1.975372e-24, 1.975373e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.975381e-24, 1.975375e-24, 1.975379e-24, 
    1.975384e-24, 1.975383e-24, 1.975383e-24, 1.975383e-24, 1.97538e-24, 
    1.975381e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 1.975382e-24, 
    1.975383e-24, 1.975383e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975381e-24, 1.97538e-24, 1.97538e-24, 
    1.975379e-24, 1.975382e-24, 1.97538e-24, 1.975382e-24, 1.975382e-24, 
    1.975381e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.97538e-24, 1.975381e-24, 1.975381e-24, 1.975382e-24, 1.975382e-24, 
    1.975383e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975378e-24, 1.975378e-24, 1.975376e-24, 1.975377e-24, 1.975375e-24, 
    1.975377e-24, 1.975374e-24, 1.975379e-24, 1.975377e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975378e-24, 
    1.975381e-24, 1.975382e-24, 1.975382e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975381e-24, 
    1.975379e-24, 1.975378e-24, 1.975376e-24, 1.975374e-24, 1.975373e-24, 
    1.975372e-24, 1.975372e-24, 1.975372e-24 ;

 CONC_CH4_SAT =
  3.269901e-08, 3.267834e-08, 3.268237e-08, 3.266568e-08, 3.267495e-08, 
    3.266401e-08, 3.269484e-08, 3.26775e-08, 3.268858e-08, 3.269717e-08, 
    3.263326e-08, 3.266494e-08, 3.260057e-08, 3.262072e-08, 3.25702e-08, 
    3.260368e-08, 3.256346e-08, 3.257121e-08, 3.2548e-08, 3.255465e-08, 
    3.252491e-08, 3.254494e-08, 3.250957e-08, 3.252971e-08, 3.252654e-08, 
    3.254559e-08, 3.26586e-08, 3.263719e-08, 3.265986e-08, 3.265681e-08, 
    3.265819e-08, 3.267474e-08, 3.268306e-08, 3.270062e-08, 3.269744e-08, 
    3.268456e-08, 3.265544e-08, 3.266535e-08, 3.264046e-08, 3.264102e-08, 
    3.261331e-08, 3.26258e-08, 3.25793e-08, 3.259252e-08, 3.255438e-08, 
    3.256395e-08, 3.255482e-08, 3.255759e-08, 3.255478e-08, 3.256883e-08, 
    3.256281e-08, 3.257519e-08, 3.262345e-08, 3.260925e-08, 3.265161e-08, 
    3.267705e-08, 3.269407e-08, 3.270611e-08, 3.270441e-08, 3.270115e-08, 
    3.268448e-08, 3.266885e-08, 3.265693e-08, 3.264896e-08, 3.26411e-08, 
    3.261724e-08, 3.260471e-08, 3.257661e-08, 3.258171e-08, 3.257309e-08, 
    3.256491e-08, 3.255113e-08, 3.255341e-08, 3.254733e-08, 3.257334e-08, 
    3.255604e-08, 3.258461e-08, 3.257679e-08, 3.263883e-08, 3.266268e-08, 
    3.267271e-08, 3.268159e-08, 3.27031e-08, 3.268823e-08, 3.269409e-08, 
    3.268019e-08, 3.267134e-08, 3.267572e-08, 3.264874e-08, 3.265922e-08, 
    3.260397e-08, 3.262775e-08, 3.256586e-08, 3.258067e-08, 3.256232e-08, 
    3.257169e-08, 3.255563e-08, 3.257008e-08, 3.254508e-08, 3.253962e-08, 
    3.254334e-08, 3.252908e-08, 3.257088e-08, 3.25548e-08, 3.267584e-08, 
    3.267512e-08, 3.267181e-08, 3.268639e-08, 3.268729e-08, 3.27007e-08, 
    3.268878e-08, 3.268369e-08, 3.267084e-08, 3.266321e-08, 3.265597e-08, 
    3.264006e-08, 3.262229e-08, 3.259748e-08, 3.257971e-08, 3.256779e-08, 
    3.257511e-08, 3.256864e-08, 3.257586e-08, 3.257925e-08, 3.254165e-08, 
    3.256275e-08, 3.253113e-08, 3.253288e-08, 3.254718e-08, 3.253269e-08, 
    3.267462e-08, 3.267874e-08, 3.269298e-08, 3.268183e-08, 3.270216e-08, 
    3.269076e-08, 3.26842e-08, 3.265897e-08, 3.265346e-08, 3.264831e-08, 
    3.263818e-08, 3.262516e-08, 3.260233e-08, 3.258251e-08, 3.256444e-08, 
    3.256577e-08, 3.25653e-08, 3.256125e-08, 3.257126e-08, 3.255961e-08, 
    3.255764e-08, 3.256276e-08, 3.253312e-08, 3.254159e-08, 3.253292e-08, 
    3.253844e-08, 3.26774e-08, 3.267049e-08, 3.267422e-08, 3.26672e-08, 
    3.267213e-08, 3.265013e-08, 3.264353e-08, 3.261274e-08, 3.262541e-08, 
    3.260529e-08, 3.262338e-08, 3.262016e-08, 3.260457e-08, 3.262241e-08, 
    3.258357e-08, 3.260984e-08, 3.256109e-08, 3.258724e-08, 3.255945e-08, 
    3.256452e-08, 3.255614e-08, 3.254863e-08, 3.253921e-08, 3.252179e-08, 
    3.252583e-08, 3.251129e-08, 3.26602e-08, 3.265122e-08, 3.265204e-08, 
    3.264266e-08, 3.263573e-08, 3.262073e-08, 3.259667e-08, 3.260573e-08, 
    3.258913e-08, 3.25858e-08, 3.261102e-08, 3.25955e-08, 3.264523e-08, 
    3.263716e-08, 3.264199e-08, 3.265947e-08, 3.26036e-08, 3.263224e-08, 
    3.257941e-08, 3.259491e-08, 3.25497e-08, 3.257214e-08, 3.252804e-08, 
    3.250914e-08, 3.24915e-08, 3.247075e-08, 3.264635e-08, 3.265244e-08, 
    3.264156e-08, 3.262645e-08, 3.261251e-08, 3.259396e-08, 3.259208e-08, 
    3.258859e-08, 3.257961e-08, 3.257204e-08, 3.258747e-08, 3.257015e-08, 
    3.263524e-08, 3.260113e-08, 3.265473e-08, 3.263854e-08, 3.262735e-08, 
    3.263228e-08, 3.260677e-08, 3.260075e-08, 3.257629e-08, 3.258895e-08, 
    3.251378e-08, 3.2547e-08, 3.245505e-08, 3.248069e-08, 3.265457e-08, 
    3.264638e-08, 3.261788e-08, 3.263144e-08, 3.259273e-08, 3.258321e-08, 
    3.257548e-08, 3.256557e-08, 3.256452e-08, 3.255866e-08, 3.256827e-08, 
    3.255904e-08, 3.259392e-08, 3.257833e-08, 3.262116e-08, 3.261072e-08, 
    3.261553e-08, 3.262079e-08, 3.260455e-08, 3.258722e-08, 3.258689e-08, 
    3.258133e-08, 3.256558e-08, 3.259258e-08, 3.250942e-08, 3.256067e-08, 
    3.263746e-08, 3.262164e-08, 3.261944e-08, 3.262555e-08, 3.258416e-08, 
    3.259914e-08, 3.255881e-08, 3.256971e-08, 3.255186e-08, 3.256072e-08, 
    3.256202e-08, 3.257343e-08, 3.258052e-08, 3.259845e-08, 3.261306e-08, 
    3.262467e-08, 3.262197e-08, 3.260922e-08, 3.258616e-08, 3.256441e-08, 
    3.256917e-08, 3.255321e-08, 3.259554e-08, 3.257776e-08, 3.258462e-08, 
    3.256675e-08, 3.260596e-08, 3.257243e-08, 3.261452e-08, 3.261083e-08, 
    3.259944e-08, 3.257652e-08, 3.257152e-08, 3.25661e-08, 3.256945e-08, 
    3.258559e-08, 3.258825e-08, 3.259973e-08, 3.260288e-08, 3.261164e-08, 
    3.261887e-08, 3.261225e-08, 3.260529e-08, 3.25856e-08, 3.256784e-08, 
    3.254852e-08, 3.25438e-08, 3.252114e-08, 3.253953e-08, 3.250912e-08, 
    3.253488e-08, 3.249036e-08, 3.257056e-08, 3.253573e-08, 3.259894e-08, 
    3.259213e-08, 3.257978e-08, 3.255156e-08, 3.256683e-08, 3.254899e-08, 
    3.258836e-08, 3.260876e-08, 3.261409e-08, 3.262396e-08, 3.261387e-08, 
    3.261469e-08, 3.260503e-08, 3.260814e-08, 3.258495e-08, 3.25974e-08, 
    3.256205e-08, 3.254914e-08, 3.251279e-08, 3.249052e-08, 3.246793e-08, 
    3.245794e-08, 3.245491e-08, 3.245363e-08,
  5.421948e-11, 5.424386e-11, 5.423915e-11, 5.426019e-11, 5.424793e-11, 
    5.426267e-11, 5.422449e-11, 5.424476e-11, 5.423187e-11, 5.422177e-11, 
    5.430773e-11, 5.426131e-11, 5.435645e-11, 5.432687e-11, 5.440126e-11, 
    5.435176e-11, 5.441125e-11, 5.44e-11, 5.443422e-11, 5.442444e-11, 
    5.446776e-11, 5.443874e-11, 5.449043e-11, 5.446093e-11, 5.446548e-11, 
    5.443775e-11, 5.427082e-11, 5.430191e-11, 5.426894e-11, 5.427339e-11, 
    5.427143e-11, 5.424809e-11, 5.423813e-11, 5.421772e-11, 5.422145e-11, 
    5.42365e-11, 5.427539e-11, 5.426085e-11, 5.429778e-11, 5.429695e-11, 
    5.433784e-11, 5.431942e-11, 5.438807e-11, 5.436863e-11, 5.442485e-11, 
    5.441072e-11, 5.442416e-11, 5.44201e-11, 5.442421e-11, 5.440348e-11, 
    5.441236e-11, 5.439416e-11, 5.432284e-11, 5.434379e-11, 5.428112e-11, 
    5.424508e-11, 5.422535e-11, 5.421122e-11, 5.421321e-11, 5.421699e-11, 
    5.423659e-11, 5.425565e-11, 5.427336e-11, 5.428518e-11, 5.429683e-11, 
    5.433162e-11, 5.435035e-11, 5.439192e-11, 5.438457e-11, 5.439713e-11, 
    5.440931e-11, 5.442956e-11, 5.442625e-11, 5.443513e-11, 5.43969e-11, 
    5.442227e-11, 5.438034e-11, 5.439181e-11, 5.429945e-11, 5.42648e-11, 
    5.425026e-11, 5.424004e-11, 5.421474e-11, 5.423219e-11, 5.42253e-11, 
    5.42418e-11, 5.425219e-11, 5.424707e-11, 5.42855e-11, 5.426994e-11, 
    5.435146e-11, 5.431641e-11, 5.440789e-11, 5.438609e-11, 5.441313e-11, 
    5.439937e-11, 5.44229e-11, 5.440173e-11, 5.443847e-11, 5.44464e-11, 
    5.444097e-11, 5.446199e-11, 5.440054e-11, 5.442411e-11, 5.42469e-11, 
    5.424773e-11, 5.425167e-11, 5.423435e-11, 5.423332e-11, 5.421759e-11, 
    5.423163e-11, 5.423757e-11, 5.425283e-11, 5.4264e-11, 5.427473e-11, 
    5.429829e-11, 5.432446e-11, 5.436113e-11, 5.43875e-11, 5.440511e-11, 
    5.439435e-11, 5.440385e-11, 5.439321e-11, 5.438824e-11, 5.444339e-11, 
    5.441241e-11, 5.445897e-11, 5.445642e-11, 5.443531e-11, 5.445671e-11, 
    5.424832e-11, 5.424352e-11, 5.422666e-11, 5.423986e-11, 5.421588e-11, 
    5.422924e-11, 5.423688e-11, 5.427014e-11, 5.427849e-11, 5.428606e-11, 
    5.430112e-11, 5.432036e-11, 5.4354e-11, 5.438329e-11, 5.441005e-11, 
    5.44081e-11, 5.440878e-11, 5.441469e-11, 5.439996e-11, 5.441711e-11, 
    5.441993e-11, 5.441247e-11, 5.445607e-11, 5.444364e-11, 5.445636e-11, 
    5.444828e-11, 5.42451e-11, 5.425322e-11, 5.424881e-11, 5.425806e-11, 
    5.42512e-11, 5.42832e-11, 5.429292e-11, 5.43385e-11, 5.431995e-11, 
    5.43496e-11, 5.432301e-11, 5.432769e-11, 5.435034e-11, 5.432448e-11, 
    5.438158e-11, 5.434269e-11, 5.441492e-11, 5.437598e-11, 5.441735e-11, 
    5.440993e-11, 5.442226e-11, 5.443323e-11, 5.444712e-11, 5.447255e-11, 
    5.44667e-11, 5.448803e-11, 5.42685e-11, 5.428168e-11, 5.428063e-11, 
    5.429448e-11, 5.43047e-11, 5.432695e-11, 5.436242e-11, 5.434913e-11, 
    5.437364e-11, 5.437852e-11, 5.434133e-11, 5.436408e-11, 5.429058e-11, 
    5.430237e-11, 5.429543e-11, 5.426948e-11, 5.435205e-11, 5.430967e-11, 
    5.438791e-11, 5.436506e-11, 5.443165e-11, 5.439848e-11, 5.446344e-11, 
    5.449084e-11, 5.451706e-11, 5.454706e-11, 5.428899e-11, 5.428002e-11, 
    5.429616e-11, 5.431827e-11, 5.433903e-11, 5.436643e-11, 5.436929e-11, 
    5.437439e-11, 5.438771e-11, 5.439884e-11, 5.43759e-11, 5.440164e-11, 
    5.43049e-11, 5.435577e-11, 5.427653e-11, 5.43003e-11, 5.431701e-11, 
    5.430979e-11, 5.434763e-11, 5.43565e-11, 5.439243e-11, 5.437393e-11, 
    5.448399e-11, 5.44354e-11, 5.457021e-11, 5.453261e-11, 5.427686e-11, 
    5.4289e-11, 5.433102e-11, 5.431106e-11, 5.436832e-11, 5.438233e-11, 
    5.439379e-11, 5.440826e-11, 5.44099e-11, 5.441848e-11, 5.44044e-11, 
    5.441796e-11, 5.436649e-11, 5.438954e-11, 5.432635e-11, 5.434169e-11, 
    5.433467e-11, 5.432689e-11, 5.435088e-11, 5.437623e-11, 5.437694e-11, 
    5.438503e-11, 5.440749e-11, 5.436855e-11, 5.448994e-11, 5.441482e-11, 
    5.430222e-11, 5.432532e-11, 5.432882e-11, 5.431984e-11, 5.438092e-11, 
    5.43588e-11, 5.441829e-11, 5.440228e-11, 5.442855e-11, 5.441549e-11, 
    5.441356e-11, 5.43968e-11, 5.43863e-11, 5.435978e-11, 5.433821e-11, 
    5.432117e-11, 5.432514e-11, 5.434387e-11, 5.437782e-11, 5.440997e-11, 
    5.440291e-11, 5.442656e-11, 5.436417e-11, 5.439028e-11, 5.438014e-11, 
    5.44066e-11, 5.434873e-11, 5.439752e-11, 5.433617e-11, 5.43416e-11, 
    5.435836e-11, 5.439194e-11, 5.43996e-11, 5.440748e-11, 5.440266e-11, 
    5.437871e-11, 5.437486e-11, 5.435799e-11, 5.435325e-11, 5.434043e-11, 
    5.432973e-11, 5.433947e-11, 5.434965e-11, 5.437879e-11, 5.44049e-11, 
    5.443336e-11, 5.444038e-11, 5.447312e-11, 5.444625e-11, 5.449033e-11, 
    5.445251e-11, 5.451807e-11, 5.440058e-11, 5.445174e-11, 5.435918e-11, 
    5.436923e-11, 5.43872e-11, 5.442867e-11, 5.440647e-11, 5.443251e-11, 
    5.437472e-11, 5.434442e-11, 5.433679e-11, 5.432217e-11, 5.433712e-11, 
    5.433591e-11, 5.435019e-11, 5.434561e-11, 5.437976e-11, 5.436144e-11, 
    5.441346e-11, 5.443234e-11, 5.448573e-11, 5.451824e-11, 5.455151e-11, 
    5.456608e-11, 5.457053e-11, 5.457237e-11,
  2.422312e-14, 2.425705e-14, 2.425048e-14, 2.428033e-14, 2.426269e-14, 
    2.428372e-14, 2.423005e-14, 2.425836e-14, 2.424031e-14, 2.422624e-14, 
    2.43458e-14, 2.428185e-14, 2.441276e-14, 2.437187e-14, 2.447476e-14, 
    2.440633e-14, 2.448858e-14, 2.447291e-14, 2.452038e-14, 2.450679e-14, 
    2.456728e-14, 2.452666e-14, 2.459883e-14, 2.455764e-14, 2.456404e-14, 
    2.45253e-14, 2.429483e-14, 2.43378e-14, 2.429225e-14, 2.429839e-14, 
    2.429566e-14, 2.426296e-14, 2.424916e-14, 2.422061e-14, 2.422581e-14, 
    2.424682e-14, 2.430115e-14, 2.428114e-14, 2.433179e-14, 2.433065e-14, 
    2.438698e-14, 2.436158e-14, 2.445638e-14, 2.442946e-14, 2.450736e-14, 
    2.448775e-14, 2.450641e-14, 2.450077e-14, 2.450649e-14, 2.447774e-14, 
    2.449005e-14, 2.446479e-14, 2.436631e-14, 2.439521e-14, 2.430898e-14, 
    2.425891e-14, 2.423127e-14, 2.421158e-14, 2.421436e-14, 2.421965e-14, 
    2.424694e-14, 2.427402e-14, 2.429828e-14, 2.431449e-14, 2.433048e-14, 
    2.43786e-14, 2.440433e-14, 2.446177e-14, 2.44515e-14, 2.446897e-14, 
    2.44858e-14, 2.451393e-14, 2.450931e-14, 2.452168e-14, 2.446858e-14, 
    2.450383e-14, 2.444563e-14, 2.446154e-14, 2.433444e-14, 2.428656e-14, 
    2.426628e-14, 2.425173e-14, 2.421649e-14, 2.42408e-14, 2.423121e-14, 
    2.425412e-14, 2.42691e-14, 2.426146e-14, 2.431494e-14, 2.42936e-14, 
    2.440586e-14, 2.435749e-14, 2.448384e-14, 2.445362e-14, 2.44911e-14, 
    2.447199e-14, 2.45047e-14, 2.447526e-14, 2.452632e-14, 2.453739e-14, 
    2.452981e-14, 2.455905e-14, 2.447362e-14, 2.450638e-14, 2.426125e-14, 
    2.426241e-14, 2.426826e-14, 2.424382e-14, 2.424237e-14, 2.422044e-14, 
    2.423999e-14, 2.424828e-14, 2.427008e-14, 2.428547e-14, 2.430018e-14, 
    2.433253e-14, 2.43686e-14, 2.441917e-14, 2.445557e-14, 2.447996e-14, 
    2.446503e-14, 2.447821e-14, 2.446346e-14, 2.445657e-14, 2.453321e-14, 
    2.449014e-14, 2.455484e-14, 2.455128e-14, 2.452196e-14, 2.455168e-14, 
    2.426324e-14, 2.425652e-14, 2.423308e-14, 2.425142e-14, 2.421806e-14, 
    2.423668e-14, 2.424737e-14, 2.429396e-14, 2.430532e-14, 2.431574e-14, 
    2.43364e-14, 2.436287e-14, 2.440931e-14, 2.444979e-14, 2.44868e-14, 
    2.448409e-14, 2.448504e-14, 2.449327e-14, 2.447284e-14, 2.449663e-14, 
    2.450058e-14, 2.449018e-14, 2.45508e-14, 2.453348e-14, 2.45512e-14, 
    2.453994e-14, 2.425871e-14, 2.42707e-14, 2.426391e-14, 2.427735e-14, 
    2.426758e-14, 2.431189e-14, 2.432526e-14, 2.438797e-14, 2.436233e-14, 
    2.440325e-14, 2.436652e-14, 2.4373e-14, 2.440442e-14, 2.436853e-14, 
    2.444748e-14, 2.43938e-14, 2.449359e-14, 2.443982e-14, 2.449695e-14, 
    2.448664e-14, 2.450375e-14, 2.451904e-14, 2.453834e-14, 2.457385e-14, 
    2.456565e-14, 2.459541e-14, 2.429162e-14, 2.430976e-14, 2.430824e-14, 
    2.432728e-14, 2.434134e-14, 2.437193e-14, 2.442091e-14, 2.440251e-14, 
    2.443637e-14, 2.444314e-14, 2.439175e-14, 2.442323e-14, 2.432196e-14, 
    2.433824e-14, 2.43286e-14, 2.429301e-14, 2.440665e-14, 2.434827e-14, 
    2.445616e-14, 2.442454e-14, 2.451685e-14, 2.447086e-14, 2.456111e-14, 
    2.459951e-14, 2.4636e-14, 2.467825e-14, 2.431974e-14, 2.430741e-14, 
    2.432956e-14, 2.436008e-14, 2.438862e-14, 2.442645e-14, 2.443036e-14, 
    2.443743e-14, 2.445583e-14, 2.447126e-14, 2.443959e-14, 2.447513e-14, 
    2.434187e-14, 2.441175e-14, 2.430268e-14, 2.433541e-14, 2.435832e-14, 
    2.434834e-14, 2.440043e-14, 2.441268e-14, 2.446245e-14, 2.443676e-14, 
    2.458997e-14, 2.452216e-14, 2.471068e-14, 2.465793e-14, 2.430308e-14, 
    2.431974e-14, 2.437761e-14, 2.435008e-14, 2.442902e-14, 2.444842e-14, 
    2.446426e-14, 2.448438e-14, 2.448661e-14, 2.449854e-14, 2.447898e-14, 
    2.44978e-14, 2.442653e-14, 2.445839e-14, 2.437108e-14, 2.439229e-14, 
    2.438256e-14, 2.437183e-14, 2.440493e-14, 2.444007e-14, 2.444094e-14, 
    2.445219e-14, 2.448368e-14, 2.442934e-14, 2.45985e-14, 2.449381e-14, 
    2.433789e-14, 2.436982e-14, 2.437453e-14, 2.436213e-14, 2.444647e-14, 
    2.441589e-14, 2.449827e-14, 2.447603e-14, 2.45125e-14, 2.449436e-14, 
    2.449169e-14, 2.446843e-14, 2.445392e-14, 2.441727e-14, 2.438749e-14, 
    2.436395e-14, 2.436943e-14, 2.43953e-14, 2.444225e-14, 2.448676e-14, 
    2.447699e-14, 2.450973e-14, 2.442329e-14, 2.445947e-14, 2.444545e-14, 
    2.448204e-14, 2.440199e-14, 2.446979e-14, 2.438463e-14, 2.439212e-14, 
    2.441528e-14, 2.446185e-14, 2.447232e-14, 2.44833e-14, 2.447655e-14, 
    2.444347e-14, 2.44381e-14, 2.441475e-14, 2.440825e-14, 2.43905e-14, 
    2.437575e-14, 2.438919e-14, 2.440329e-14, 2.444353e-14, 2.447972e-14, 
    2.451924e-14, 2.452895e-14, 2.457483e-14, 2.453732e-14, 2.459906e-14, 
    2.454632e-14, 2.463775e-14, 2.44739e-14, 2.454501e-14, 2.441638e-14, 
    2.443026e-14, 2.445525e-14, 2.451282e-14, 2.448186e-14, 2.451813e-14, 
    2.44379e-14, 2.439613e-14, 2.438548e-14, 2.436536e-14, 2.438594e-14, 
    2.438427e-14, 2.440396e-14, 2.439764e-14, 2.444487e-14, 2.44195e-14, 
    2.449159e-14, 2.451787e-14, 2.459225e-14, 2.463778e-14, 2.468434e-14, 
    2.470483e-14, 2.471108e-14, 2.471369e-14,
  3.219115e-18, 3.226515e-18, 3.22508e-18, 3.231465e-18, 3.227743e-18, 
    3.232164e-18, 3.220622e-18, 3.226802e-18, 3.22286e-18, 3.219792e-18, 
    3.244979e-18, 3.231778e-18, 3.258817e-18, 3.250353e-18, 3.271669e-18, 
    3.257487e-18, 3.274537e-18, 3.27128e-18, 3.281139e-18, 3.278314e-18, 
    3.291344e-18, 3.282444e-18, 3.298332e-18, 3.289205e-18, 3.290624e-18, 
    3.282162e-18, 3.23445e-18, 3.243327e-18, 3.23392e-18, 3.235186e-18, 
    3.234622e-18, 3.227805e-18, 3.224796e-18, 3.218563e-18, 3.219697e-18, 
    3.224283e-18, 3.235756e-18, 3.23163e-18, 3.242073e-18, 3.241837e-18, 
    3.253479e-18, 3.248226e-18, 3.267852e-18, 3.26227e-18, 3.278432e-18, 
    3.27436e-18, 3.278237e-18, 3.277064e-18, 3.278253e-18, 3.272282e-18, 
    3.274838e-18, 3.269595e-18, 3.249205e-18, 3.255182e-18, 3.23737e-18, 
    3.226928e-18, 3.22089e-18, 3.216597e-18, 3.217204e-18, 3.218356e-18, 
    3.224309e-18, 3.230163e-18, 3.235161e-18, 3.238504e-18, 3.241803e-18, 
    3.251753e-18, 3.257072e-18, 3.268971e-18, 3.266839e-18, 3.270465e-18, 
    3.273956e-18, 3.279799e-18, 3.278839e-18, 3.281411e-18, 3.270382e-18, 
    3.277703e-18, 3.265621e-18, 3.26892e-18, 3.242633e-18, 3.232746e-18, 
    3.228532e-18, 3.225353e-18, 3.217669e-18, 3.22297e-18, 3.220877e-18, 
    3.225872e-18, 3.229135e-18, 3.227475e-18, 3.238596e-18, 3.234197e-18, 
    3.257388e-18, 3.247384e-18, 3.273548e-18, 3.267278e-18, 3.275055e-18, 
    3.271088e-18, 3.277881e-18, 3.271768e-18, 3.282374e-18, 3.284723e-18, 
    3.283102e-18, 3.289514e-18, 3.271427e-18, 3.278231e-18, 3.227428e-18, 
    3.227683e-18, 3.228953e-18, 3.223628e-18, 3.223311e-18, 3.218529e-18, 
    3.22279e-18, 3.224601e-18, 3.229346e-18, 3.232522e-18, 3.235553e-18, 
    3.242226e-18, 3.249679e-18, 3.260142e-18, 3.267684e-18, 3.272741e-18, 
    3.269644e-18, 3.272378e-18, 3.269319e-18, 3.267889e-18, 3.283811e-18, 
    3.274858e-18, 3.288583e-18, 3.287793e-18, 3.28147e-18, 3.287882e-18, 
    3.227863e-18, 3.226395e-18, 3.221284e-18, 3.225283e-18, 3.218009e-18, 
    3.222071e-18, 3.224403e-18, 3.234274e-18, 3.236613e-18, 3.238762e-18, 
    3.243025e-18, 3.248494e-18, 3.2581e-18, 3.266486e-18, 3.274162e-18, 
    3.2736e-18, 3.273797e-18, 3.275506e-18, 3.271264e-18, 3.276204e-18, 
    3.277027e-18, 3.274865e-18, 3.287687e-18, 3.283864e-18, 3.287776e-18, 
    3.285283e-18, 3.226874e-18, 3.22948e-18, 3.228009e-18, 3.23085e-18, 
    3.228808e-18, 3.237972e-18, 3.240732e-18, 3.253687e-18, 3.248383e-18, 
    3.256847e-18, 3.249247e-18, 3.250589e-18, 3.257094e-18, 3.249662e-18, 
    3.26601e-18, 3.254894e-18, 3.275573e-18, 3.264425e-18, 3.276271e-18, 
    3.274128e-18, 3.277683e-18, 3.280861e-18, 3.284931e-18, 3.292796e-18, 
    3.290976e-18, 3.297572e-18, 3.233789e-18, 3.237531e-18, 3.237214e-18, 
    3.241142e-18, 3.244047e-18, 3.250364e-18, 3.260501e-18, 3.25669e-18, 
    3.263702e-18, 3.265106e-18, 3.254463e-18, 3.260982e-18, 3.240047e-18, 
    3.24341e-18, 3.241416e-18, 3.234077e-18, 3.25755e-18, 3.24548e-18, 
    3.267806e-18, 3.261251e-18, 3.280406e-18, 3.270858e-18, 3.289972e-18, 
    3.298489e-18, 3.306577e-18, 3.315974e-18, 3.239589e-18, 3.237043e-18, 
    3.241613e-18, 3.247921e-18, 3.253817e-18, 3.261648e-18, 3.262457e-18, 
    3.263922e-18, 3.267735e-18, 3.270936e-18, 3.264373e-18, 3.27174e-18, 
    3.244164e-18, 3.258605e-18, 3.23607e-18, 3.242826e-18, 3.247554e-18, 
    3.245493e-18, 3.256258e-18, 3.258795e-18, 3.269112e-18, 3.263783e-18, 
    3.296374e-18, 3.281515e-18, 3.323183e-18, 3.311454e-18, 3.236151e-18, 
    3.239586e-18, 3.251542e-18, 3.245851e-18, 3.262178e-18, 3.266201e-18, 
    3.269483e-18, 3.273662e-18, 3.274123e-18, 3.276602e-18, 3.272538e-18, 
    3.276446e-18, 3.261665e-18, 3.268268e-18, 3.250189e-18, 3.254575e-18, 
    3.252561e-18, 3.250344e-18, 3.25719e-18, 3.264473e-18, 3.26465e-18, 
    3.266984e-18, 3.273531e-18, 3.262245e-18, 3.298277e-18, 3.275632e-18, 
    3.243333e-18, 3.249934e-18, 3.250903e-18, 3.24834e-18, 3.265797e-18, 
    3.259461e-18, 3.276545e-18, 3.271926e-18, 3.279501e-18, 3.275733e-18, 
    3.275178e-18, 3.27035e-18, 3.26734e-18, 3.259747e-18, 3.253584e-18, 
    3.248714e-18, 3.249847e-18, 3.2552e-18, 3.264924e-18, 3.274155e-18, 
    3.272129e-18, 3.278925e-18, 3.260992e-18, 3.268494e-18, 3.265586e-18, 
    3.273174e-18, 3.256584e-18, 3.270646e-18, 3.25299e-18, 3.254539e-18, 
    3.259335e-18, 3.268989e-18, 3.271157e-18, 3.273437e-18, 3.272035e-18, 
    3.265175e-18, 3.264061e-18, 3.259224e-18, 3.257879e-18, 3.254203e-18, 
    3.251153e-18, 3.253935e-18, 3.256854e-18, 3.265186e-18, 3.272696e-18, 
    3.280903e-18, 3.282922e-18, 3.293022e-18, 3.284715e-18, 3.298402e-18, 
    3.28672e-18, 3.30698e-18, 3.271492e-18, 3.286419e-18, 3.25956e-18, 
    3.262437e-18, 3.267621e-18, 3.279573e-18, 3.273138e-18, 3.280675e-18, 
    3.264019e-18, 3.255374e-18, 3.253166e-18, 3.249006e-18, 3.253261e-18, 
    3.252915e-18, 3.256989e-18, 3.255681e-18, 3.265464e-18, 3.260207e-18, 
    3.275159e-18, 3.280621e-18, 3.296872e-18, 3.306978e-18, 3.317319e-18, 
    3.321879e-18, 3.323269e-18, 3.32385e-18,
  1.347684e-22, 1.352459e-22, 1.351532e-22, 1.355537e-22, 1.353251e-22, 
    1.35596e-22, 1.348655e-22, 1.352646e-22, 1.350099e-22, 1.348119e-22, 
    1.363713e-22, 1.355726e-22, 1.372091e-22, 1.36696e-22, 1.379891e-22, 
    1.371286e-22, 1.381633e-22, 1.379652e-22, 1.385665e-22, 1.383927e-22, 
    1.392145e-22, 1.38649e-22, 1.396586e-22, 1.390782e-22, 1.391685e-22, 
    1.386312e-22, 1.357339e-22, 1.362714e-22, 1.357019e-22, 1.357785e-22, 
    1.357443e-22, 1.353292e-22, 1.351352e-22, 1.347326e-22, 1.348058e-22, 
    1.351019e-22, 1.35813e-22, 1.355636e-22, 1.361947e-22, 1.361804e-22, 
    1.368853e-22, 1.365671e-22, 1.37757e-22, 1.374181e-22, 1.383999e-22, 
    1.381523e-22, 1.383881e-22, 1.383166e-22, 1.38389e-22, 1.380261e-22, 
    1.381814e-22, 1.378628e-22, 1.366264e-22, 1.369885e-22, 1.359104e-22, 
    1.352731e-22, 1.348828e-22, 1.346059e-22, 1.34645e-22, 1.347194e-22, 
    1.351036e-22, 1.35475e-22, 1.357768e-22, 1.359789e-22, 1.361783e-22, 
    1.367812e-22, 1.371033e-22, 1.378251e-22, 1.376954e-22, 1.379158e-22, 
    1.381277e-22, 1.38483e-22, 1.384246e-22, 1.385839e-22, 1.379106e-22, 
    1.383557e-22, 1.376214e-22, 1.378219e-22, 1.362294e-22, 1.35631e-22, 
    1.353756e-22, 1.351709e-22, 1.34675e-22, 1.350171e-22, 1.348821e-22, 
    1.352042e-22, 1.354124e-22, 1.353077e-22, 1.359844e-22, 1.357186e-22, 
    1.371224e-22, 1.365163e-22, 1.38103e-22, 1.377221e-22, 1.381945e-22, 
    1.379535e-22, 1.383665e-22, 1.379947e-22, 1.386447e-22, 1.387935e-22, 
    1.386908e-22, 1.390976e-22, 1.379741e-22, 1.383877e-22, 1.353047e-22, 
    1.353212e-22, 1.354012e-22, 1.350596e-22, 1.350391e-22, 1.347305e-22, 
    1.350054e-22, 1.351223e-22, 1.354254e-22, 1.356174e-22, 1.358006e-22, 
    1.36204e-22, 1.366552e-22, 1.372892e-22, 1.377468e-22, 1.380539e-22, 
    1.378657e-22, 1.380318e-22, 1.37846e-22, 1.377591e-22, 1.387357e-22, 
    1.381827e-22, 1.390385e-22, 1.389883e-22, 1.385876e-22, 1.38994e-22, 
    1.353328e-22, 1.35238e-22, 1.349082e-22, 1.351662e-22, 1.346969e-22, 
    1.34959e-22, 1.351097e-22, 1.357234e-22, 1.358646e-22, 1.359945e-22, 
    1.362523e-22, 1.365833e-22, 1.371654e-22, 1.376741e-22, 1.381402e-22, 
    1.381061e-22, 1.381181e-22, 1.38222e-22, 1.379642e-22, 1.382644e-22, 
    1.383145e-22, 1.38183e-22, 1.389815e-22, 1.387388e-22, 1.389872e-22, 
    1.388289e-22, 1.352689e-22, 1.354337e-22, 1.353423e-22, 1.355165e-22, 
    1.353923e-22, 1.35947e-22, 1.361139e-22, 1.368981e-22, 1.365766e-22, 
    1.370895e-22, 1.366289e-22, 1.367102e-22, 1.371049e-22, 1.36654e-22, 
    1.376454e-22, 1.369714e-22, 1.382261e-22, 1.375494e-22, 1.382685e-22, 
    1.381382e-22, 1.383543e-22, 1.385491e-22, 1.388066e-22, 1.393064e-22, 
    1.391907e-22, 1.3961e-22, 1.35694e-22, 1.359202e-22, 1.359009e-22, 
    1.361384e-22, 1.363142e-22, 1.366965e-22, 1.373109e-22, 1.370798e-22, 
    1.37505e-22, 1.375903e-22, 1.369447e-22, 1.373402e-22, 1.360723e-22, 
    1.362758e-22, 1.361551e-22, 1.357115e-22, 1.371322e-22, 1.364011e-22, 
    1.377542e-22, 1.373564e-22, 1.385203e-22, 1.379397e-22, 1.391269e-22, 
    1.396688e-22, 1.401832e-22, 1.407827e-22, 1.360445e-22, 1.358905e-22, 
    1.361668e-22, 1.365488e-22, 1.369057e-22, 1.373805e-22, 1.374295e-22, 
    1.375185e-22, 1.377498e-22, 1.379442e-22, 1.37546e-22, 1.379931e-22, 
    1.363219e-22, 1.371961e-22, 1.358318e-22, 1.362406e-22, 1.365266e-22, 
    1.364017e-22, 1.370536e-22, 1.372074e-22, 1.378336e-22, 1.375099e-22, 
    1.395344e-22, 1.385907e-22, 1.412425e-22, 1.404943e-22, 1.358366e-22, 
    1.360443e-22, 1.36768e-22, 1.364234e-22, 1.374126e-22, 1.376567e-22, 
    1.37856e-22, 1.3811e-22, 1.381379e-22, 1.382887e-22, 1.380416e-22, 
    1.382791e-22, 1.373815e-22, 1.377822e-22, 1.366859e-22, 1.369517e-22, 
    1.368296e-22, 1.366952e-22, 1.3711e-22, 1.375521e-22, 1.375625e-22, 
    1.377044e-22, 1.381029e-22, 1.374166e-22, 1.39656e-22, 1.382305e-22, 
    1.362709e-22, 1.366708e-22, 1.367292e-22, 1.365739e-22, 1.376322e-22, 
    1.372478e-22, 1.382851e-22, 1.380044e-22, 1.384649e-22, 1.382358e-22, 
    1.382021e-22, 1.379086e-22, 1.377259e-22, 1.372652e-22, 1.368917e-22, 
    1.365965e-22, 1.366652e-22, 1.369896e-22, 1.375794e-22, 1.3814e-22, 
    1.380169e-22, 1.384298e-22, 1.373406e-22, 1.37796e-22, 1.376196e-22, 
    1.380802e-22, 1.370734e-22, 1.379275e-22, 1.368555e-22, 1.369494e-22, 
    1.372402e-22, 1.378263e-22, 1.379577e-22, 1.380963e-22, 1.38011e-22, 
    1.375946e-22, 1.375269e-22, 1.372334e-22, 1.371519e-22, 1.36929e-22, 
    1.367443e-22, 1.369128e-22, 1.370899e-22, 1.375952e-22, 1.380513e-22, 
    1.385518e-22, 1.386793e-22, 1.393214e-22, 1.387934e-22, 1.396641e-22, 
    1.389215e-22, 1.402098e-22, 1.379785e-22, 1.389017e-22, 1.372538e-22, 
    1.374282e-22, 1.377432e-22, 1.384697e-22, 1.380781e-22, 1.385376e-22, 
    1.375243e-22, 1.370003e-22, 1.368662e-22, 1.366143e-22, 1.368719e-22, 
    1.36851e-22, 1.370979e-22, 1.370186e-22, 1.37612e-22, 1.37293e-22, 
    1.38201e-22, 1.38534e-22, 1.395657e-22, 1.402091e-22, 1.40868e-22, 
    1.411591e-22, 1.412479e-22, 1.41285e-22,
  1.8411e-27, 1.85035e-27, 1.84855e-27, 1.856196e-27, 1.851885e-27, 
    1.856985e-27, 1.84297e-27, 1.850714e-27, 1.84577e-27, 1.84193e-27, 
    1.871502e-27, 1.856549e-27, 1.887205e-27, 1.877575e-27, 1.901867e-27, 
    1.885696e-27, 1.905144e-27, 1.901412e-27, 1.912742e-27, 1.90946e-27, 
    1.924866e-27, 1.914306e-27, 1.933133e-27, 1.922327e-27, 1.924009e-27, 
    1.913969e-27, 1.859562e-27, 1.86963e-27, 1.858964e-27, 1.860397e-27, 
    1.859757e-27, 1.851966e-27, 1.848205e-27, 1.840426e-27, 1.841812e-27, 
    1.847555e-27, 1.861042e-27, 1.856377e-27, 1.868181e-27, 1.867914e-27, 
    1.881124e-27, 1.875157e-27, 1.897496e-27, 1.891126e-27, 1.909595e-27, 
    1.904933e-27, 1.909373e-27, 1.908028e-27, 1.909391e-27, 1.902559e-27, 
    1.905483e-27, 1.899486e-27, 1.876271e-27, 1.883063e-27, 1.862864e-27, 
    1.850883e-27, 1.843306e-27, 1.838054e-27, 1.838786e-27, 1.840181e-27, 
    1.847589e-27, 1.854721e-27, 1.860362e-27, 1.864142e-27, 1.867875e-27, 
    1.879181e-27, 1.885219e-27, 1.89878e-27, 1.896338e-27, 1.900485e-27, 
    1.904471e-27, 1.911164e-27, 1.910062e-27, 1.913072e-27, 1.900384e-27, 
    1.908765e-27, 1.894945e-27, 1.898715e-27, 1.868846e-27, 1.857636e-27, 
    1.852861e-27, 1.848894e-27, 1.839349e-27, 1.845911e-27, 1.843293e-27, 
    1.849537e-27, 1.853549e-27, 1.851546e-27, 1.864246e-27, 1.859274e-27, 
    1.885578e-27, 1.874208e-27, 1.904006e-27, 1.89684e-27, 1.905728e-27, 
    1.901191e-27, 1.908968e-27, 1.901967e-27, 1.914225e-27, 1.917033e-27, 
    1.9151e-27, 1.922686e-27, 1.901578e-27, 1.909369e-27, 1.851489e-27, 
    1.851808e-27, 1.853336e-27, 1.846736e-27, 1.846337e-27, 1.840387e-27, 
    1.845681e-27, 1.847951e-27, 1.853793e-27, 1.857384e-27, 1.860808e-27, 
    1.868357e-27, 1.876813e-27, 1.888708e-27, 1.897303e-27, 1.903081e-27, 
    1.899539e-27, 1.902665e-27, 1.899169e-27, 1.897535e-27, 1.915953e-27, 
    1.905507e-27, 1.921586e-27, 1.920652e-27, 1.913144e-27, 1.920757e-27, 
    1.852034e-27, 1.850192e-27, 1.843798e-27, 1.8488e-27, 1.839758e-27, 
    1.844784e-27, 1.847709e-27, 1.859368e-27, 1.862004e-27, 1.864437e-27, 
    1.86926e-27, 1.875462e-27, 1.886383e-27, 1.895939e-27, 1.904705e-27, 
    1.904062e-27, 1.904288e-27, 1.906246e-27, 1.901393e-27, 1.907044e-27, 
    1.90799e-27, 1.905512e-27, 1.920526e-27, 1.91601e-27, 1.920632e-27, 
    1.917687e-27, 1.850792e-27, 1.85395e-27, 1.852217e-27, 1.855498e-27, 
    1.85317e-27, 1.86355e-27, 1.866674e-27, 1.881369e-27, 1.875337e-27, 
    1.884958e-27, 1.876316e-27, 1.877842e-27, 1.885254e-27, 1.876785e-27, 
    1.895402e-27, 1.882745e-27, 1.906322e-27, 1.893602e-27, 1.907121e-27, 
    1.904667e-27, 1.908736e-27, 1.912412e-27, 1.917273e-27, 1.926574e-27, 
    1.924418e-27, 1.932226e-27, 1.858814e-27, 1.863048e-27, 1.862683e-27, 
    1.867128e-27, 1.87042e-27, 1.877583e-27, 1.889113e-27, 1.884773e-27, 
    1.892758e-27, 1.894361e-27, 1.882238e-27, 1.889665e-27, 1.865893e-27, 
    1.869706e-27, 1.867441e-27, 1.859143e-27, 1.885761e-27, 1.872052e-27, 
    1.897444e-27, 1.889967e-27, 1.911867e-27, 1.900936e-27, 1.923231e-27, 
    1.933328e-27, 1.942911e-27, 1.954365e-27, 1.865371e-27, 1.862489e-27, 
    1.86766e-27, 1.874819e-27, 1.881508e-27, 1.890421e-27, 1.89134e-27, 
    1.893012e-27, 1.89736e-27, 1.901017e-27, 1.893532e-27, 1.901936e-27, 
    1.870575e-27, 1.886959e-27, 1.861393e-27, 1.869047e-27, 1.8744e-27, 
    1.872059e-27, 1.88428e-27, 1.887167e-27, 1.898939e-27, 1.892851e-27, 
    1.930824e-27, 1.913206e-27, 1.963201e-27, 1.948825e-27, 1.861481e-27, 
    1.865365e-27, 1.878927e-27, 1.872465e-27, 1.891022e-27, 1.895611e-27, 
    1.899356e-27, 1.904138e-27, 1.904662e-27, 1.907502e-27, 1.902848e-27, 
    1.907321e-27, 1.89044e-27, 1.897969e-27, 1.877383e-27, 1.88237e-27, 
    1.880077e-27, 1.877559e-27, 1.88534e-27, 1.893648e-27, 1.89384e-27, 
    1.896508e-27, 1.90402e-27, 1.891098e-27, 1.933099e-27, 1.90642e-27, 
    1.869608e-27, 1.877106e-27, 1.878196e-27, 1.875284e-27, 1.89515e-27, 
    1.887928e-27, 1.907434e-27, 1.902149e-27, 1.91082e-27, 1.906505e-27, 
    1.905871e-27, 1.900347e-27, 1.896911e-27, 1.888256e-27, 1.881245e-27, 
    1.875708e-27, 1.876995e-27, 1.883082e-27, 1.89416e-27, 1.904703e-27, 
    1.902387e-27, 1.91016e-27, 1.88967e-27, 1.898232e-27, 1.894914e-27, 
    1.903577e-27, 1.884655e-27, 1.900716e-27, 1.880564e-27, 1.882326e-27, 
    1.887785e-27, 1.898804e-27, 1.90127e-27, 1.903881e-27, 1.902272e-27, 
    1.894445e-27, 1.893171e-27, 1.887656e-27, 1.886129e-27, 1.881943e-27, 
    1.878478e-27, 1.88164e-27, 1.884964e-27, 1.894454e-27, 1.903034e-27, 
    1.912464e-27, 1.91488e-27, 1.92686e-27, 1.917036e-27, 1.93325e-27, 
    1.919428e-27, 1.943421e-27, 1.901671e-27, 1.919051e-27, 1.888039e-27, 
    1.891315e-27, 1.897239e-27, 1.910917e-27, 1.903536e-27, 1.912198e-27, 
    1.893122e-27, 1.883285e-27, 1.880765e-27, 1.876041e-27, 1.880873e-27, 
    1.88048e-27, 1.885111e-27, 1.883623e-27, 1.89477e-27, 1.888775e-27, 
    1.905851e-27, 1.91213e-27, 1.931401e-27, 1.943401e-27, 1.955997e-27, 
    1.961594e-27, 1.963301e-27, 1.964014e-27,
  8.105283e-33, 8.160627e-33, 8.14984e-33, 8.195232e-33, 8.169814e-33, 
    8.199858e-33, 8.116445e-33, 8.162813e-33, 8.133197e-33, 8.110224e-33, 
    8.286118e-33, 8.197298e-33, 8.381051e-33, 8.322751e-33, 8.470025e-33, 
    8.371918e-33, 8.489948e-33, 8.467239e-33, 8.536091e-33, 8.516189e-33, 
    8.608125e-33, 8.545482e-33, 8.657065e-33, 8.593084e-33, 8.603041e-33, 
    8.54346e-33, 8.214974e-33, 8.27482e-33, 8.211465e-33, 8.219885e-33, 
    8.216119e-33, 8.170307e-33, 8.1478e-33, 8.101276e-33, 8.109517e-33, 
    8.143894e-33, 8.223675e-33, 8.196275e-33, 8.266006e-33, 8.264395e-33, 
    8.344215e-33, 8.308133e-33, 8.443449e-33, 8.404789e-33, 8.517013e-33, 
    8.488647e-33, 8.515668e-33, 8.507474e-33, 8.515775e-33, 8.474214e-33, 
    8.491993e-33, 8.455529e-33, 8.314868e-33, 8.355954e-33, 8.234372e-33, 
    8.163848e-33, 8.118464e-33, 8.087205e-33, 8.09155e-33, 8.099828e-33, 
    8.144094e-33, 8.186566e-33, 8.219668e-33, 8.241873e-33, 8.264162e-33, 
    8.332503e-33, 8.369023e-33, 8.451257e-33, 8.436411e-33, 8.461615e-33, 
    8.485833e-33, 8.526573e-33, 8.519862e-33, 8.538081e-33, 8.460986e-33, 
    8.511974e-33, 8.427952e-33, 8.450849e-33, 8.270094e-33, 8.203667e-33, 
    8.175656e-33, 8.151905e-33, 8.094888e-33, 8.134051e-33, 8.118383e-33, 
    8.155747e-33, 8.179682e-33, 8.167777e-33, 8.242481e-33, 8.213282e-33, 
    8.371192e-33, 8.302406e-33, 8.483005e-33, 8.43946e-33, 8.493482e-33, 
    8.465885e-33, 8.513206e-33, 8.470606e-33, 8.545e-33, 8.561787e-33, 
    8.550263e-33, 8.595193e-33, 8.468245e-33, 8.515648e-33, 8.167438e-33, 
    8.169356e-33, 8.178423e-33, 8.138989e-33, 8.136601e-33, 8.101043e-33, 
    8.132665e-33, 8.146259e-33, 8.181109e-33, 8.202187e-33, 8.22229e-33, 
    8.267078e-33, 8.318156e-33, 8.39015e-33, 8.442274e-33, 8.477374e-33, 
    8.455849e-33, 8.474849e-33, 8.453604e-33, 8.443672e-33, 8.555392e-33, 
    8.492147e-33, 8.588691e-33, 8.583163e-33, 8.538514e-33, 8.583787e-33, 
    8.170705e-33, 8.159668e-33, 8.121401e-33, 8.151334e-33, 8.097315e-33, 
    8.127303e-33, 8.144817e-33, 8.213848e-33, 8.229309e-33, 8.243609e-33, 
    8.272524e-33, 8.309975e-33, 8.376058e-33, 8.433999e-33, 8.487252e-33, 
    8.483344e-33, 8.484717e-33, 8.496633e-33, 8.467119e-33, 8.50149e-33, 
    8.507252e-33, 8.492164e-33, 8.582422e-33, 8.55572e-33, 8.583045e-33, 
    8.565638e-33, 8.163259e-33, 8.182039e-33, 8.171799e-33, 8.191123e-33, 
    8.177453e-33, 8.238415e-33, 8.256949e-33, 8.345717e-33, 8.309225e-33, 
    8.36743e-33, 8.315136e-33, 8.324368e-33, 8.369251e-33, 8.317967e-33, 
    8.430756e-33, 8.354053e-33, 8.497097e-33, 8.419848e-33, 8.501955e-33, 
    8.487021e-33, 8.511782e-33, 8.534115e-33, 8.563194e-33, 8.61821e-33, 
    8.605449e-33, 8.651679e-33, 8.210579e-33, 8.235455e-33, 8.233298e-33, 
    8.259661e-33, 8.279527e-33, 8.322792e-33, 8.392595e-33, 8.366292e-33, 
    8.414683e-33, 8.424417e-33, 8.350945e-33, 8.395946e-33, 8.252218e-33, 
    8.275239e-33, 8.261552e-33, 8.212517e-33, 8.372295e-33, 8.2894e-33, 
    8.443131e-33, 8.397767e-33, 8.530845e-33, 8.464362e-33, 8.598423e-33, 
    8.658237e-33, 8.715064e-33, 8.783505e-33, 8.249101e-33, 8.23216e-33, 
    8.262864e-33, 8.306111e-33, 8.346538e-33, 8.40052e-33, 8.406083e-33, 
    8.416228e-33, 8.442611e-33, 8.464831e-33, 8.419403e-33, 8.470414e-33, 
    8.280511e-33, 8.379545e-33, 8.22573e-33, 8.271264e-33, 8.303572e-33, 
    8.289422e-33, 8.363301e-33, 8.380792e-33, 8.452219e-33, 8.415245e-33, 
    8.643405e-33, 8.538901e-33, 8.837109e-33, 8.750351e-33, 8.22624e-33, 
    8.24906e-33, 8.330935e-33, 8.291872e-33, 8.404156e-33, 8.432002e-33, 
    8.454735e-33, 8.483817e-33, 8.48699e-33, 8.504278e-33, 8.475962e-33, 
    8.503172e-33, 8.400635e-33, 8.446318e-33, 8.321578e-33, 8.351752e-33, 
    8.337871e-33, 8.322642e-33, 8.369725e-33, 8.420106e-33, 8.421247e-33, 
    8.437455e-33, 8.483176e-33, 8.404615e-33, 8.656928e-33, 8.497762e-33, 
    8.274619e-33, 8.319937e-33, 8.326503e-33, 8.308893e-33, 8.429204e-33, 
    8.38541e-33, 8.503864e-33, 8.471708e-33, 8.524473e-33, 8.498208e-33, 
    8.494348e-33, 8.460757e-33, 8.439892e-33, 8.387402e-33, 8.344943e-33, 
    8.311453e-33, 8.319233e-33, 8.356063e-33, 8.423211e-33, 8.48725e-33, 
    8.473174e-33, 8.520453e-33, 8.395963e-33, 8.447922e-33, 8.427783e-33, 
    8.480398e-33, 8.36558e-33, 8.463075e-33, 8.340813e-33, 8.351477e-33, 
    8.384543e-33, 8.451416e-33, 8.466369e-33, 8.482252e-33, 8.472461e-33, 
    8.424934e-33, 8.417199e-33, 8.383754e-33, 8.374511e-33, 8.349159e-33, 
    8.328196e-33, 8.347332e-33, 8.36746e-33, 8.42498e-33, 8.477102e-33, 
    8.534432e-33, 8.54893e-33, 8.619937e-33, 8.561831e-33, 8.657824e-33, 
    8.57602e-33, 8.718149e-33, 8.468848e-33, 8.573751e-33, 8.386071e-33, 
    8.405933e-33, 8.441906e-33, 8.525094e-33, 8.480151e-33, 8.53285e-33, 
    8.416901e-33, 8.357306e-33, 8.342029e-33, 8.313474e-33, 8.342683e-33, 
    8.340307e-33, 8.368338e-33, 8.359324e-33, 8.426896e-33, 8.390537e-33, 
    8.494235e-33, 8.532435e-33, 8.646801e-33, 8.717994e-33, 8.793245e-33, 
    8.827244e-33, 8.837711e-33, 8.842089e-33,
  1.16866e-38, 1.179981e-38, 1.177771e-38, 1.187028e-38, 1.181863e-38, 
    1.187966e-38, 1.170941e-38, 1.180431e-38, 1.174365e-38, 1.169671e-38, 
    1.205556e-38, 1.187447e-38, 1.225076e-38, 1.213064e-38, 1.243891e-38, 
    1.223193e-38, 1.248139e-38, 1.243293e-38, 1.257987e-38, 1.253742e-38, 
    1.273131e-38, 1.259973e-38, 1.283425e-38, 1.26997e-38, 1.272061e-38, 
    1.259546e-38, 1.191032e-38, 1.203242e-38, 1.19032e-38, 1.192031e-38, 
    1.191265e-38, 1.181965e-38, 1.177357e-38, 1.167829e-38, 1.169526e-38, 
    1.176555e-38, 1.192802e-38, 1.187237e-38, 1.201426e-38, 1.201096e-38, 
    1.217479e-38, 1.210061e-38, 1.23823e-38, 1.230024e-38, 1.253918e-38, 
    1.247857e-38, 1.253631e-38, 1.251878e-38, 1.253654e-38, 1.244779e-38, 
    1.248572e-38, 1.240799e-38, 1.211445e-38, 1.219897e-38, 1.194975e-38, 
    1.180646e-38, 1.171354e-38, 1.164921e-38, 1.165819e-38, 1.167531e-38, 
    1.176596e-38, 1.185269e-38, 1.191984e-38, 1.196499e-38, 1.201049e-38, 
    1.215076e-38, 1.222594e-38, 1.239893e-38, 1.236733e-38, 1.242097e-38, 
    1.247257e-38, 1.255966e-38, 1.254529e-38, 1.258409e-38, 1.24196e-38, 
    1.252843e-38, 1.234936e-38, 1.239803e-38, 1.202275e-38, 1.188737e-38, 
    1.183062e-38, 1.178194e-38, 1.166509e-38, 1.174541e-38, 1.171339e-38, 
    1.178979e-38, 1.183873e-38, 1.181444e-38, 1.196623e-38, 1.190688e-38, 
    1.223041e-38, 1.208887e-38, 1.246653e-38, 1.237382e-38, 1.248889e-38, 
    1.243003e-38, 1.253106e-38, 1.244009e-38, 1.259872e-38, 1.263415e-38, 
    1.260987e-38, 1.27041e-38, 1.243506e-38, 1.253629e-38, 1.181375e-38, 
    1.181769e-38, 1.183618e-38, 1.175551e-38, 1.175062e-38, 1.167781e-38, 
    1.174256e-38, 1.177038e-38, 1.184162e-38, 1.188436e-38, 1.192518e-38, 
    1.201647e-38, 1.212121e-38, 1.226953e-38, 1.23798e-38, 1.245452e-38, 
    1.240866e-38, 1.244913e-38, 1.240388e-38, 1.238276e-38, 1.262075e-38, 
    1.248606e-38, 1.269047e-38, 1.267888e-38, 1.258501e-38, 1.268018e-38, 
    1.182046e-38, 1.179782e-38, 1.171954e-38, 1.178075e-38, 1.16701e-38, 
    1.173161e-38, 1.176745e-38, 1.190806e-38, 1.193944e-38, 1.196853e-38, 
    1.202761e-38, 1.210439e-38, 1.224042e-38, 1.236223e-38, 1.247559e-38, 
    1.246725e-38, 1.247018e-38, 1.249563e-38, 1.243266e-38, 1.2506e-38, 
    1.251833e-38, 1.248608e-38, 1.267732e-38, 1.262141e-38, 1.267863e-38, 
    1.264218e-38, 1.180518e-38, 1.184352e-38, 1.18227e-38, 1.186193e-38, 
    1.183422e-38, 1.195799e-38, 1.199578e-38, 1.217791e-38, 1.210286e-38, 
    1.222263e-38, 1.211499e-38, 1.213397e-38, 1.222644e-38, 1.212079e-38, 
    1.235537e-38, 1.219509e-38, 1.249662e-38, 1.233225e-38, 1.2507e-38, 
    1.247509e-38, 1.252799e-38, 1.25757e-38, 1.263707e-38, 1.275245e-38, 
    1.272564e-38, 1.282287e-38, 1.190139e-38, 1.195196e-38, 1.194755e-38, 
    1.200128e-38, 1.204195e-38, 1.213071e-38, 1.227456e-38, 1.222026e-38, 
    1.232121e-38, 1.234187e-38, 1.218863e-38, 1.228154e-38, 1.198608e-38, 
    1.20332e-38, 1.200516e-38, 1.190534e-38, 1.223267e-38, 1.206221e-38, 
    1.238163e-38, 1.228537e-38, 1.256879e-38, 1.242683e-38, 1.271089e-38, 
    1.283676e-38, 1.295682e-38, 1.310233e-38, 1.197971e-38, 1.194523e-38, 
    1.200783e-38, 1.209649e-38, 1.217957e-38, 1.229121e-38, 1.230298e-38, 
    1.23245e-38, 1.23805e-38, 1.242779e-38, 1.233126e-38, 1.243968e-38, 
    1.204406e-38, 1.224762e-38, 1.193218e-38, 1.202507e-38, 1.209126e-38, 
    1.206223e-38, 1.221408e-38, 1.225017e-38, 1.240097e-38, 1.23224e-38, 
    1.280551e-38, 1.258586e-38, 1.321825e-38, 1.303121e-38, 1.19332e-38, 
    1.197962e-38, 1.214748e-38, 1.206725e-38, 1.22989e-38, 1.235797e-38, 
    1.240629e-38, 1.246828e-38, 1.247503e-38, 1.251196e-38, 1.245151e-38, 
    1.250959e-38, 1.229145e-38, 1.238839e-38, 1.212821e-38, 1.21903e-38, 
    1.216171e-38, 1.21304e-38, 1.222733e-38, 1.233276e-38, 1.233513e-38, 
    1.236957e-38, 1.246706e-38, 1.229987e-38, 1.283409e-38, 1.249817e-38, 
    1.203189e-38, 1.212489e-38, 1.213834e-38, 1.210216e-38, 1.235203e-38, 
    1.225972e-38, 1.251107e-38, 1.244244e-38, 1.255515e-38, 1.249899e-38, 
    1.249074e-38, 1.241911e-38, 1.237474e-38, 1.226384e-38, 1.217629e-38, 
    1.210741e-38, 1.212339e-38, 1.219919e-38, 1.233934e-38, 1.24756e-38, 
    1.244559e-38, 1.254655e-38, 1.228155e-38, 1.239182e-38, 1.234904e-38, 
    1.246097e-38, 1.22188e-38, 1.242419e-38, 1.216776e-38, 1.218972e-38, 
    1.225793e-38, 1.239928e-38, 1.243106e-38, 1.246494e-38, 1.244404e-38, 
    1.234299e-38, 1.232656e-38, 1.225628e-38, 1.223723e-38, 1.218494e-38, 
    1.214181e-38, 1.218119e-38, 1.222269e-38, 1.234307e-38, 1.245396e-38, 
    1.257638e-38, 1.260703e-38, 1.275615e-38, 1.263429e-38, 1.283599e-38, 
    1.266409e-38, 1.296348e-38, 1.243643e-38, 1.265925e-38, 1.226107e-38, 
    1.230266e-38, 1.237905e-38, 1.255655e-38, 1.246044e-38, 1.257306e-38, 
    1.232592e-38, 1.220177e-38, 1.217027e-38, 1.211157e-38, 1.217162e-38, 
    1.216672e-38, 1.222447e-38, 1.220588e-38, 1.234713e-38, 1.227029e-38, 
    1.249051e-38, 1.257218e-38, 1.281261e-38, 1.296308e-38, 1.312328e-38, 
    1.319683e-38, 1.321953e-38, 1.322904e-38,
  5.605194e-45, 5.605194e-45, 5.605194e-45, 7.006492e-45, 5.605194e-45, 
    7.006492e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  8.930465e-06, 8.770834e-06, 8.801885e-06, 8.673013e-06, 8.744523e-06, 
    8.660111e-06, 8.898124e-06, 8.764486e-06, 8.849817e-06, 8.916111e-06, 
    8.422535e-06, 8.667264e-06, 8.167904e-06, 8.324334e-06, 7.931022e-06, 
    8.192249e-06, 7.878283e-06, 7.938584e-06, 7.757048e-06, 7.809082e-06, 
    7.576555e-06, 7.733024e-06, 7.455871e-06, 7.61395e-06, 7.589228e-06, 
    7.738179e-06, 8.618066e-06, 8.453023e-06, 8.627834e-06, 8.604315e-06, 
    8.614872e-06, 8.743041e-06, 8.807571e-06, 8.942669e-06, 8.918156e-06, 
    8.818932e-06, 8.593737e-06, 8.670236e-06, 8.47739e-06, 8.481748e-06, 
    8.266713e-06, 8.363711e-06, 8.001754e-06, 8.104739e-06, 7.806912e-06, 
    7.881878e-06, 7.810431e-06, 7.832103e-06, 7.810148e-06, 7.920078e-06, 
    7.87299e-06, 7.969684e-06, 8.345548e-06, 8.235194e-06, 8.564032e-06, 
    8.761334e-06, 8.892262e-06, 8.985081e-06, 8.971962e-06, 8.946949e-06, 
    8.818351e-06, 8.697344e-06, 8.605048e-06, 8.543271e-06, 8.482375e-06, 
    8.297827e-06, 8.20008e-06, 7.98091e-06, 8.020507e-06, 7.953429e-06, 
    7.889334e-06, 7.781628e-06, 7.799365e-06, 7.751886e-06, 7.955211e-06, 
    7.820113e-06, 8.043053e-06, 7.982117e-06, 8.465756e-06, 8.649605e-06, 
    8.727621e-06, 8.795915e-06, 8.961874e-06, 8.847284e-06, 8.892467e-06, 
    8.784962e-06, 8.716599e-06, 8.750417e-06, 8.541581e-06, 8.622808e-06, 
    8.194284e-06, 8.379039e-06, 7.896812e-06, 8.012383e-06, 7.869097e-06, 
    7.942236e-06, 7.816885e-06, 7.929706e-06, 7.734217e-06, 7.6916e-06, 
    7.720723e-06, 7.608835e-06, 7.935956e-06, 7.810426e-06, 8.751362e-06, 
    8.745847e-06, 8.720156e-06, 8.833048e-06, 8.839955e-06, 8.943338e-06, 
    8.851356e-06, 8.812163e-06, 8.71264e-06, 8.653726e-06, 8.597701e-06, 
    8.474435e-06, 8.336622e-06, 8.143681e-06, 8.004894e-06, 7.911767e-06, 
    7.968883e-06, 7.918458e-06, 7.974824e-06, 8.001237e-06, 7.707566e-06, 
    7.872547e-06, 7.624934e-06, 7.638651e-06, 7.750755e-06, 7.637106e-06, 
    8.741975e-06, 8.773709e-06, 8.883811e-06, 8.797654e-06, 8.954593e-06, 
    8.866761e-06, 8.816229e-06, 8.621098e-06, 8.578202e-06, 8.538394e-06, 
    8.459752e-06, 8.358748e-06, 8.181368e-06, 8.02684e-06, 7.885607e-06, 
    7.895962e-06, 7.892316e-06, 7.860739e-06, 7.938935e-06, 7.847897e-06, 
    7.832606e-06, 7.872574e-06, 7.640488e-06, 7.706839e-06, 7.638942e-06, 
    7.682151e-06, 8.763396e-06, 8.709993e-06, 8.738852e-06, 8.684577e-06, 
    8.722812e-06, 8.552694e-06, 8.501647e-06, 8.262533e-06, 8.360735e-06, 
    8.204426e-06, 8.344869e-06, 8.319992e-06, 8.199299e-06, 8.337288e-06, 
    8.035354e-06, 8.240112e-06, 7.859511e-06, 8.064258e-06, 7.846668e-06, 
    7.886219e-06, 7.820735e-06, 7.762051e-06, 7.688194e-06, 7.551783e-06, 
    7.583387e-06, 7.469229e-06, 8.630346e-06, 8.561e-06, 8.567118e-06, 
    8.49452e-06, 8.440799e-06, 8.324302e-06, 8.137222e-06, 8.207608e-06, 
    8.078372e-06, 8.052408e-06, 8.248743e-06, 8.128221e-06, 8.514578e-06, 
    8.452223e-06, 8.489361e-06, 8.624871e-06, 8.191376e-06, 8.414022e-06, 
    8.002597e-06, 8.123441e-06, 7.770418e-06, 7.946101e-06, 7.600779e-06, 
    7.452826e-06, 7.313469e-06, 7.150341e-06, 8.52315e-06, 8.570286e-06, 
    8.485886e-06, 8.369005e-06, 8.260493e-06, 8.116072e-06, 8.101292e-06, 
    8.074211e-06, 8.004052e-06, 7.945022e-06, 8.065636e-06, 7.930221e-06, 
    8.437736e-06, 8.172037e-06, 8.588092e-06, 8.462935e-06, 8.375902e-06, 
    8.414099e-06, 8.215653e-06, 8.168832e-06, 7.978387e-06, 8.07688e-06, 
    7.489349e-06, 7.749635e-06, 7.026023e-06, 7.228675e-06, 8.586748e-06, 
    8.523318e-06, 8.302302e-06, 8.40751e-06, 8.106431e-06, 8.032206e-06, 
    7.971841e-06, 7.894613e-06, 7.886281e-06, 7.840499e-06, 7.915511e-06, 
    7.843468e-06, 8.115764e-06, 7.99416e-06, 8.327597e-06, 8.246515e-06, 
    8.283826e-06, 8.324731e-06, 8.198441e-06, 8.063736e-06, 8.060874e-06, 
    8.017646e-06, 7.895711e-06, 8.105209e-06, 7.455678e-06, 7.85719e-06, 
    8.454115e-06, 8.331762e-06, 8.314298e-06, 8.361711e-06, 8.039648e-06, 
    8.156435e-06, 7.841618e-06, 7.926787e-06, 7.787214e-06, 7.856588e-06, 
    7.866791e-06, 7.955833e-06, 8.011231e-06, 8.151079e-06, 8.264757e-06, 
    8.354838e-06, 8.333898e-06, 8.234928e-06, 8.055496e-06, 7.885518e-06, 
    7.92277e-06, 7.797827e-06, 8.128285e-06, 7.98982e-06, 8.043349e-06, 
    7.903724e-06, 8.209474e-06, 7.949104e-06, 8.275932e-06, 8.247315e-06, 
    8.158752e-06, 7.980409e-06, 7.940944e-06, 7.898757e-06, 7.924794e-06, 
    8.050941e-06, 8.071603e-06, 8.160911e-06, 8.185548e-06, 8.253548e-06, 
    8.309809e-06, 8.258402e-06, 8.204389e-06, 8.050895e-06, 7.912392e-06, 
    7.761212e-06, 7.724195e-06, 7.547219e-06, 7.691278e-06, 7.453434e-06, 
    7.655637e-06, 7.305418e-06, 7.934025e-06, 7.661616e-06, 8.154727e-06, 
    8.101704e-06, 8.005723e-06, 7.785329e-06, 7.90438e-06, 7.765148e-06, 
    8.072413e-06, 8.231503e-06, 8.272654e-06, 8.349359e-06, 8.270899e-06, 
    8.277284e-06, 8.202163e-06, 8.22631e-06, 8.045796e-06, 8.142792e-06, 
    7.867042e-06, 7.766253e-06, 7.481191e-06, 7.306096e-06, 7.127626e-06, 
    7.048739e-06, 7.02472e-06, 7.014676e-06,
  3.671203e-06, 3.539144e-06, 3.56468e-06, 3.459195e-06, 3.517571e-06, 
    3.448707e-06, 3.644294e-06, 3.53393e-06, 3.604244e-06, 3.659255e-06, 
    3.257937e-06, 3.45452e-06, 3.058637e-06, 3.180453e-06, 2.878136e-06, 
    3.077455e-06, 2.838613e-06, 2.883831e-06, 2.748687e-06, 2.787128e-06, 
    2.61721e-06, 2.731021e-06, 2.530961e-06, 2.644214e-06, 2.626349e-06, 
    2.734807e-06, 3.414624e-06, 3.282161e-06, 3.42253e-06, 3.403502e-06, 
    3.41204e-06, 3.516353e-06, 3.569355e-06, 3.681386e-06, 3.660956e-06, 
    3.578727e-06, 3.394959e-06, 3.456942e-06, 3.301603e-06, 3.305081e-06, 
    3.135347e-06, 3.211439e-06, 2.931535e-06, 3.010046e-06, 2.785519e-06, 
    2.841306e-06, 2.788126e-06, 2.80421e-06, 2.787917e-06, 2.869921e-06, 
    2.834664e-06, 2.907274e-06, 3.197129e-06, 3.110789e-06, 3.371021e-06, 
    3.531335e-06, 3.639423e-06, 3.716839e-06, 3.705858e-06, 3.684953e-06, 
    3.578247e-06, 3.479016e-06, 3.404101e-06, 3.354335e-06, 3.305581e-06, 
    3.159653e-06, 3.083524e-06, 2.915751e-06, 2.945764e-06, 2.895007e-06, 
    2.846882e-06, 2.766815e-06, 2.77993e-06, 2.744884e-06, 2.896355e-06, 
    2.795303e-06, 2.962912e-06, 2.916669e-06, 3.292298e-06, 3.440182e-06, 
    3.503724e-06, 3.559763e-06, 3.697421e-06, 3.602145e-06, 3.639592e-06, 
    3.550758e-06, 3.49473e-06, 3.522402e-06, 3.352978e-06, 3.418463e-06, 
    3.079035e-06, 3.22353e-06, 2.852478e-06, 2.939596e-06, 2.83176e-06, 
    2.886582e-06, 2.79291e-06, 2.877157e-06, 2.731894e-06, 2.700675e-06, 
    2.721991e-06, 2.640518e-06, 2.881856e-06, 2.788119e-06, 3.523175e-06, 
    3.518655e-06, 3.497637e-06, 3.590379e-06, 3.596086e-06, 3.681943e-06, 
    3.605517e-06, 3.573148e-06, 3.491499e-06, 3.443526e-06, 3.398164e-06, 
    3.299243e-06, 3.190105e-06, 3.039963e-06, 2.933915e-06, 2.863687e-06, 
    2.906672e-06, 2.868708e-06, 2.911158e-06, 2.931146e-06, 2.71235e-06, 
    2.834332e-06, 2.652172e-06, 2.66212e-06, 2.74405e-06, 2.660998e-06, 
    3.515484e-06, 3.541511e-06, 3.632407e-06, 3.5612e-06, 3.691339e-06, 
    3.618269e-06, 3.576495e-06, 3.417073e-06, 3.382437e-06, 3.350417e-06, 
    3.287543e-06, 3.207527e-06, 3.069045e-06, 2.950572e-06, 2.844095e-06, 
    2.851843e-06, 2.849114e-06, 2.825524e-06, 2.884096e-06, 2.815957e-06, 
    2.804581e-06, 2.834355e-06, 2.663453e-06, 2.711823e-06, 2.662332e-06, 
    2.69378e-06, 3.533045e-06, 3.489336e-06, 3.512928e-06, 3.468611e-06, 
    3.499804e-06, 3.361897e-06, 3.320966e-06, 3.132078e-06, 3.20909e-06, 
    3.086896e-06, 3.196598e-06, 3.177044e-06, 3.082911e-06, 3.190636e-06, 
    2.957041e-06, 3.114606e-06, 2.824609e-06, 2.979061e-06, 2.815042e-06, 
    2.844552e-06, 2.795769e-06, 2.75237e-06, 2.698191e-06, 2.599404e-06, 
    2.622142e-06, 2.540446e-06, 3.424567e-06, 3.368581e-06, 3.37351e-06, 
    3.315278e-06, 3.272463e-06, 3.180432e-06, 3.034994e-06, 3.089369e-06, 
    2.989859e-06, 2.970037e-06, 3.121341e-06, 3.028069e-06, 3.331321e-06, 
    3.281541e-06, 3.311155e-06, 3.420129e-06, 3.076786e-06, 3.251203e-06, 
    2.932173e-06, 3.024399e-06, 2.758539e-06, 2.889484e-06, 2.634693e-06, 
    2.528795e-06, 2.430911e-06, 2.318613e-06, 3.338191e-06, 3.37606e-06, 
    3.308384e-06, 3.215606e-06, 3.130495e-06, 3.018738e-06, 3.007404e-06, 
    2.986677e-06, 2.933279e-06, 2.888679e-06, 2.980122e-06, 2.877544e-06, 
    3.270009e-06, 3.061834e-06, 3.390407e-06, 3.290067e-06, 3.221053e-06, 
    3.251271e-06, 3.095612e-06, 3.059364e-06, 2.913845e-06, 2.988718e-06, 
    2.554746e-06, 2.743221e-06, 2.234738e-06, 2.372223e-06, 3.389327e-06, 
    3.338328e-06, 3.163171e-06, 3.246051e-06, 3.011343e-06, 2.954654e-06, 
    2.908906e-06, 2.85083e-06, 2.844598e-06, 2.810451e-06, 2.866496e-06, 
    2.812661e-06, 3.018502e-06, 2.925783e-06, 3.183021e-06, 3.119602e-06, 
    3.148719e-06, 3.18077e-06, 3.082265e-06, 2.97867e-06, 2.976495e-06, 
    2.943588e-06, 2.851625e-06, 3.010407e-06, 2.530802e-06, 2.822855e-06, 
    3.283056e-06, 3.186281e-06, 3.172579e-06, 3.209864e-06, 2.960317e-06, 
    3.049796e-06, 2.811284e-06, 2.874963e-06, 2.770943e-06, 2.822431e-06, 
    2.830039e-06, 2.896825e-06, 2.938722e-06, 3.045665e-06, 3.13382e-06, 
    3.204448e-06, 3.187972e-06, 3.110583e-06, 2.972386e-06, 2.844024e-06, 
    2.87194e-06, 2.778792e-06, 3.028123e-06, 2.922493e-06, 2.963131e-06, 
    2.857655e-06, 3.090814e-06, 2.891728e-06, 3.14255e-06, 3.120228e-06, 
    3.051583e-06, 2.915369e-06, 2.885609e-06, 2.853932e-06, 2.873466e-06, 
    2.968914e-06, 2.984683e-06, 3.053249e-06, 3.07228e-06, 3.125084e-06, 
    3.169062e-06, 3.128866e-06, 3.086869e-06, 2.968883e-06, 2.864151e-06, 
    2.751751e-06, 2.72454e-06, 2.596116e-06, 2.700431e-06, 2.529209e-06, 
    2.674431e-06, 2.425292e-06, 2.880389e-06, 2.678797e-06, 3.048481e-06, 
    3.00772e-06, 2.934537e-06, 2.769539e-06, 2.858148e-06, 2.754647e-06, 
    2.985303e-06, 3.107915e-06, 3.139988e-06, 3.200132e-06, 3.138619e-06, 
    3.143605e-06, 3.08515e-06, 3.103888e-06, 2.964998e-06, 3.039286e-06, 
    2.830224e-06, 2.755463e-06, 2.548948e-06, 2.425774e-06, 2.303185e-06, 
    2.249957e-06, 2.233869e-06, 2.227158e-06,
  1.690738e-06, 1.622556e-06, 1.635712e-06, 1.581455e-06, 1.611452e-06, 
    1.576073e-06, 1.676816e-06, 1.619872e-06, 1.656122e-06, 1.684555e-06, 
    1.478595e-06, 1.579056e-06, 1.377615e-06, 1.439229e-06, 1.286946e-06, 
    1.387111e-06, 1.267195e-06, 1.289795e-06, 1.222396e-06, 1.241522e-06, 
    1.157261e-06, 1.213619e-06, 1.11477e-06, 1.170603e-06, 1.161774e-06, 
    1.215499e-06, 1.5586e-06, 1.490928e-06, 1.562651e-06, 1.552904e-06, 
    1.557276e-06, 1.610826e-06, 1.638123e-06, 1.696011e-06, 1.685435e-06, 
    1.642955e-06, 1.54853e-06, 1.580299e-06, 1.500836e-06, 1.50261e-06, 
    1.416375e-06, 1.454955e-06, 1.313691e-06, 1.353132e-06, 1.240721e-06, 
    1.268539e-06, 1.242019e-06, 1.250033e-06, 1.241915e-06, 1.282838e-06, 
    1.265224e-06, 1.301531e-06, 1.44769e-06, 1.403952e-06, 1.536282e-06, 
    1.618536e-06, 1.674298e-06, 1.714383e-06, 1.70869e-06, 1.697858e-06, 
    1.642708e-06, 1.591632e-06, 1.55321e-06, 1.527753e-06, 1.502865e-06, 
    1.428685e-06, 1.390175e-06, 1.305779e-06, 1.320829e-06, 1.295389e-06, 
    1.271324e-06, 1.231411e-06, 1.237938e-06, 1.220506e-06, 1.296063e-06, 
    1.245594e-06, 1.329436e-06, 1.306239e-06, 1.496094e-06, 1.5717e-06, 
    1.604331e-06, 1.633178e-06, 1.704317e-06, 1.655039e-06, 1.674385e-06, 
    1.628538e-06, 1.599707e-06, 1.613938e-06, 1.527059e-06, 1.560567e-06, 
    1.387908e-06, 1.461097e-06, 1.274119e-06, 1.317734e-06, 1.263774e-06, 
    1.291172e-06, 1.244402e-06, 1.286456e-06, 1.214053e-06, 1.19856e-06, 
    1.209136e-06, 1.168776e-06, 1.288807e-06, 1.242016e-06, 1.614336e-06, 
    1.61201e-06, 1.601201e-06, 1.648966e-06, 1.651911e-06, 1.696299e-06, 
    1.65678e-06, 1.640078e-06, 1.598046e-06, 1.573416e-06, 1.55017e-06, 
    1.499634e-06, 1.444125e-06, 1.3682e-06, 1.314885e-06, 1.279721e-06, 
    1.30123e-06, 1.282231e-06, 1.303477e-06, 1.313496e-06, 1.204351e-06, 
    1.265058e-06, 1.174538e-06, 1.179461e-06, 1.220092e-06, 1.178906e-06, 
    1.610379e-06, 1.623775e-06, 1.670671e-06, 1.633918e-06, 1.701166e-06, 
    1.663365e-06, 1.641804e-06, 1.559855e-06, 1.542121e-06, 1.525751e-06, 
    1.49367e-06, 1.452968e-06, 1.382866e-06, 1.323242e-06, 1.269932e-06, 
    1.273802e-06, 1.272439e-06, 1.260662e-06, 1.289928e-06, 1.25589e-06, 
    1.250218e-06, 1.265069e-06, 1.18012e-06, 1.204089e-06, 1.179565e-06, 
    1.195141e-06, 1.619416e-06, 1.596935e-06, 1.609064e-06, 1.586288e-06, 
    1.602315e-06, 1.531618e-06, 1.510713e-06, 1.414721e-06, 1.453762e-06, 
    1.391878e-06, 1.44742e-06, 1.4375e-06, 1.389866e-06, 1.444395e-06, 
    1.326489e-06, 1.405882e-06, 1.260205e-06, 1.33755e-06, 1.255433e-06, 
    1.27016e-06, 1.245827e-06, 1.224227e-06, 1.197328e-06, 1.148473e-06, 
    1.159696e-06, 1.119433e-06, 1.563695e-06, 1.535035e-06, 1.537555e-06, 
    1.507811e-06, 1.485989e-06, 1.439218e-06, 1.365695e-06, 1.393127e-06, 
    1.342977e-06, 1.333015e-06, 1.409288e-06, 1.362207e-06, 1.515998e-06, 
    1.490612e-06, 1.505708e-06, 1.561421e-06, 1.386773e-06, 1.475168e-06, 
    1.314011e-06, 1.360358e-06, 1.227295e-06, 1.292624e-06, 1.165896e-06, 
    1.113706e-06, 1.065726e-06, 1.010997e-06, 1.519506e-06, 1.53886e-06, 
    1.504294e-06, 1.457072e-06, 1.41392e-06, 1.357508e-06, 1.351803e-06, 
    1.341378e-06, 1.314566e-06, 1.292221e-06, 1.338083e-06, 1.28665e-06, 
    1.48474e-06, 1.379227e-06, 1.5462e-06, 1.494957e-06, 1.459839e-06, 
    1.475202e-06, 1.396281e-06, 1.377982e-06, 1.304824e-06, 1.342404e-06, 
    1.126469e-06, 1.21968e-06, 9.703491e-07, 1.037081e-06, 1.545647e-06, 
    1.519576e-06, 1.430468e-06, 1.472547e-06, 1.353785e-06, 1.32529e-06, 
    1.302349e-06, 1.273296e-06, 1.270183e-06, 1.253144e-06, 1.281125e-06, 
    1.254246e-06, 1.357389e-06, 1.310807e-06, 1.440531e-06, 1.408409e-06, 
    1.423146e-06, 1.43939e-06, 1.389539e-06, 1.337353e-06, 1.33626e-06, 
    1.319737e-06, 1.273694e-06, 1.353314e-06, 1.114693e-06, 1.25933e-06, 
    1.491384e-06, 1.442185e-06, 1.435236e-06, 1.454155e-06, 1.328134e-06, 
    1.373156e-06, 1.253559e-06, 1.285359e-06, 1.233465e-06, 1.259119e-06, 
    1.262915e-06, 1.296299e-06, 1.317296e-06, 1.371074e-06, 1.415603e-06, 
    1.451405e-06, 1.443043e-06, 1.403848e-06, 1.334195e-06, 1.269897e-06, 
    1.283847e-06, 1.237372e-06, 1.362234e-06, 1.309158e-06, 1.329547e-06, 
    1.276706e-06, 1.393857e-06, 1.293747e-06, 1.420022e-06, 1.408725e-06, 
    1.374057e-06, 1.305587e-06, 1.290685e-06, 1.274846e-06, 1.28461e-06, 
    1.332451e-06, 1.340375e-06, 1.374898e-06, 1.384499e-06, 1.411182e-06, 
    1.433453e-06, 1.413095e-06, 1.391865e-06, 1.332436e-06, 1.279953e-06, 
    1.22392e-06, 1.210401e-06, 1.146851e-06, 1.198439e-06, 1.11391e-06, 
    1.185555e-06, 1.062979e-06, 1.288073e-06, 1.187718e-06, 1.372493e-06, 
    1.351962e-06, 1.315197e-06, 1.232767e-06, 1.276952e-06, 1.225359e-06, 
    1.340687e-06, 1.402499e-06, 1.418725e-06, 1.449214e-06, 1.418032e-06, 
    1.420556e-06, 1.390996e-06, 1.400463e-06, 1.330484e-06, 1.367858e-06, 
    1.263007e-06, 1.225765e-06, 1.123616e-06, 1.063215e-06, 1.003506e-06, 
    9.777102e-07, 9.699291e-07, 9.666854e-07,
  4.260761e-07, 4.054311e-07, 4.093989e-07, 3.930841e-07, 4.020879e-07, 
    3.914729e-07, 4.218442e-07, 4.046224e-07, 4.155693e-07, 4.241953e-07, 
    3.62517e-07, 3.923656e-07, 3.329851e-07, 3.509467e-07, 3.068893e-07, 
    3.357416e-07, 3.012593e-07, 3.077029e-07, 2.885635e-07, 2.939711e-07, 
    2.702913e-07, 2.860882e-07, 2.584937e-07, 2.740157e-07, 2.715501e-07, 
    2.866182e-07, 3.862507e-07, 3.661568e-07, 3.874602e-07, 3.845513e-07, 
    3.858557e-07, 4.018996e-07, 4.101268e-07, 4.276807e-07, 4.244629e-07, 
    4.115865e-07, 3.832475e-07, 3.927377e-07, 3.690852e-07, 3.696099e-07, 
    3.442632e-07, 3.5556e-07, 3.145439e-07, 3.258983e-07, 2.937442e-07, 
    3.016418e-07, 2.941119e-07, 2.963834e-07, 2.940824e-07, 3.057165e-07, 
    3.006984e-07, 3.110592e-07, 3.534273e-07, 3.406406e-07, 3.796008e-07, 
    4.042204e-07, 4.210795e-07, 4.332821e-07, 4.315447e-07, 4.282434e-07, 
    4.115118e-07, 3.961343e-07, 3.846426e-07, 3.77065e-07, 3.696854e-07, 
    3.478605e-07, 3.366319e-07, 3.122756e-07, 3.16593e-07, 3.093018e-07, 
    3.024345e-07, 2.9111e-07, 2.929563e-07, 2.880303e-07, 3.094946e-07, 
    2.951249e-07, 3.190675e-07, 3.124073e-07, 3.676833e-07, 3.901646e-07, 
    3.999471e-07, 4.08634e-07, 4.302115e-07, 4.152415e-07, 4.211061e-07, 
    4.072342e-07, 3.985577e-07, 4.028358e-07, 3.768591e-07, 3.868378e-07, 
    3.359732e-07, 3.57365e-07, 3.032307e-07, 3.157042e-07, 3.002861e-07, 
    3.080962e-07, 2.94787e-07, 3.067492e-07, 2.862106e-07, 2.818509e-07, 
    2.848255e-07, 2.73505e-07, 3.074205e-07, 2.94111e-07, 4.029555e-07, 
    4.022558e-07, 3.990065e-07, 4.134038e-07, 4.142948e-07, 4.277685e-07, 
    4.157685e-07, 4.107172e-07, 3.980589e-07, 3.906777e-07, 3.837362e-07, 
    3.687295e-07, 3.523819e-07, 3.302563e-07, 3.148864e-07, 3.048274e-07, 
    3.109728e-07, 3.055433e-07, 3.116163e-07, 3.144878e-07, 2.834791e-07, 
    3.006513e-07, 2.751161e-07, 2.764936e-07, 2.879134e-07, 2.763382e-07, 
    4.017651e-07, 4.057982e-07, 4.199788e-07, 4.088573e-07, 4.29251e-07, 
    4.177636e-07, 4.112389e-07, 3.866253e-07, 3.813383e-07, 3.764705e-07, 
    3.669664e-07, 3.549765e-07, 3.345087e-07, 3.172863e-07, 3.020382e-07, 
    3.031404e-07, 3.02752e-07, 2.994014e-07, 3.077407e-07, 2.980456e-07, 
    2.964359e-07, 3.006545e-07, 2.766783e-07, 2.834053e-07, 2.765229e-07, 
    2.808905e-07, 4.04485e-07, 3.977253e-07, 4.013696e-07, 3.945321e-07, 
    3.993412e-07, 3.782138e-07, 3.720099e-07, 3.437806e-07, 3.552097e-07, 
    3.371269e-07, 3.533482e-07, 3.504403e-07, 3.365422e-07, 3.524607e-07, 
    3.182199e-07, 3.412031e-07, 2.992717e-07, 3.214035e-07, 2.979161e-07, 
    3.021032e-07, 2.951907e-07, 2.890805e-07, 2.815048e-07, 2.678431e-07, 
    2.709702e-07, 2.597836e-07, 3.877719e-07, 3.792296e-07, 3.799793e-07, 
    3.711499e-07, 3.646977e-07, 3.509435e-07, 3.295312e-07, 3.374899e-07, 
    3.229675e-07, 3.200973e-07, 3.421956e-07, 3.285217e-07, 3.735763e-07, 
    3.660631e-07, 3.705271e-07, 3.870928e-07, 3.356433e-07, 3.615066e-07, 
    3.146357e-07, 3.279869e-07, 2.899467e-07, 3.085114e-07, 2.727008e-07, 
    2.581995e-07, 2.449997e-07, 2.301029e-07, 3.746166e-07, 3.803674e-07, 
    3.701085e-07, 3.56182e-07, 3.435466e-07, 3.271627e-07, 3.255143e-07, 
    3.225063e-07, 3.147947e-07, 3.08396e-07, 3.215569e-07, 3.068045e-07, 
    3.643295e-07, 3.334527e-07, 3.825531e-07, 3.673468e-07, 3.569951e-07, 
    3.615166e-07, 3.384072e-07, 3.330912e-07, 3.12002e-07, 3.228022e-07, 
    2.617322e-07, 2.877973e-07, 2.191509e-07, 2.371815e-07, 3.823883e-07, 
    3.746373e-07, 3.483816e-07, 3.607343e-07, 3.260869e-07, 3.178752e-07, 
    3.112931e-07, 3.029962e-07, 3.021098e-07, 2.972662e-07, 3.052278e-07, 
    2.975789e-07, 3.271284e-07, 3.137166e-07, 3.513282e-07, 3.419393e-07, 
    3.462405e-07, 3.509937e-07, 3.364468e-07, 3.213467e-07, 3.210316e-07, 
    3.162794e-07, 3.031101e-07, 3.259508e-07, 2.584727e-07, 2.990236e-07, 
    3.662909e-07, 3.518132e-07, 3.497772e-07, 3.553249e-07, 3.186927e-07, 
    3.316921e-07, 2.973841e-07, 3.06436e-07, 2.916907e-07, 2.989629e-07, 
    3.000418e-07, 3.095618e-07, 3.155784e-07, 3.310887e-07, 3.440377e-07, 
    3.545175e-07, 3.520644e-07, 3.406101e-07, 3.204372e-07, 3.020283e-07, 
    3.060046e-07, 2.92796e-07, 3.285294e-07, 3.132439e-07, 3.190993e-07, 
    3.039679e-07, 3.377022e-07, 3.088329e-07, 3.453279e-07, 3.420315e-07, 
    3.319533e-07, 3.122209e-07, 3.07957e-07, 3.034378e-07, 3.062222e-07, 
    3.199351e-07, 3.222174e-07, 3.321969e-07, 3.349827e-07, 3.427478e-07, 
    3.492551e-07, 3.43306e-07, 3.371228e-07, 3.199305e-07, 3.048936e-07, 
    2.889936e-07, 2.851818e-07, 2.673921e-07, 2.818171e-07, 2.582563e-07, 
    2.782017e-07, 2.442484e-07, 3.072113e-07, 2.788076e-07, 3.315e-07, 
    3.255603e-07, 3.149761e-07, 2.914935e-07, 3.04038e-07, 2.894002e-07, 
    3.223072e-07, 3.402174e-07, 3.449491e-07, 3.538745e-07, 3.447467e-07, 
    3.454839e-07, 3.368704e-07, 3.396244e-07, 3.19369e-07, 3.301572e-07, 
    3.000682e-07, 2.895148e-07, 2.609415e-07, 2.443127e-07, 2.280769e-07, 
    2.211268e-07, 2.190382e-07, 2.181685e-07,
  3.882819e-08, 3.648678e-08, 3.693427e-08, 3.510205e-08, 3.611067e-08, 
    3.492222e-08, 3.83456e-08, 3.639573e-08, 3.763255e-08, 3.861354e-08, 
    3.17257e-08, 3.502183e-08, 2.853646e-08, 3.046742e-08, 2.5781e-08, 
    2.883103e-08, 2.519453e-08, 2.586596e-08, 2.388276e-08, 2.443964e-08, 
    2.20217e-08, 2.362877e-08, 2.083738e-08, 2.239841e-08, 2.214886e-08, 
    2.368311e-08, 3.434075e-08, 3.21238e-08, 3.447524e-08, 3.415202e-08, 
    3.429686e-08, 3.608951e-08, 3.701652e-08, 3.90115e-08, 3.864406e-08, 
    3.718151e-08, 3.400736e-08, 3.506335e-08, 3.244481e-08, 3.250241e-08, 
    2.97457e-08, 3.096776e-08, 2.658294e-08, 2.778219e-08, 2.441623e-08, 
    2.523426e-08, 2.445418e-08, 2.468895e-08, 2.445114e-08, 2.565857e-08, 
    2.513625e-08, 2.621719e-08, 3.073624e-08, 2.93561e-08, 3.360347e-08, 
    3.635051e-08, 3.825856e-08, 3.965295e-08, 3.945375e-08, 3.907584e-08, 
    3.717306e-08, 3.544302e-08, 3.416213e-08, 3.332325e-08, 3.251069e-08, 
    3.013373e-08, 2.892629e-08, 2.634476e-08, 2.679852e-08, 2.603316e-08, 
    2.531669e-08, 2.414466e-08, 2.433494e-08, 2.382801e-08, 2.605333e-08, 
    2.455883e-08, 2.705934e-08, 2.635855e-08, 3.229109e-08, 3.477633e-08, 
    3.587031e-08, 3.684791e-08, 3.930104e-08, 3.759538e-08, 3.826158e-08, 
    3.668996e-08, 3.571444e-08, 3.619472e-08, 3.330051e-08, 3.440602e-08, 
    2.885579e-08, 3.116402e-08, 2.539954e-08, 2.670497e-08, 2.509343e-08, 
    2.590706e-08, 2.452391e-08, 2.576634e-08, 2.364132e-08, 2.319534e-08, 
    2.349944e-08, 2.234666e-08, 2.583645e-08, 2.44541e-08, 3.620818e-08, 
    3.612953e-08, 3.576476e-08, 3.738717e-08, 3.748809e-08, 3.902154e-08, 
    3.765513e-08, 3.708321e-08, 3.565853e-08, 3.483352e-08, 3.406156e-08, 
    3.240577e-08, 3.06229e-08, 2.824551e-08, 2.661895e-08, 2.556584e-08, 
    2.620814e-08, 2.56405e-08, 2.627559e-08, 2.657704e-08, 2.336169e-08, 
    2.513136e-08, 2.250996e-08, 2.264979e-08, 2.381601e-08, 2.2634e-08, 
    3.607439e-08, 3.652812e-08, 3.813333e-08, 3.68731e-08, 3.919109e-08, 
    3.788157e-08, 3.71422e-08, 3.438241e-08, 3.379577e-08, 3.325763e-08, 
    3.221242e-08, 3.090438e-08, 2.869918e-08, 2.687155e-08, 2.527547e-08, 
    2.539013e-08, 2.534972e-08, 2.500162e-08, 2.586991e-08, 2.486105e-08, 
    2.469439e-08, 2.513168e-08, 2.266855e-08, 2.335414e-08, 2.265276e-08, 
    2.309732e-08, 3.638023e-08, 3.562116e-08, 3.602996e-08, 3.526382e-08, 
    3.58023e-08, 3.345016e-08, 3.276619e-08, 2.969375e-08, 3.092971e-08, 
    2.897928e-08, 3.072764e-08, 3.04126e-08, 2.89167e-08, 3.063141e-08, 
    2.696997e-08, 2.941655e-08, 2.498816e-08, 2.730612e-08, 2.484763e-08, 
    2.528223e-08, 2.456562e-08, 2.393589e-08, 2.316e-08, 2.177478e-08, 
    2.209025e-08, 2.096619e-08, 3.450991e-08, 3.356243e-08, 3.364533e-08, 
    3.26716e-08, 3.196402e-08, 3.046706e-08, 2.81683e-08, 2.901814e-08, 
    2.747155e-08, 2.716807e-08, 2.952318e-08, 2.806091e-08, 3.293858e-08, 
    3.211349e-08, 3.260316e-08, 3.443438e-08, 2.882049e-08, 3.161534e-08, 
    2.659259e-08, 2.800403e-08, 2.402495e-08, 2.595049e-08, 2.226524e-08, 
    2.080805e-08, 1.950004e-08, 1.804579e-08, 3.305318e-08, 3.368828e-08, 
    3.255716e-08, 3.103537e-08, 2.966854e-08, 2.791645e-08, 2.774144e-08, 
    2.742274e-08, 2.66093e-08, 2.593841e-08, 2.732233e-08, 2.577211e-08, 
    3.192379e-08, 2.858637e-08, 3.393037e-08, 3.225415e-08, 3.112377e-08, 
    3.161641e-08, 2.911644e-08, 2.854776e-08, 2.631605e-08, 2.745404e-08, 
    2.116112e-08, 2.38041e-08, 1.699192e-08, 1.873387e-08, 3.391209e-08, 
    3.305545e-08, 3.018999e-08, 3.153106e-08, 2.780221e-08, 2.693361e-08, 
    2.624171e-08, 2.537513e-08, 2.528292e-08, 2.478032e-08, 2.560759e-08, 
    2.481271e-08, 2.79128e-08, 2.649601e-08, 3.050872e-08, 2.949563e-08, 
    2.995882e-08, 3.04725e-08, 2.890645e-08, 2.730011e-08, 2.726677e-08, 
    2.676551e-08, 2.538705e-08, 2.778776e-08, 2.083534e-08, 2.496249e-08, 
    3.213842e-08, 3.056127e-08, 3.034085e-08, 3.094221e-08, 2.701981e-08, 
    2.83985e-08, 2.479253e-08, 2.573364e-08, 2.420447e-08, 2.495613e-08, 
    2.506807e-08, 2.606037e-08, 2.669173e-08, 2.833418e-08, 2.972142e-08, 
    3.085453e-08, 3.058846e-08, 2.935282e-08, 2.720398e-08, 2.527445e-08, 
    2.568864e-08, 2.43184e-08, 2.806171e-08, 2.644638e-08, 2.706272e-08, 
    2.547629e-08, 2.90409e-08, 2.598416e-08, 2.98604e-08, 2.950554e-08, 
    2.842635e-08, 2.633903e-08, 2.589251e-08, 2.54211e-08, 2.571133e-08, 
    2.715095e-08, 2.739217e-08, 2.845233e-08, 2.874983e-08, 2.958257e-08, 
    3.028438e-08, 2.964264e-08, 2.897884e-08, 2.715046e-08, 2.557277e-08, 
    2.392697e-08, 2.353591e-08, 2.172939e-08, 2.319191e-08, 2.081375e-08, 
    2.28235e-08, 1.942618e-08, 2.581464e-08, 2.288512e-08, 2.837801e-08, 
    2.774632e-08, 2.66284e-08, 2.418419e-08, 2.54836e-08, 2.396877e-08, 
    2.740167e-08, 2.931066e-08, 2.981959e-08, 3.078474e-08, 2.979777e-08, 
    2.987723e-08, 2.895179e-08, 2.9247e-08, 2.709117e-08, 2.823494e-08, 
    2.507081e-08, 2.398054e-08, 2.108196e-08, 1.943247e-08, 1.784984e-08, 
    1.718108e-08, 1.698114e-08, 1.689804e-08,
  1.121087e-09, 1.036321e-09, 1.052411e-09, 9.86869e-10, 1.022838e-09, 
    9.804847e-10, 1.1035e-09, 1.033054e-09, 1.077623e-09, 1.113256e-09, 
    8.68511e-10, 9.8402e-10, 7.597664e-10, 8.252387e-10, 6.68384e-10, 
    7.696802e-10, 6.492592e-10, 6.711638e-10, 6.069127e-10, 6.248161e-10, 
    5.478942e-10, 5.987836e-10, 5.110126e-10, 5.597372e-10, 5.518858e-10, 
    6.005207e-10, 9.599024e-10, 8.822982e-10, 9.646545e-10, 9.532419e-10, 
    9.583526e-10, 1.022081e-09, 1.055375e-09, 1.127782e-09, 1.114369e-09, 
    1.061323e-09, 9.481438e-10, 9.854937e-10, 8.934464e-10, 8.954505e-10, 
    8.006337e-10, 8.423883e-10, 6.947226e-10, 7.345064e-10, 6.24061e-10, 
    6.505508e-10, 6.252852e-10, 6.328665e-10, 6.251868e-10, 6.643815e-10, 
    6.473647e-10, 6.826833e-10, 8.344435e-10, 7.874172e-10, 9.339397e-10, 
    1.031433e-09, 1.100334e-09, 1.151279e-09, 1.143971e-09, 1.130135e-09, 
    1.061019e-09, 9.989972e-10, 9.535981e-10, 9.241111e-10, 8.957388e-10, 
    8.138439e-10, 7.728915e-10, 6.868777e-10, 7.018394e-10, 6.766427e-10, 
    6.532327e-10, 6.153192e-10, 6.214416e-10, 6.051585e-10, 6.773038e-10, 
    6.286625e-10, 7.104705e-10, 6.873311e-10, 8.881056e-10, 9.753116e-10, 
    1.014243e-09, 1.049302e-09, 1.138376e-09, 1.076278e-09, 1.100444e-09, 
    1.04362e-09, 1.008675e-09, 1.025847e-09, 9.233146e-10, 9.622078e-10, 
    7.705144e-10, 8.491362e-10, 6.559308e-10, 6.987491e-10, 6.459737e-10, 
    6.725094e-10, 6.275351e-10, 6.679041e-10, 5.991846e-10, 5.849655e-10, 
    5.946535e-10, 5.581068e-10, 6.701978e-10, 6.252827e-10, 1.02633e-09, 
    1.023513e-09, 1.010471e-09, 1.068749e-09, 1.072397e-09, 1.128149e-09, 
    1.078441e-09, 1.057778e-09, 1.00668e-09, 9.773387e-10, 9.500528e-10, 
    8.920891e-10, 8.305601e-10, 7.500012e-10, 6.959102e-10, 6.613536e-10, 
    6.823856e-10, 6.637911e-10, 6.846024e-10, 6.945278e-10, 5.90261e-10, 
    6.47206e-10, 5.632542e-10, 5.676693e-10, 6.047742e-10, 5.671705e-10, 
    1.021539e-09, 1.037804e-09, 1.095783e-09, 1.050208e-09, 1.13435e-09, 
    1.086645e-09, 1.059905e-09, 9.613743e-10, 9.406963e-10, 9.218132e-10, 
    8.853714e-10, 8.402117e-10, 7.652389e-10, 7.042543e-10, 6.518913e-10, 
    6.556241e-10, 6.543079e-10, 6.429938e-10, 6.712931e-10, 6.384367e-10, 
    6.330427e-10, 6.472162e-10, 5.682625e-10, 5.900199e-10, 5.677634e-10, 
    5.818497e-10, 1.032497e-09, 1.005347e-09, 1.019949e-09, 9.926191e-10, 
    1.011812e-09, 9.285602e-10, 9.046408e-10, 7.988691e-10, 8.410816e-10, 
    7.746789e-10, 8.341486e-10, 8.233644e-10, 7.725689e-10, 8.308512e-10, 
    7.075112e-10, 7.894655e-10, 6.425571e-10, 7.186585e-10, 6.380019e-10, 
    6.521111e-10, 6.288812e-10, 6.08616e-10, 5.838415e-10, 5.4016e-10, 
    5.500448e-10, 5.149972e-10, 9.658802e-10, 9.32499e-10, 9.354091e-10, 
    9.013423e-10, 8.767572e-10, 8.25226e-10, 7.474141e-10, 7.759903e-10, 
    7.241564e-10, 7.14075e-10, 7.93079e-10, 7.438195e-10, 9.106563e-10, 
    8.819394e-10, 8.989582e-10, 9.632104e-10, 7.693245e-10, 8.64696e-10, 
    6.95041e-10, 7.419169e-10, 6.114738e-10, 6.739329e-10, 5.555442e-10, 
    5.101064e-10, 4.700292e-10, 4.263013e-10, 9.146604e-10, 9.369179e-10, 
    8.973563e-10, 8.44712e-10, 7.980122e-10, 7.389895e-10, 7.33147e-10, 
    7.225331e-10, 6.95592e-10, 6.735363e-10, 7.191961e-10, 6.680927e-10, 
    8.753654e-10, 7.614439e-10, 9.454322e-10, 8.86821e-10, 8.477514e-10, 
    8.647324e-10, 7.793101e-10, 7.601454e-10, 6.859333e-10, 7.23574e-10, 
    5.210408e-10, 6.043934e-10, 3.951837e-10, 4.468799e-10, 9.447886e-10, 
    9.147396e-10, 8.15762e-10, 8.61785e-10, 7.351745e-10, 7.06307e-10, 
    6.834887e-10, 6.55136e-10, 6.521335e-10, 6.358228e-10, 6.627164e-10, 
    6.368709e-10, 7.388675e-10, 6.918571e-10, 8.266509e-10, 7.921451e-10, 
    8.078824e-10, 8.254119e-10, 7.722216e-10, 7.184581e-10, 7.173506e-10, 
    7.00749e-10, 6.555261e-10, 7.346924e-10, 5.109507e-10, 6.417262e-10, 
    8.828029e-10, 8.284506e-10, 8.209121e-10, 8.415107e-10, 7.091612e-10, 
    7.551323e-10, 6.362177e-10, 6.668348e-10, 6.172421e-10, 6.415183e-10, 
    6.451503e-10, 6.775345e-10, 6.983122e-10, 7.529743e-10, 7.998085e-10, 
    8.385004e-10, 8.293802e-10, 7.873062e-10, 7.152668e-10, 6.518582e-10, 
    6.653642e-10, 6.209088e-10, 7.438459e-10, 6.902224e-10, 7.105828e-10, 
    6.584324e-10, 7.767587e-10, 6.750375e-10, 8.045331e-10, 7.924809e-10, 
    7.560674e-10, 6.866893e-10, 6.72033e-10, 6.566334e-10, 6.661053e-10, 
    7.135077e-10, 7.215168e-10, 7.569393e-10, 7.669441e-10, 7.950938e-10, 
    8.189832e-10, 7.971327e-10, 7.746641e-10, 7.13491e-10, 6.615798e-10, 
    6.083301e-10, 5.958173e-10, 5.387417e-10, 5.848571e-10, 5.102836e-10, 
    5.731669e-10, 4.677879e-10, 6.69485e-10, 5.75118e-10, 7.544445e-10, 
    7.333096e-10, 6.962224e-10, 6.165904e-10, 6.586707e-10, 6.096711e-10, 
    7.218326e-10, 7.858793e-10, 8.03145e-10, 8.361064e-10, 8.024031e-10, 
    8.051055e-10, 7.737508e-10, 7.837241e-10, 7.115253e-10, 7.496465e-10, 
    6.452395e-10, 6.100488e-10, 5.185847e-10, 4.679782e-10, 4.204776e-10, 
    4.007321e-10, 3.948678e-10, 3.924357e-10,
  9.033904e-12, 8.13938e-12, 8.307563e-12, 7.62736e-12, 7.999038e-12, 
    7.561804e-12, 8.846605e-12, 8.10533e-12, 8.572637e-12, 8.9504e-12, 
    6.433369e-12, 7.598089e-12, 5.378786e-12, 6.008593e-12, 4.527471e-12, 
    5.473127e-12, 4.353667e-12, 4.552858e-12, 3.974536e-12, 4.133847e-12, 
    3.459982e-12, 3.902684e-12, 3.147137e-12, 3.561889e-12, 3.49425e-12, 
    3.918013e-12, 7.351326e-12, 6.57007e-12, 7.399802e-12, 7.283506e-12, 
    7.335531e-12, 7.99118e-12, 8.338638e-12, 9.105425e-12, 8.962255e-12, 
    8.40106e-12, 7.231689e-12, 7.613222e-12, 6.681055e-12, 6.701056e-12, 
    5.770048e-12, 6.176144e-12, 4.769359e-12, 5.14012e-12, 4.127099e-12, 
    4.365351e-12, 4.138041e-12, 4.205953e-12, 4.137162e-12, 4.490963e-12, 
    4.336533e-12, 4.65843e-12, 6.098393e-12, 5.64283e-12, 7.087756e-12, 
    8.088451e-12, 8.812988e-12, 9.357449e-12, 9.278904e-12, 9.130593e-12, 
    8.397859e-12, 7.752238e-12, 7.287125e-12, 6.988542e-12, 6.703934e-12, 
    5.897859e-12, 5.503762e-12, 4.697012e-12, 4.835213e-12, 4.603004e-12, 
    4.389644e-12, 4.049161e-12, 4.10371e-12, 3.959007e-12, 4.609059e-12, 
    4.168265e-12, 4.915355e-12, 4.701184e-12, 6.627845e-12, 7.508774e-12, 
    7.909872e-12, 8.275008e-12, 9.218861e-12, 8.558455e-12, 8.814158e-12, 
    8.215574e-12, 7.852214e-12, 8.030315e-12, 6.980516e-12, 7.374833e-12, 
    5.481079e-12, 6.242358e-12, 4.414115e-12, 4.806592e-12, 4.323964e-12, 
    4.56516e-12, 4.15817e-12, 4.523084e-12, 3.906223e-12, 3.781254e-12, 
    3.866297e-12, 3.547815e-12, 4.54403e-12, 4.13802e-12, 8.035333e-12, 
    8.006053e-12, 7.870798e-12, 8.479131e-12, 8.517541e-12, 9.109355e-12, 
    8.581262e-12, 8.363838e-12, 7.831577e-12, 7.529541e-12, 7.251079e-12, 
    6.667521e-12, 6.060474e-12, 5.286227e-12, 4.780334e-12, 4.463392e-12, 
    4.655694e-12, 4.485582e-12, 4.676072e-12, 4.767557e-12, 3.827685e-12, 
    4.335099e-12, 3.592283e-12, 3.630527e-12, 3.955608e-12, 3.626202e-12, 
    7.98555e-12, 8.154851e-12, 8.764702e-12, 8.284492e-12, 9.175722e-12, 
    8.667941e-12, 8.386172e-12, 7.366338e-12, 7.156136e-12, 6.965394e-12, 
    6.600609e-12, 6.154821e-12, 5.430812e-12, 4.857608e-12, 4.377489e-12, 
    4.41133e-12, 4.399391e-12, 4.297068e-12, 4.554039e-12, 4.256013e-12, 
    4.207536e-12, 4.33519e-12, 3.635672e-12, 3.825566e-12, 3.631343e-12, 
    3.753994e-12, 8.09952e-12, 7.8178e-12, 7.969043e-12, 7.686508e-12, 
    7.884684e-12, 7.033421e-12, 6.792953e-12, 5.75303e-12, 6.163342e-12, 
    5.52083e-12, 6.095511e-12, 5.990345e-12, 5.500689e-12, 6.063309e-12, 
    4.88785e-12, 5.66251e-12, 4.29313e-12, 4.991675e-12, 4.2521e-12, 
    4.37948e-12, 4.170221e-12, 3.989632e-12, 3.771414e-12, 3.393801e-12, 
    3.478432e-12, 3.180596e-12, 7.412316e-12, 7.073194e-12, 7.102612e-12, 
    6.759932e-12, 6.515034e-12, 6.008467e-12, 5.261766e-12, 5.533358e-12, 
    5.043053e-12, 4.948917e-12, 5.697246e-12, 5.227826e-12, 6.853246e-12, 
    6.56649e-12, 6.736097e-12, 7.385065e-12, 5.469732e-12, 6.395645e-12, 
    4.772301e-12, 5.209879e-12, 4.014986e-12, 4.578189e-12, 3.525727e-12, 
    3.139543e-12, 2.807922e-12, 2.456452e-12, 6.893446e-12, 7.117877e-12, 
    6.720088e-12, 6.198932e-12, 5.744762e-12, 5.182297e-12, 5.127346e-12, 
    5.027869e-12, 4.777391e-12, 4.574555e-12, 4.99669e-12, 4.524805e-12, 
    6.501246e-12, 5.39472e-12, 7.20416e-12, 6.615043e-12, 6.228758e-12, 
    6.396e-12, 5.565109e-12, 5.382379e-12, 4.688318e-12, 5.037603e-12, 
    3.231512e-12, 3.952241e-12, 2.213373e-12, 2.620462e-12, 7.197627e-12, 
    6.89424e-12, 5.916458e-12, 6.366899e-12, 5.1464e-12, 4.87666e-12, 
    4.665831e-12, 4.406904e-12, 4.379684e-12, 4.232505e-12, 4.475795e-12, 
    4.241927e-12, 5.181148e-12, 4.742902e-12, 6.022347e-12, 5.688264e-12, 
    5.840092e-12, 6.010277e-12, 5.497361e-12, 4.989799e-12, 4.979458e-12, 
    4.825112e-12, 4.41046e-12, 5.141868e-12, 3.14663e-12, 4.285654e-12, 
    6.575066e-12, 6.039899e-12, 5.966486e-12, 6.167543e-12, 4.903181e-12, 
    5.334812e-12, 4.236054e-12, 4.513328e-12, 4.066274e-12, 4.283765e-12, 
    4.316528e-12, 4.611174e-12, 4.802549e-12, 5.314366e-12, 5.762086e-12, 
    6.138065e-12, 6.048956e-12, 5.641764e-12, 4.960028e-12, 4.377192e-12, 
    4.49992e-12, 4.098955e-12, 5.228072e-12, 4.727827e-12, 4.916405e-12, 
    4.436832e-12, 5.540705e-12, 4.588312e-12, 5.807703e-12, 5.691491e-12, 
    5.343677e-12, 4.69528e-12, 4.560803e-12, 4.420494e-12, 4.506674e-12, 
    4.943634e-12, 5.018368e-12, 5.351945e-12, 5.447046e-12, 5.71664e-12, 
    5.947735e-12, 5.736284e-12, 5.520687e-12, 4.943476e-12, 4.465452e-12, 
    3.987098e-12, 3.876541e-12, 3.381705e-12, 3.78031e-12, 3.141038e-12, 
    3.678299e-12, 2.789649e-12, 4.537528e-12, 3.695272e-12, 5.328291e-12, 
    5.128874e-12, 4.783225e-12, 4.060478e-12, 4.438996e-12, 3.998992e-12, 
    5.02132e-12, 5.62807e-12, 5.794291e-12, 6.114647e-12, 5.787126e-12, 
    5.813235e-12, 5.51196e-12, 5.607392e-12, 4.925173e-12, 5.282868e-12, 
    4.317335e-12, 4.002341e-12, 3.210795e-12, 2.791193e-12, 2.410496e-12, 
    2.256265e-12, 2.210935e-12, 2.192201e-12,
  1.140901e-14, 9.431197e-15, 9.794042e-15, 8.353593e-15, 9.13172e-15, 
    8.218653e-15, 1.09853e-14, 9.358269e-15, 1.037454e-14, 1.121948e-14, 
    6.011736e-15, 8.293255e-15, 4.168972e-15, 5.241947e-15, 2.862697e-15, 
    4.324242e-15, 2.618482e-15, 2.899029e-15, 2.114732e-15, 2.321429e-15, 
    1.499738e-15, 2.023944e-15, 1.168206e-15, 1.614872e-15, 1.538072e-15, 
    2.043185e-15, 7.79019e-15, 6.266885e-15, 7.888215e-15, 7.653726e-15, 
    7.758338e-15, 9.11505e-15, 9.861578e-15, 1.157207e-14, 1.124633e-14, 
    9.997613e-15, 7.549984e-15, 8.324417e-15, 6.476551e-15, 6.514586e-15, 
    4.825609e-15, 5.541311e-15, 3.215735e-15, 3.785183e-15, 2.312525e-15, 
    2.634635e-15, 2.326971e-15, 2.417377e-15, 2.325809e-15, 2.81072e-15, 
    2.59484e-15, 3.051962e-15, 5.401695e-15, 4.608459e-15, 7.264227e-15, 
    9.322202e-15, 1.090978e-14, 1.215234e-14, 1.197057e-14, 1.162964e-14, 
    9.990622e-15, 8.61256e-15, 7.660973e-15, 7.069346e-15, 6.520067e-15, 
    5.047244e-15, 4.375079e-15, 3.108576e-15, 3.314424e-15, 2.971316e-15, 
    2.668357e-15, 2.210638e-15, 2.281766e-15, 2.094984e-15, 2.980082e-15, 
    2.36705e-15, 3.435975e-15, 3.114711e-15, 6.37578e-15, 8.109997e-15, 
    8.943081e-15, 9.723477e-15, 1.183218e-14, 1.034323e-14, 1.091241e-14, 
    9.595038e-15, 8.821703e-15, 9.19819e-15, 7.053659e-15, 7.83767e-15, 
    4.337412e-15, 5.66117e-15, 2.70249e-15, 3.271399e-15, 2.577551e-15, 
    2.916697e-15, 2.353635e-15, 2.856419e-15, 2.028381e-15, 1.874052e-15, 
    1.978561e-15, 1.598763e-15, 2.886369e-15, 2.326947e-15, 9.208874e-15, 
    9.146615e-15, 8.860752e-15, 1.016859e-14, 1.025303e-14, 1.158106e-14, 
    1.03936e-14, 9.916411e-15, 8.778397e-15, 8.152489e-15, 7.58874e-15, 
    6.450859e-15, 5.334048e-15, 4.01858e-15, 3.232106e-15, 2.771705e-15, 
    3.047958e-15, 2.803087e-15, 3.077795e-15, 3.213045e-15, 1.930839e-15, 
    2.592868e-15, 1.649865e-15, 1.694322e-15, 2.090671e-15, 1.68927e-15, 
    9.103097e-15, 9.46438e-15, 1.080158e-14, 9.744004e-15, 1.173305e-14, 
    1.058578e-14, 9.965118e-15, 7.820515e-15, 7.399526e-15, 7.024136e-15, 
    6.32431e-15, 5.502901e-15, 4.254338e-15, 3.348238e-15, 2.651462e-15, 
    2.698594e-15, 2.68193e-15, 2.540708e-15, 2.900723e-15, 2.484851e-15, 
    2.419505e-15, 2.592989e-15, 1.700339e-15, 1.928227e-15, 1.695276e-15, 
    1.841016e-15, 9.345817e-15, 8.749532e-15, 9.068109e-15, 8.475934e-15, 
    8.889978e-15, 7.157301e-15, 6.690323e-15, 4.796374e-15, 5.518242e-15, 
    4.403489e-15, 5.396538e-15, 5.209684e-15, 4.369983e-15, 5.339081e-15, 
    3.394096e-15, 4.641842e-15, 2.53533e-15, 3.553219e-15, 2.479552e-15, 
    2.654226e-15, 2.369645e-15, 2.134004e-15, 1.862098e-15, 1.426799e-15, 
    1.520321e-15, 1.202028e-15, 7.913576e-15, 7.23552e-15, 7.293543e-15, 
    6.626987e-15, 6.163687e-15, 5.241716e-15, 3.979157e-15, 4.424375e-15, 
    3.632891e-15, 3.48735e-15, 4.700912e-15, 3.924698e-15, 6.806423e-15, 
    6.260124e-15, 6.581412e-15, 7.858377e-15, 4.318608e-15, 5.941917e-15, 
    3.220121e-15, 3.895999e-15, 2.166517e-15, 2.935467e-15, 1.573622e-15, 
    1.160591e-15, 8.485952e-16, 5.652149e-16, 6.884201e-15, 7.323716e-15, 
    6.55085e-15, 5.582475e-15, 4.782173e-15, 3.85205e-15, 3.765015e-15, 
    3.609275e-15, 3.227709e-15, 2.93022e-15, 3.560954e-15, 2.858876e-15, 
    6.137979e-15, 4.195046e-15, 7.495046e-15, 6.35156e-15, 5.636483e-15, 
    5.942557e-15, 4.477493e-15, 4.174828e-15, 3.095786e-15, 3.624407e-15, 
    1.254278e-15, 2.08641e-15, 4.001545e-16, 6.911144e-16, 7.48202e-15, 
    6.885734e-15, 5.079752e-15, 5.888907e-15, 3.795112e-15, 3.377093e-15, 
    3.062787e-15, 2.692418e-15, 2.65451e-15, 2.45308e-15, 2.78923e-15, 
    2.465794e-15, 3.850224e-15, 3.176389e-15, 5.266299e-15, 4.685611e-15, 
    4.946625e-15, 5.244917e-15, 4.364417e-15, 3.550307e-15, 3.534334e-15, 
    3.299222e-15, 2.697422e-15, 3.787945e-15, 1.167717e-15, 2.525167e-15, 
    6.276218e-15, 5.297466e-15, 5.1676e-15, 5.525802e-15, 3.417413e-15, 
    4.097268e-15, 2.457866e-15, 2.842509e-15, 2.232858e-15, 2.522557e-15, 
    2.567346e-15, 2.983146e-15, 3.265337e-15, 4.064088e-15, 4.811918e-15, 
    5.472775e-15, 5.31354e-15, 4.606652e-15, 3.504427e-15, 2.651055e-15, 
    2.823442e-15, 2.27553e-15, 3.925083e-15, 3.154056e-15, 3.437589e-15, 
    2.734318e-15, 4.436651e-15, 2.950101e-15, 4.890534e-15, 4.691103e-15, 
    4.111685e-15, 3.106033e-15, 2.910434e-15, 2.711416e-15, 2.833037e-15, 
    3.479252e-15, 3.594524e-15, 4.125144e-15, 4.281099e-15, 4.734018e-15, 
    5.134604e-15, 4.767636e-15, 4.403247e-15, 3.479004e-15, 2.77462e-15, 
    2.130765e-15, 1.991295e-15, 1.413641e-15, 1.872916e-15, 1.162105e-15, 
    1.750548e-15, 8.326406e-16, 2.877082e-15, 1.770668e-15, 4.086669e-15, 
    3.767423e-15, 3.236434e-15, 2.225336e-15, 2.737358e-15, 2.145992e-15, 
    3.599104e-15, 4.583496e-15, 4.867374e-15, 5.430777e-15, 4.855016e-15, 
    4.9001e-15, 4.388698e-15, 4.548574e-15, 3.450979e-15, 4.013146e-15, 
    2.568455e-15, 2.150284e-15, 1.232903e-15, 8.339763e-16, 5.31994e-16, 
    4.273464e-16, 3.986326e-16, 3.870426e-16,
  3.859466e-20, 3.197366e-20, 3.318957e-20, 2.835901e-20, 3.096967e-20, 
    2.790597e-20, 3.717757e-20, 3.172921e-20, 3.513364e-20, 3.796089e-20, 
    2.048221e-20, 2.815644e-20, 1.425774e-20, 1.788534e-20, 9.826356e-21, 
    1.478333e-20, 8.995481e-21, 9.949891e-21, 7.278588e-21, 7.983586e-21, 
    5.175844e-21, 6.968677e-21, 4.038358e-21, 5.57016e-21, 5.307167e-21, 
    7.034371e-21, 2.646687e-20, 2.134202e-20, 2.679619e-20, 2.600831e-20, 
    2.635985e-20, 3.091377e-20, 3.341582e-20, 3.913985e-20, 3.805067e-20, 
    3.387149e-20, 2.565964e-20, 2.826106e-20, 2.204825e-20, 2.217633e-20, 
    1.647893e-20, 1.889576e-20, 1.102599e-20, 1.295769e-20, 7.95323e-21, 
    9.050464e-21, 8.002476e-21, 8.310587e-21, 7.998517e-21, 9.649593e-21, 
    8.914999e-21, 1.046969e-20, 1.842461e-20, 1.574481e-20, 2.469892e-20, 
    3.160831e-20, 3.692493e-20, 4.107912e-20, 4.047177e-20, 3.93323e-20, 
    3.384807e-20, 2.922818e-20, 2.603266e-20, 2.404346e-20, 2.219478e-20, 
    1.72278e-20, 1.495536e-20, 1.066203e-20, 1.136104e-20, 1.019562e-20, 
    9.165241e-21, 7.605799e-21, 7.848362e-21, 7.211189e-21, 1.022542e-20, 
    8.139086e-21, 1.177355e-20, 1.068288e-20, 2.170885e-20, 2.754111e-20, 
    3.033704e-20, 3.295314e-20, 4.00093e-20, 3.502882e-20, 3.693372e-20, 
    3.252277e-20, 2.99299e-20, 3.119254e-20, 2.399069e-20, 2.662639e-20, 
    1.482789e-20, 1.930012e-20, 9.281394e-21, 1.121499e-20, 8.856137e-21, 
    1.000996e-20, 8.093362e-21, 9.805008e-21, 6.983829e-21, 6.456656e-21, 
    6.813702e-21, 5.515009e-21, 9.906847e-21, 8.002394e-21, 3.122836e-20, 
    3.101961e-20, 3.006088e-20, 3.444409e-20, 3.472684e-20, 3.916989e-20, 
    3.519745e-20, 3.35995e-20, 2.978461e-20, 2.768381e-20, 2.57899e-20, 
    2.196172e-20, 1.819628e-20, 1.374844e-20, 1.108158e-20, 9.516883e-21, 
    1.045608e-20, 9.623628e-21, 1.055746e-20, 1.101685e-20, 6.65069e-21, 
    8.908286e-21, 5.689938e-21, 5.842073e-21, 7.19647e-21, 5.824789e-21, 
    3.087369e-20, 3.208489e-20, 3.656291e-20, 3.302192e-20, 3.967798e-20, 
    3.584074e-20, 3.376265e-20, 2.656875e-20, 2.515385e-20, 2.389137e-20, 
    2.153548e-20, 1.876616e-20, 1.454673e-20, 1.147581e-20, 9.107737e-21, 
    9.268139e-21, 9.211432e-21, 8.730686e-21, 9.955649e-21, 8.540452e-21, 
    8.317836e-21, 8.908697e-21, 5.86266e-21, 6.641769e-21, 5.845337e-21, 
    6.343742e-21, 3.168747e-20, 2.968777e-20, 3.075636e-20, 2.876967e-20, 
    3.015892e-20, 2.433931e-20, 2.2768e-20, 1.638012e-20, 1.881792e-20, 
    1.505149e-20, 1.840721e-20, 1.77764e-20, 1.493811e-20, 1.821327e-20, 
    1.163144e-20, 1.58577e-20, 8.712373e-21, 1.217127e-20, 8.522404e-21, 
    9.117148e-21, 8.147931e-21, 7.344352e-21, 6.415801e-21, 4.925861e-21, 
    5.246363e-21, 4.154551e-21, 2.688139e-20, 2.460238e-20, 2.47975e-20, 
    2.255478e-20, 2.099432e-20, 1.788456e-20, 1.361489e-20, 1.512215e-20, 
    1.244145e-20, 1.194785e-20, 1.605742e-20, 1.34304e-20, 2.315879e-20, 
    2.131925e-20, 2.240134e-20, 2.669596e-20, 1.476426e-20, 2.024685e-20, 
    1.104088e-20, 1.333318e-20, 7.455288e-21, 1.007377e-20, 5.428922e-21, 
    4.012189e-21, 2.938294e-21, 1.95914e-21, 2.342053e-20, 2.489896e-20, 
    2.229844e-20, 1.903465e-20, 1.633212e-20, 1.318428e-20, 1.288934e-20, 
    1.236137e-20, 1.106664e-20, 1.005593e-20, 1.219751e-20, 9.813363e-21, 
    2.090768e-20, 1.434601e-20, 2.547497e-20, 2.162727e-20, 1.921685e-20, 
    2.024901e-20, 1.530186e-20, 1.427756e-20, 1.061858e-20, 1.241269e-20, 
    4.333986e-21, 7.181925e-21, 1.386536e-21, 2.394665e-21, 2.543119e-20, 
    2.342569e-20, 1.733761e-20, 2.006814e-20, 1.299134e-20, 1.157374e-20, 
    1.050647e-20, 9.247123e-21, 9.118114e-21, 8.432227e-21, 9.576496e-21, 
    8.475536e-21, 1.317809e-20, 1.089237e-20, 1.796756e-20, 1.600569e-20, 
    1.688788e-20, 1.789537e-20, 1.491928e-20, 1.21614e-20, 1.210722e-20, 
    1.130944e-20, 9.264151e-21, 1.296705e-20, 4.036677e-21, 8.67776e-21, 
    2.137347e-20, 1.807278e-20, 1.76343e-20, 1.884343e-20, 1.171057e-20, 
    1.401494e-20, 8.448531e-21, 9.757704e-21, 7.681584e-21, 8.668873e-21, 
    8.82139e-21, 1.023583e-20, 1.11944e-20, 1.390257e-20, 1.643266e-20, 
    1.86645e-20, 1.812705e-20, 1.57387e-20, 1.200578e-20, 9.106355e-21, 
    9.69286e-21, 7.8271e-21, 1.343171e-20, 1.081652e-20, 1.177903e-20, 
    9.389691e-21, 1.516368e-20, 1.012351e-20, 1.669835e-20, 1.602426e-20, 
    1.406376e-20, 1.065339e-20, 9.988667e-21, 9.311768e-21, 9.725491e-21, 
    1.192038e-20, 1.231135e-20, 1.410934e-20, 1.463731e-20, 1.616934e-20, 
    1.752287e-20, 1.628298e-20, 1.505067e-20, 1.191954e-20, 9.526799e-21, 
    7.333301e-21, 6.85719e-21, 4.880749e-21, 6.452773e-21, 4.017393e-21, 
    6.034414e-21, 2.883271e-21, 9.875268e-21, 6.103224e-21, 1.397905e-20, 
    1.289751e-20, 1.109627e-20, 7.655931e-21, 9.400035e-21, 7.38526e-21, 
    1.232689e-20, 1.566039e-20, 1.662008e-20, 1.852276e-20, 1.657832e-20, 
    1.673067e-20, 1.500144e-20, 1.554229e-20, 1.182446e-20, 1.373003e-20, 
    8.825167e-21, 7.399903e-21, 4.260591e-21, 2.887878e-21, 1.844055e-21, 
    1.481013e-21, 1.381246e-21, 1.340955e-21,
  2.833738e-26, 2.349564e-26, 2.438506e-26, 2.085076e-26, 2.276113e-26, 
    2.051918e-26, 2.730139e-26, 2.331681e-26, 2.580687e-26, 2.787407e-26, 
    1.508225e-26, 2.070251e-26, 1.05172e-26, 1.317857e-26, 7.261474e-27, 
    1.090297e-26, 6.650332e-27, 7.352317e-27, 5.386588e-27, 5.905672e-27, 
    3.836718e-27, 5.158324e-27, 2.996983e-27, 4.127572e-27, 3.933597e-27, 
    5.206716e-27, 1.946574e-26, 1.571232e-26, 1.970683e-26, 1.913003e-26, 
    1.938739e-26, 2.272023e-26, 2.455054e-26, 2.873592e-26, 2.79397e-26, 
    2.488382e-26, 1.887475e-26, 2.077908e-26, 1.622976e-26, 1.63236e-26, 
    1.214708e-26, 1.391941e-26, 8.143423e-27, 9.562673e-27, 5.883326e-27, 
    6.690782e-27, 5.919578e-27, 6.146361e-27, 5.916663e-27, 7.131479e-27, 
    6.591119e-27, 7.734501e-27, 1.357398e-26, 1.160851e-26, 1.817127e-26, 
    2.322836e-26, 2.711667e-26, 3.015336e-26, 2.970947e-26, 2.88766e-26, 
    2.486669e-26, 2.148686e-26, 1.914786e-26, 1.769126e-26, 1.633712e-26, 
    1.269636e-26, 1.102922e-26, 7.8759e-27, 8.389668e-27, 7.533005e-27, 
    6.775218e-27, 5.62754e-27, 5.806126e-27, 5.33695e-27, 7.554911e-27, 
    6.020133e-27, 8.692791e-27, 7.891221e-27, 1.59811e-26, 2.025212e-26, 
    2.229826e-26, 2.421213e-26, 2.937145e-26, 2.573021e-26, 2.71231e-26, 
    2.389732e-26, 2.200035e-26, 2.292419e-26, 1.765261e-26, 1.958253e-26, 
    1.093568e-26, 1.421584e-26, 6.860661e-27, 8.28233e-27, 6.547813e-27, 
    7.396488e-27, 5.986478e-27, 7.245774e-27, 5.169486e-27, 4.781085e-27, 
    5.044159e-27, 4.086899e-27, 7.320664e-27, 5.919516e-27, 2.29504e-26, 
    2.279767e-26, 2.209619e-26, 2.530259e-26, 2.550938e-26, 2.875788e-26, 
    2.585353e-26, 2.468489e-26, 2.189404e-26, 2.035657e-26, 1.897012e-26, 
    1.616637e-26, 1.340656e-26, 1.014333e-26, 8.184281e-27, 7.033874e-27, 
    7.724499e-27, 7.112383e-27, 7.799029e-27, 8.13671e-27, 4.92406e-27, 
    6.586181e-27, 4.215901e-27, 4.328076e-27, 5.326109e-27, 4.315333e-27, 
    2.26909e-26, 2.3577e-26, 2.685198e-26, 2.426244e-26, 2.912927e-26, 
    2.632393e-26, 2.480422e-26, 1.954033e-26, 1.850441e-26, 1.757987e-26, 
    1.585407e-26, 1.382439e-26, 1.072932e-26, 8.474011e-27, 6.732916e-27, 
    6.850911e-27, 6.809198e-27, 6.455509e-27, 7.356552e-27, 6.315527e-27, 
    6.151697e-27, 6.586483e-27, 4.343256e-27, 4.917487e-27, 4.330483e-27, 
    4.697874e-27, 2.328627e-26, 2.182317e-26, 2.260506e-26, 2.115131e-26, 
    2.216793e-26, 1.790793e-26, 1.675704e-26, 1.20746e-26, 1.386234e-26, 
    1.109977e-26, 1.356122e-26, 1.309868e-26, 1.101657e-26, 1.341902e-26, 
    8.588373e-27, 1.169133e-26, 6.442033e-27, 8.985003e-27, 6.302245e-27, 
    6.739838e-27, 6.026644e-27, 5.435019e-27, 4.750978e-27, 3.652265e-27, 
    3.888742e-27, 3.082815e-27, 1.97692e-26, 1.810058e-26, 1.824346e-26, 
    1.660085e-26, 1.545754e-26, 1.3178e-26, 1.004529e-26, 1.115162e-26, 
    9.183485e-27, 8.820855e-27, 1.183786e-26, 9.909825e-27, 1.70433e-26, 
    1.569564e-26, 1.648844e-26, 1.963345e-26, 1.088897e-26, 1.490977e-26, 
    8.15437e-27, 9.838433e-27, 5.516713e-27, 7.443406e-27, 4.023406e-27, 
    2.97765e-27, 2.18361e-27, 1.458113e-27, 1.723502e-26, 1.831776e-26, 
    1.641306e-26, 1.402123e-26, 1.203939e-26, 9.729085e-27, 9.512472e-27, 
    9.124659e-27, 8.173306e-27, 7.43029e-27, 9.004279e-27, 7.251919e-27, 
    1.539405e-26, 1.0582e-26, 1.873953e-26, 1.592133e-26, 1.415479e-26, 
    1.491135e-26, 1.128349e-26, 1.053176e-26, 7.843959e-27, 9.162353e-27, 
    3.215338e-27, 5.315396e-27, 1.032859e-27, 1.781039e-27, 1.870747e-26, 
    1.72388e-26, 1.277689e-26, 1.477878e-26, 9.587386e-27, 8.545974e-27, 
    7.761541e-27, 6.835452e-27, 6.740549e-27, 6.235884e-27, 7.077719e-27, 
    6.267755e-27, 9.72454e-27, 8.045213e-27, 1.323886e-26, 1.179991e-26, 
    1.244705e-26, 1.318592e-26, 1.100274e-26, 8.97775e-27, 8.937947e-27, 
    8.351745e-27, 6.847977e-27, 9.569549e-27, 2.99574e-27, 6.416565e-27, 
    1.573536e-26, 1.331601e-26, 1.299447e-26, 1.388104e-26, 8.646513e-27, 
    1.033898e-26, 6.247882e-27, 7.210987e-27, 5.68334e-27, 6.410026e-27, 
    6.522248e-27, 7.562569e-27, 8.267205e-27, 1.025649e-26, 1.211314e-26, 
    1.374986e-26, 1.33558e-26, 1.160403e-26, 8.863418e-27, 6.731899e-27, 
    7.163299e-27, 5.790473e-27, 9.910785e-27, 7.989458e-27, 8.696816e-27, 
    6.940321e-27, 1.11821e-26, 7.479984e-27, 1.230803e-26, 1.181353e-26, 
    1.037481e-26, 7.869549e-27, 7.38083e-27, 6.883004e-27, 7.187297e-27, 
    8.800673e-27, 9.087913e-27, 1.040827e-26, 1.07958e-26, 1.191997e-26, 
    1.291276e-26, 1.200334e-26, 1.109916e-26, 8.800055e-27, 7.041167e-27, 
    5.426881e-27, 5.076197e-27, 3.618973e-27, 4.778223e-27, 2.981494e-27, 
    4.469876e-27, 2.142885e-27, 7.297443e-27, 4.520599e-27, 1.031263e-26, 
    9.518467e-27, 8.195081e-27, 5.664452e-27, 6.94793e-27, 5.465145e-27, 
    9.099324e-27, 1.154657e-26, 1.225062e-26, 1.364595e-26, 1.221999e-26, 
    1.233174e-26, 1.106304e-26, 1.145991e-26, 8.730197e-27, 1.012982e-26, 
    6.525027e-27, 5.475928e-27, 3.161135e-27, 2.146295e-27, 1.372713e-27, 
    1.103088e-27, 1.028926e-27, 9.989671e-28,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.004388433, 0.004385842, 0.004386347, 0.004384255, 0.004385417, 
    0.004384046, 0.00438791, 0.004385737, 0.004387126, 0.004388203, 
    0.004380189, 0.004384162, 0.004376089, 0.004378616, 0.004372278, 
    0.004376479, 0.004371433, 0.004372405, 0.004369493, 0.004370327, 
    0.004366594, 0.004369108, 0.004364669, 0.004367197, 0.004366799, 
    0.00436919, 0.004383367, 0.004380682, 0.004383525, 0.004383143, 
    0.004383316, 0.004385392, 0.004386434, 0.004388635, 0.004388236, 
    0.004386622, 0.004382971, 0.004384214, 0.004381092, 0.004381163, 
    0.004377687, 0.004379254, 0.00437342, 0.004375078, 0.004370292, 
    0.004371495, 0.004370348, 0.004370696, 0.004370343, 0.004372107, 
    0.004371351, 0.004372905, 0.004378959, 0.004377177, 0.004382491, 
    0.004385681, 0.004387814, 0.004389324, 0.00438911, 0.004388703, 
    0.004386613, 0.004384653, 0.004383158, 0.004382158, 0.004381173, 
    0.00437818, 0.004376608, 0.004373082, 0.004373723, 0.004372641, 
    0.004371615, 0.004369886, 0.004370171, 0.004369408, 0.004372673, 
    0.004370501, 0.004374086, 0.004373105, 0.004380887, 0.004383879, 
    0.004385136, 0.004386249, 0.004388946, 0.004387083, 0.004387817, 
    0.004386074, 0.004384965, 0.004385515, 0.00438213, 0.004383445, 
    0.004376515, 0.004379498, 0.004371734, 0.004373591, 0.00437129, 
    0.004372465, 0.00437045, 0.004372264, 0.004369126, 0.004368441, 
    0.004368908, 0.004367118, 0.004372363, 0.004370346, 0.004385529, 
    0.004385439, 0.004385023, 0.004386851, 0.004386964, 0.004388645, 
    0.004387151, 0.004386513, 0.004384902, 0.004383946, 0.004383038, 
    0.004381043, 0.004378813, 0.004375702, 0.004373471, 0.004371976, 
    0.004372894, 0.004372083, 0.004372988, 0.004373414, 0.004368696, 
    0.004371343, 0.004367376, 0.004367596, 0.004369389, 0.004367571, 
    0.004385377, 0.004385892, 0.004387677, 0.00438628, 0.004388829, 
    0.0043874, 0.004386577, 0.004383414, 0.004382723, 0.004382077, 
    0.004380806, 0.004379173, 0.004376309, 0.004373822, 0.004371556, 
    0.004371722, 0.004371663, 0.004371155, 0.004372411, 0.004370949, 
    0.004370702, 0.004371346, 0.004367625, 0.004368688, 0.004367601, 
    0.004368293, 0.004385725, 0.004384859, 0.004385327, 0.004384445, 
    0.004385064, 0.004382305, 0.004381478, 0.004377615, 0.004379204, 
    0.00437668, 0.004378949, 0.004378546, 0.00437659, 0.004378828, 
    0.004373956, 0.004377251, 0.004371135, 0.004374417, 0.00437093, 
    0.004371565, 0.004370514, 0.004369571, 0.004368389, 0.004366203, 
    0.004366709, 0.004364885, 0.004383567, 0.004382442, 0.004382544, 
    0.004381368, 0.004380499, 0.004378618, 0.0043756, 0.004376736, 
    0.004374654, 0.004374235, 0.0043774, 0.004375453, 0.004381691, 
    0.004380679, 0.004381284, 0.004383476, 0.004376469, 0.004380062, 
    0.004373434, 0.004375379, 0.004369705, 0.004372522, 0.004366988, 
    0.004364616, 0.004362401, 0.004359795, 0.004381831, 0.004382595, 
    0.00438123, 0.004379335, 0.004377587, 0.004375259, 0.004375023, 
    0.004374586, 0.004373459, 0.00437251, 0.004374444, 0.004372272, 
    0.004380437, 0.004376159, 0.004382881, 0.004380852, 0.004379448, 
    0.004380067, 0.004376866, 0.004376111, 0.004373042, 0.00437463, 
    0.004365198, 0.004369367, 0.004357825, 0.004361044, 0.004382862, 
    0.004381835, 0.00437826, 0.004379961, 0.004375106, 0.00437391, 
    0.004372941, 0.004371698, 0.004371566, 0.00437083, 0.004372036, 
    0.004370878, 0.004375254, 0.004373299, 0.004378672, 0.004377361, 
    0.004377965, 0.004378626, 0.004376588, 0.004374413, 0.004374372, 
    0.004373674, 0.004371698, 0.004375086, 0.00436465, 0.004371082, 
    0.004380716, 0.004378732, 0.004378456, 0.004379223, 0.00437403, 
    0.00437591, 0.004370848, 0.004372217, 0.004369976, 0.004371089, 
    0.004371252, 0.004372683, 0.004373573, 0.004375822, 0.004377655, 
    0.004379112, 0.004378774, 0.004377174, 0.004374282, 0.004371551, 
    0.004372149, 0.004370146, 0.004375457, 0.004373227, 0.004374087, 
    0.004371846, 0.004376764, 0.004372559, 0.004377838, 0.004377376, 
    0.004375947, 0.004373072, 0.004372444, 0.004371764, 0.004372185, 
    0.004374209, 0.004374544, 0.004375983, 0.004376378, 0.004377477, 
    0.004378385, 0.004377554, 0.004376681, 0.004374211, 0.004371983, 
    0.004369557, 0.004368966, 0.004366121, 0.004368429, 0.004364613, 
    0.004367846, 0.004362258, 0.004372323, 0.004367952, 0.004375884, 
    0.00437503, 0.00437348, 0.004369939, 0.004371856, 0.004369617, 
    0.004374557, 0.004377116, 0.004377785, 0.004379022, 0.004377757, 
    0.00437786, 0.004376648, 0.004377038, 0.004374129, 0.004375692, 
    0.004371255, 0.004369636, 0.004365074, 0.004362277, 0.004359441, 
    0.004358187, 0.004357806, 0.004357647,
  8.330007e-06, 8.329982e-06, 8.329994e-06, 8.330192e-06, 8.329985e-06, 
    8.330273e-06, 8.330014e-06, 8.329971e-06, 8.330006e-06, 8.33002e-06, 
    8.331656e-06, 8.330229e-06, 8.33318e-06, 8.332298e-06, 8.3345e-06, 
    8.33303e-06, 8.334793e-06, 8.334483e-06, 8.335464e-06, 8.335188e-06, 
    8.336357e-06, 8.335592e-06, 8.336983e-06, 8.33619e-06, 8.336307e-06, 
    8.335562e-06, 8.330545e-06, 8.331474e-06, 8.330483e-06, 8.330619e-06, 
    8.330564e-06, 8.329976e-06, 8.329971e-06, 8.330025e-06, 8.33002e-06, 
    8.329989e-06, 8.33068e-06, 8.330228e-06, 8.331406e-06, 8.331381e-06, 
    8.332636e-06, 8.332075e-06, 8.334137e-06, 8.333569e-06, 8.335201e-06, 
    8.334794e-06, 8.335177e-06, 8.335065e-06, 8.335179e-06, 8.334582e-06, 
    8.334838e-06, 8.334317e-06, 8.332176e-06, 8.332811e-06, 8.330869e-06, 
    8.329947e-06, 8.330008e-06, 8.330026e-06, 8.330024e-06, 8.330015e-06, 
    8.329989e-06, 8.330059e-06, 8.330632e-06, 8.331007e-06, 8.331376e-06, 
    8.332409e-06, 8.332996e-06, 8.334238e-06, 8.334038e-06, 8.334391e-06, 
    8.334755e-06, 8.335328e-06, 8.335237e-06, 8.335482e-06, 8.334398e-06, 
    8.335115e-06, 8.333918e-06, 8.334248e-06, 8.331393e-06, 8.330354e-06, 
    8.329944e-06, 8.329988e-06, 8.33002e-06, 8.329996e-06, 8.330005e-06, 
    8.329998e-06, 8.329978e-06, 8.329992e-06, 8.331017e-06, 8.330519e-06, 
    8.333031e-06, 8.331971e-06, 8.334713e-06, 8.334081e-06, 8.334865e-06, 
    8.334471e-06, 8.335136e-06, 8.334539e-06, 8.335579e-06, 8.335792e-06, 
    8.335644e-06, 8.336232e-06, 8.334503e-06, 8.335169e-06, 8.329988e-06, 
    8.329986e-06, 8.329983e-06, 8.329992e-06, 8.329996e-06, 8.330021e-06, 
    8.330007e-06, 8.329993e-06, 8.329983e-06, 8.330328e-06, 8.33067e-06, 
    8.331415e-06, 8.332217e-06, 8.33333e-06, 8.334122e-06, 8.334637e-06, 
    8.334328e-06, 8.3346e-06, 8.334292e-06, 8.33415e-06, 8.335706e-06, 
    8.334835e-06, 8.336148e-06, 8.336079e-06, 8.335484e-06, 8.336087e-06, 
    8.329986e-06, 8.329998e-06, 8.33001e-06, 8.330001e-06, 8.330024e-06, 
    8.330004e-06, 8.329983e-06, 8.330512e-06, 8.330794e-06, 8.331029e-06, 
    8.331508e-06, 8.332103e-06, 8.333119e-06, 8.333992e-06, 8.33478e-06, 
    8.334724e-06, 8.334742e-06, 8.334908e-06, 8.334486e-06, 8.334977e-06, 
    8.335051e-06, 8.334845e-06, 8.33607e-06, 8.335726e-06, 8.336078e-06, 
    8.335857e-06, 8.329996e-06, 8.329981e-06, 8.329986e-06, 8.330133e-06, 
    8.329974e-06, 8.330924e-06, 8.331228e-06, 8.332639e-06, 8.332087e-06, 
    8.332983e-06, 8.332186e-06, 8.332324e-06, 8.332977e-06, 8.332235e-06, 
    8.333928e-06, 8.332758e-06, 8.334914e-06, 8.333748e-06, 8.334984e-06, 
    8.334776e-06, 8.335128e-06, 8.335431e-06, 8.335822e-06, 8.336507e-06, 
    8.336353e-06, 8.33693e-06, 8.330474e-06, 8.330884e-06, 8.330863e-06, 
    8.3313e-06, 8.331614e-06, 8.332308e-06, 8.333377e-06, 8.332984e-06, 
    8.333718e-06, 8.333858e-06, 8.33275e-06, 8.333421e-06, 8.331168e-06, 
    8.331525e-06, 8.331324e-06, 8.330498e-06, 8.333053e-06, 8.331755e-06, 
    8.334132e-06, 8.333458e-06, 8.335385e-06, 8.334427e-06, 8.336265e-06, 
    8.336976e-06, 8.337699e-06, 8.338437e-06, 8.331123e-06, 8.330845e-06, 
    8.331355e-06, 8.332022e-06, 8.332673e-06, 8.333497e-06, 8.333589e-06, 
    8.333735e-06, 8.334133e-06, 8.334455e-06, 8.333767e-06, 8.334537e-06, 
    8.331576e-06, 8.333172e-06, 8.330724e-06, 8.331458e-06, 8.33199e-06, 
    8.331773e-06, 8.332942e-06, 8.333208e-06, 8.334257e-06, 8.333727e-06, 
    8.336789e-06, 8.335472e-06, 8.339034e-06, 8.338077e-06, 8.330743e-06, 
    8.33113e-06, 8.33242e-06, 8.331815e-06, 8.33356e-06, 8.333969e-06, 
    8.334311e-06, 8.334718e-06, 8.334773e-06, 8.335012e-06, 8.334617e-06, 
    8.335003e-06, 8.333499e-06, 8.334183e-06, 8.332294e-06, 8.332754e-06, 
    8.332549e-06, 8.33231e-06, 8.33304e-06, 8.333775e-06, 8.333815e-06, 
    8.334043e-06, 8.334629e-06, 8.333567e-06, 8.336907e-06, 8.334848e-06, 
    8.331544e-06, 8.332235e-06, 8.332363e-06, 8.332093e-06, 8.333927e-06, 
    8.333271e-06, 8.335011e-06, 8.334555e-06, 8.335304e-06, 8.334932e-06, 
    8.334876e-06, 8.334397e-06, 8.334087e-06, 8.333296e-06, 8.332646e-06, 
    8.332135e-06, 8.332257e-06, 8.332816e-06, 8.333825e-06, 8.334767e-06, 
    8.334559e-06, 8.335248e-06, 8.333435e-06, 8.334196e-06, 8.333895e-06, 
    8.334676e-06, 8.332968e-06, 8.334352e-06, 8.332595e-06, 8.332759e-06, 
    8.333258e-06, 8.334229e-06, 8.334478e-06, 8.334695e-06, 8.334567e-06, 
    8.333855e-06, 8.333747e-06, 8.333252e-06, 8.333102e-06, 8.332725e-06, 
    8.332398e-06, 8.33269e-06, 8.33299e-06, 8.333865e-06, 8.334619e-06, 
    8.335431e-06, 8.335635e-06, 8.336488e-06, 8.335762e-06, 8.336913e-06, 
    8.335885e-06, 8.337667e-06, 8.334468e-06, 8.335905e-06, 8.333289e-06, 
    8.333588e-06, 8.334096e-06, 8.33528e-06, 8.334673e-06, 8.335393e-06, 
    8.333745e-06, 8.332823e-06, 8.332611e-06, 8.332162e-06, 8.332622e-06, 
    8.332586e-06, 8.33302e-06, 8.332882e-06, 8.333894e-06, 8.333355e-06, 
    8.334868e-06, 8.335394e-06, 8.33686e-06, 8.337706e-06, 8.338578e-06, 
    8.33894e-06, 8.339052e-06, 8.339097e-06,
  1.682193e-10, 1.682733e-10, 1.68263e-10, 1.68323e-10, 1.682826e-10, 
    1.683319e-10, 1.682306e-10, 1.682752e-10, 1.682468e-10, 1.682246e-10, 
    1.68492e-10, 1.68327e-10, 1.686673e-10, 1.68561e-10, 1.688294e-10, 
    1.686503e-10, 1.688657e-10, 1.68825e-10, 1.689495e-10, 1.689139e-10, 
    1.69072e-10, 1.68966e-10, 1.691554e-10, 1.690471e-10, 1.690637e-10, 
    1.689624e-10, 1.683609e-10, 1.684712e-10, 1.683542e-10, 1.683699e-10, 
    1.68363e-10, 1.682828e-10, 1.682603e-10, 1.682157e-10, 1.682239e-10, 
    1.68257e-10, 1.68377e-10, 1.683255e-10, 1.68457e-10, 1.68454e-10, 
    1.686004e-10, 1.685343e-10, 1.687817e-10, 1.687114e-10, 1.689154e-10, 
    1.688639e-10, 1.689128e-10, 1.688981e-10, 1.68913e-10, 1.688376e-10, 
    1.688698e-10, 1.688038e-10, 1.685466e-10, 1.686218e-10, 1.683975e-10, 
    1.682756e-10, 1.682324e-10, 1.682014e-10, 1.682058e-10, 1.68214e-10, 
    1.682571e-10, 1.68307e-10, 1.6837e-10, 1.68412e-10, 1.684536e-10, 
    1.685778e-10, 1.686453e-10, 1.687956e-10, 1.68769e-10, 1.688145e-10, 
    1.688588e-10, 1.689325e-10, 1.689204e-10, 1.689528e-10, 1.688137e-10, 
    1.689059e-10, 1.687538e-10, 1.687953e-10, 1.684624e-10, 1.683395e-10, 
    1.682883e-10, 1.682649e-10, 1.682091e-10, 1.682474e-10, 1.682322e-10, 
    1.68269e-10, 1.68295e-10, 1.682807e-10, 1.684132e-10, 1.683578e-10, 
    1.686493e-10, 1.685235e-10, 1.688536e-10, 1.687745e-10, 1.688727e-10, 
    1.688227e-10, 1.689082e-10, 1.688313e-10, 1.68965e-10, 1.689939e-10, 
    1.689741e-10, 1.690511e-10, 1.688269e-10, 1.689126e-10, 1.682803e-10, 
    1.682821e-10, 1.682933e-10, 1.682522e-10, 1.6825e-10, 1.682154e-10, 
    1.682463e-10, 1.682594e-10, 1.682972e-10, 1.683367e-10, 1.683748e-10, 
    1.684587e-10, 1.685523e-10, 1.686842e-10, 1.687796e-10, 1.688436e-10, 
    1.688045e-10, 1.68839e-10, 1.688004e-10, 1.687824e-10, 1.689829e-10, 
    1.6887e-10, 1.6904e-10, 1.690306e-10, 1.689534e-10, 1.690317e-10, 
    1.682835e-10, 1.682728e-10, 1.682353e-10, 1.682647e-10, 1.682117e-10, 
    1.68241e-10, 1.682577e-10, 1.683584e-10, 1.683882e-10, 1.684151e-10, 
    1.684689e-10, 1.685377e-10, 1.686585e-10, 1.687643e-10, 1.688615e-10, 
    1.688544e-10, 1.688569e-10, 1.688783e-10, 1.688249e-10, 1.688872e-10, 
    1.688974e-10, 1.688703e-10, 1.690294e-10, 1.689839e-10, 1.690304e-10, 
    1.690009e-10, 1.682764e-10, 1.682985e-10, 1.682846e-10, 1.683156e-10, 
    1.682917e-10, 1.684048e-10, 1.684394e-10, 1.686026e-10, 1.685362e-10, 
    1.686427e-10, 1.685472e-10, 1.68564e-10, 1.686451e-10, 1.685525e-10, 
    1.68758e-10, 1.686176e-10, 1.688792e-10, 1.687377e-10, 1.68888e-10, 
    1.688611e-10, 1.689059e-10, 1.689459e-10, 1.689966e-10, 1.690897e-10, 
    1.690682e-10, 1.691466e-10, 1.683527e-10, 1.683995e-10, 1.683958e-10, 
    1.684452e-10, 1.684816e-10, 1.685613e-10, 1.686889e-10, 1.686411e-10, 
    1.687295e-10, 1.687471e-10, 1.68613e-10, 1.686949e-10, 1.684312e-10, 
    1.684732e-10, 1.684485e-10, 1.683561e-10, 1.686514e-10, 1.684993e-10, 
    1.687811e-10, 1.686985e-10, 1.689401e-10, 1.688193e-10, 1.690563e-10, 
    1.691568e-10, 1.692537e-10, 1.693647e-10, 1.684256e-10, 1.683937e-10, 
    1.684512e-10, 1.685301e-10, 1.686047e-10, 1.687034e-10, 1.687138e-10, 
    1.687322e-10, 1.687804e-10, 1.688208e-10, 1.687375e-10, 1.688309e-10, 
    1.68482e-10, 1.686649e-10, 1.683812e-10, 1.684658e-10, 1.685256e-10, 
    1.684998e-10, 1.686357e-10, 1.686676e-10, 1.687974e-10, 1.687306e-10, 
    1.691316e-10, 1.689536e-10, 1.694509e-10, 1.693111e-10, 1.683824e-10, 
    1.684257e-10, 1.685758e-10, 1.685044e-10, 1.687103e-10, 1.687609e-10, 
    1.688025e-10, 1.688549e-10, 1.688609e-10, 1.688921e-10, 1.68841e-10, 
    1.688903e-10, 1.687036e-10, 1.68787e-10, 1.685592e-10, 1.686143e-10, 
    1.685891e-10, 1.685612e-10, 1.686474e-10, 1.687387e-10, 1.687415e-10, 
    1.687706e-10, 1.688516e-10, 1.687111e-10, 1.691532e-10, 1.688784e-10, 
    1.684728e-10, 1.685553e-10, 1.68568e-10, 1.685359e-10, 1.687558e-10, 
    1.686759e-10, 1.688914e-10, 1.688333e-10, 1.689288e-10, 1.688813e-10, 
    1.688742e-10, 1.688134e-10, 1.687753e-10, 1.686794e-10, 1.686017e-10, 
    1.685406e-10, 1.685549e-10, 1.68622e-10, 1.687445e-10, 1.688611e-10, 
    1.688355e-10, 1.689216e-10, 1.686953e-10, 1.687897e-10, 1.687529e-10, 
    1.688489e-10, 1.686396e-10, 1.688155e-10, 1.685945e-10, 1.68614e-10, 
    1.686743e-10, 1.687956e-10, 1.688236e-10, 1.688521e-10, 1.688346e-10, 
    1.687478e-10, 1.687339e-10, 1.68673e-10, 1.686559e-10, 1.686098e-10, 
    1.685714e-10, 1.686063e-10, 1.686428e-10, 1.687481e-10, 1.688427e-10, 
    1.689463e-10, 1.68972e-10, 1.690915e-10, 1.689932e-10, 1.691545e-10, 
    1.690157e-10, 1.692571e-10, 1.688268e-10, 1.690132e-10, 1.686773e-10, 
    1.687136e-10, 1.687784e-10, 1.689291e-10, 1.688485e-10, 1.689431e-10, 
    1.687334e-10, 1.68624e-10, 1.685967e-10, 1.685442e-10, 1.685979e-10, 
    1.685935e-10, 1.686449e-10, 1.686284e-10, 1.687516e-10, 1.686854e-10, 
    1.688738e-10, 1.689426e-10, 1.691381e-10, 1.692579e-10, 1.693814e-10, 
    1.694356e-10, 1.694522e-10, 1.694591e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  1.047567, 1.028503, 1.03221, 1.016824, 1.025361, 1.015284, 1.043704, 
    1.027745, 1.037935, 1.045853, 0.986935, 1.016138, 0.956573, 0.9752231, 
    0.9283484, 0.9594749, 0.9220675, 0.9292492, 0.9076329, 0.9138277, 
    0.8861535, 0.9047733, 0.8717993, 0.8906027, 0.8876613, 0.905387, 
    1.010266, 0.9905719, 1.011432, 1.008625, 1.009885, 1.025184, 1.032889, 
    1.049025, 1.046097, 1.034246, 1.007362, 1.016493, 0.9934793, 0.9939992, 
    0.9683524, 0.9799193, 0.9367741, 0.9490449, 0.9135692, 0.9224957, 
    0.9139882, 0.9165685, 0.9139546, 0.9270451, 0.9214372, 0.9329537, 
    0.9777529, 0.9645946, 1.003817, 1.027368, 1.043004, 1.054092, 1.052524, 
    1.049536, 1.034177, 1.019729, 1.008712, 1.00134, 0.994074, 0.972062, 
    0.9604083, 0.9342909, 0.9390084, 0.9310175, 0.9233837, 0.9105592, 
    0.9126707, 0.9070185, 0.9312297, 0.9151409, 0.9416945, 0.9344347, 
    0.9920909, 1.01403, 1.023343, 1.031497, 1.051319, 1.037632, 1.043028, 
    1.03019, 1.022027, 1.026065, 1.001138, 1.010832, 0.9597175, 0.9817472, 
    0.9242741, 0.9380404, 0.9209737, 0.9296843, 0.9147566, 0.9281918, 
    0.9049152, 0.8998429, 0.9033091, 0.8899942, 0.9289362, 0.9139875, 
    1.026178, 1.025519, 1.022452, 1.035932, 1.036757, 1.049105, 1.038118, 
    1.033438, 1.021555, 1.014522, 1.007835, 0.9931267, 0.9766885, 0.9536859, 
    0.9371482, 0.9260553, 0.9328584, 0.9268522, 0.9335661, 0.9367126, 
    0.9017431, 0.9213845, 0.8919098, 0.8935419, 0.9068838, 0.893358, 
    1.025057, 1.028846, 1.041994, 1.031705, 1.050449, 1.039958, 1.033923, 
    1.010628, 1.005508, 1.000758, 0.991375, 0.9793273, 0.958178, 0.9397627, 
    0.9229398, 0.9241729, 0.9237387, 0.9199783, 0.929291, 0.9184492, 
    0.9166284, 0.9213877, 0.8937604, 0.9016566, 0.8935766, 0.8987184, 
    1.027615, 1.021239, 1.024684, 1.018205, 1.022769, 1.002464, 0.9963732, 
    0.9678538, 0.9795641, 0.9609265, 0.9776721, 0.9747053, 0.9603152, 
    0.976768, 0.940777, 0.9651807, 0.9198321, 0.9442208, 0.9183028, 
    0.9230126, 0.915215, 0.9082285, 0.8994377, 0.8832067, 0.8869665, 
    0.8733879, 1.011732, 1.003455, 1.004186, 0.9955229, 0.989114, 0.9752194, 
    0.9529161, 0.9613059, 0.9459029, 0.9428091, 0.9662099, 0.9518434, 
    0.9979162, 0.9904768, 0.9949074, 1.011078, 0.9593709, 0.9859198, 
    0.9368745, 0.9512738, 0.9092246, 0.9301445, 0.8890356, 0.871437, 
    0.8548695, 0.8354861, 0.998939, 1.004564, 0.9944929, 0.9805503, 
    0.9676108, 0.9503955, 0.9486342, 0.9454071, 0.9370478, 0.930016, 
    0.9443853, 0.9282531, 0.9887484, 0.9570658, 1.006688, 0.9917545, 
    0.9813731, 0.9859291, 0.962265, 0.9566838, 0.9339904, 0.9457251, 
    0.8757804, 0.9067505, 0.8207223, 0.8447925, 1.006528, 0.998959, 
    0.9725959, 0.9851432, 0.9492466, 0.9404021, 0.9332107, 0.9240122, 
    0.92302, 0.9175683, 0.9265011, 0.9179217, 0.9503588, 0.9358695, 
    0.9756123, 0.9659443, 0.9703929, 0.9752706, 0.9602131, 0.9441588, 
    0.943818, 0.9386674, 0.9241425, 0.9491011, 0.8717759, 0.9195554, 
    0.9907026, 0.9761087, 0.9740263, 0.9796805, 0.9412888, 0.9552062, 
    0.9177015, 0.9278442, 0.911224, 0.9194841, 0.920699, 0.9313039, 
    0.9379032, 0.9545678, 0.9681191, 0.9788609, 0.9763637, 0.9645628, 
    0.9431769, 0.9229291, 0.9273657, 0.9124876, 0.9518511, 0.9353523, 
    0.9417297, 0.9250972, 0.9615283, 0.9305019, 0.9694517, 0.9660397, 
    0.9554824, 0.9342312, 0.9295303, 0.9245057, 0.9276068, 0.9426342, 
    0.9450963, 0.9557396, 0.9586763, 0.9667827, 0.9734911, 0.9673615, 
    0.9609221, 0.9426289, 0.9261296, 0.9081287, 0.9037223, 0.8826637, 
    0.8998045, 0.8715091, 0.8955626, 0.8539122, 0.928706, 0.8962744, 
    0.9550026, 0.9486834, 0.9372469, 0.9109995, 0.9251755, 0.9085971, 
    0.9451929, 0.9641544, 0.9690608, 0.9782075, 0.9688516, 0.9696128, 
    0.960657, 0.9635354, 0.9420213, 0.9535801, 0.9207289, 0.9087286, 
    0.8748105, 0.853993, 0.8327881, 0.8234196, 0.8205676, 0.8193752,
  0.4324116, 0.4167897, 0.41981, 0.4073347, 0.4142381, 0.4060945, 0.4292279, 
    0.416173, 0.4244899, 0.4309978, 0.3835423, 0.4067819, 0.3599938, 
    0.3743855, 0.3386776, 0.3622167, 0.3340116, 0.33935, 0.323397, 0.3279341, 
    0.3078829, 0.3213121, 0.2977086, 0.3110688, 0.308961, 0.3217589, 
    0.4020644, 0.3864053, 0.4029993, 0.4007495, 0.401759, 0.4140942, 
    0.420363, 0.4336163, 0.4311991, 0.4214715, 0.3997395, 0.4070683, 
    0.3887032, 0.3891143, 0.369056, 0.3780471, 0.3449826, 0.3542544, 
    0.3277443, 0.3343295, 0.3280519, 0.3299505, 0.3280272, 0.3377078, 
    0.3335455, 0.3421179, 0.3763561, 0.3661546, 0.3969093, 0.4158661, 
    0.4286516, 0.4378112, 0.4365118, 0.4340384, 0.4214148, 0.4096786, 
    0.4008203, 0.3949367, 0.3891734, 0.3719279, 0.3629336, 0.3431189, 
    0.3466629, 0.3406696, 0.3349878, 0.3255365, 0.3270845, 0.3229482, 
    0.3408287, 0.3288991, 0.3486879, 0.3432272, 0.3876036, 0.4050864, 
    0.4126006, 0.4192284, 0.4355136, 0.4242417, 0.4286716, 0.4181633, 
    0.4115369, 0.4148095, 0.3947763, 0.4025184, 0.3624033, 0.3794759, 
    0.3356484, 0.3459345, 0.3332026, 0.3396748, 0.3286166, 0.338562, 
    0.3214152, 0.317731, 0.3202465, 0.3106327, 0.3391168, 0.3280512, 
    0.4149009, 0.4143664, 0.4118807, 0.4228498, 0.4235249, 0.4336822, 
    0.4246406, 0.4208116, 0.4111547, 0.4054819, 0.4001183, 0.3884243, 
    0.375526, 0.357788, 0.3452637, 0.3369718, 0.3420469, 0.3375645, 
    0.3425765, 0.3449367, 0.3191088, 0.3335063, 0.3120077, 0.3131815, 
    0.3228498, 0.3130492, 0.4139914, 0.4170696, 0.4278216, 0.4193983, 
    0.4347939, 0.4261491, 0.4212076, 0.402354, 0.3982589, 0.3944735, 
    0.3870414, 0.3775847, 0.3612233, 0.3472307, 0.3346588, 0.3355735, 
    0.3352513, 0.3324665, 0.3393813, 0.3313371, 0.3299942, 0.333509, 
    0.3133388, 0.3190465, 0.3132065, 0.3169172, 0.4160683, 0.410899, 
    0.413689, 0.4084481, 0.4121369, 0.3958307, 0.3909921, 0.3686698, 
    0.3777695, 0.363332, 0.3762933, 0.3739827, 0.3628613, 0.3755887, 
    0.3479946, 0.3666056, 0.3323584, 0.350595, 0.3312291, 0.3347127, 
    0.3289541, 0.3238317, 0.3174378, 0.3057821, 0.3084647, 0.2988274, 
    0.4032401, 0.3966208, 0.3972035, 0.3903197, 0.385259, 0.374383, 0.357201, 
    0.3636241, 0.3518702, 0.3495292, 0.3674012, 0.3563832, 0.3922161, 
    0.386332, 0.3898323, 0.4027154, 0.3621376, 0.3827464, 0.345058, 
    0.3559496, 0.3245598, 0.3400175, 0.3099454, 0.2974532, 0.2859097, 
    0.2726704, 0.3930282, 0.397505, 0.3895047, 0.3785395, 0.3684827, 
    0.355281, 0.3539423, 0.3514944, 0.3451885, 0.3399224, 0.3507204, 
    0.3386077, 0.3849691, 0.3603714, 0.3992012, 0.3873398, 0.3791831, 
    0.3827544, 0.3643616, 0.3600797, 0.3428938, 0.3517355, 0.3005142, 
    0.322752, 0.262785, 0.2789902, 0.3990735, 0.3930444, 0.3723435, 
    0.3821375, 0.3544076, 0.3477127, 0.3423106, 0.3354538, 0.3347182, 
    0.3306871, 0.3373033, 0.330948, 0.3552531, 0.3443034, 0.3746889, 
    0.3671958, 0.3706359, 0.374423, 0.3627849, 0.3505489, 0.3502919, 
    0.3464059, 0.3355479, 0.354297, 0.29769, 0.3321514, 0.3865111, 0.3750742, 
    0.3734551, 0.3778609, 0.3483814, 0.3589494, 0.3307855, 0.3383031, 
    0.3260237, 0.3321013, 0.3329994, 0.3408841, 0.3458313, 0.3584615, 
    0.3688756, 0.3772209, 0.3752739, 0.3661302, 0.3498066, 0.3346505, 
    0.3379461, 0.3269502, 0.3563895, 0.343915, 0.3487138, 0.3362596, 
    0.3637949, 0.3402825, 0.369907, 0.3672697, 0.3591605, 0.3430738, 
    0.3395599, 0.3358201, 0.3381262, 0.3493967, 0.3512589, 0.3593574, 
    0.3616054, 0.3678434, 0.3730395, 0.3682902, 0.3633288, 0.349393, 
    0.3370266, 0.3237587, 0.3205473, 0.3053943, 0.3177021, 0.2975022, 
    0.3146342, 0.2852471, 0.3389437, 0.3151493, 0.3587942, 0.3539797, 
    0.3453372, 0.3258582, 0.3363178, 0.3241004, 0.3513322, 0.365815, 
    0.3696043, 0.3767109, 0.3694425, 0.3700317, 0.3631257, 0.3653393, 
    0.3489342, 0.3577079, 0.3330213, 0.3241968, 0.2998303, 0.285304, 
    0.2708519, 0.2645785, 0.2626826, 0.2618917,
  0.1957281, 0.1877837, 0.1893164, 0.1829964, 0.1864902, 0.1823697, 
    0.1941056, 0.187471, 0.1916943, 0.1950074, 0.1710214, 0.182717, 
    0.1592735, 0.1664407, 0.1487324, 0.160378, 0.146437, 0.1490635, 
    0.1412321, 0.143454, 0.1336675, 0.1402125, 0.1287349, 0.1352167, 
    0.1341915, 0.1404309, 0.1803349, 0.1724569, 0.1808066, 0.1796716, 
    0.1801808, 0.1864173, 0.1895972, 0.1963425, 0.19511, 0.1901602, 
    0.1791624, 0.1828618, 0.1736101, 0.1738165, 0.1637819, 0.1682705, 
    0.151841, 0.1564265, 0.1433609, 0.1465932, 0.1435118, 0.1444428, 
    0.1434996, 0.1482549, 0.1462079, 0.1504276, 0.1674251, 0.1623368, 
    0.1777364, 0.1873154, 0.1938121, 0.1984839, 0.1978203, 0.1965578, 
    0.1901314, 0.1841817, 0.1797073, 0.1767433, 0.1738462, 0.165214, 
    0.1607343, 0.1509213, 0.1526707, 0.1497136, 0.1469168, 0.1422793, 
    0.1430376, 0.1410125, 0.149792, 0.1439271, 0.1536714, 0.1509747, 
    0.1730581, 0.1818604, 0.1856608, 0.1890211, 0.1973107, 0.1915681, 
    0.1938223, 0.1884806, 0.1851221, 0.1867798, 0.1766626, 0.1805639, 
    0.1604707, 0.1689852, 0.1472417, 0.152311, 0.1460395, 0.1492235, 
    0.1437886, 0.1486754, 0.1402629, 0.1384634, 0.1396918, 0.1350045, 
    0.1489486, 0.1435114, 0.1868261, 0.1865552, 0.1852962, 0.1908605, 
    0.1912036, 0.1963761, 0.1917709, 0.1898249, 0.1849287, 0.1820602, 
    0.1793534, 0.1734701, 0.1670104, 0.1581786, 0.1519798, 0.1478927, 
    0.1503925, 0.1481844, 0.1506537, 0.1518183, 0.139136, 0.1461887, 
    0.1356737, 0.1362453, 0.1409644, 0.1361808, 0.1863652, 0.1879257, 
    0.1933895, 0.1891074, 0.1969434, 0.1925383, 0.1900261, 0.180481, 
    0.1784162, 0.1765103, 0.172776, 0.1680393, 0.1598842, 0.1529512, 
    0.1467551, 0.1472048, 0.1470464, 0.1456779, 0.1490789, 0.1451233, 
    0.1444643, 0.14619, 0.1363219, 0.1391056, 0.1362574, 0.1380663, 
    0.1874179, 0.1847993, 0.186212, 0.1835593, 0.1854259, 0.1771934, 
    0.1747598, 0.1635894, 0.1681317, 0.1609324, 0.1673937, 0.1662395, 
    0.1606984, 0.1670417, 0.1533288, 0.1625613, 0.1456248, 0.1546147, 
    0.1450703, 0.1467816, 0.1439541, 0.1414448, 0.1383203, 0.1326472, 
    0.1339502, 0.1292761, 0.1809282, 0.1775911, 0.1778846, 0.1744219, 
    0.1718819, 0.1664394, 0.1578874, 0.1610776, 0.1552457, 0.1540875, 
    0.1629574, 0.1574817, 0.175375, 0.1724201, 0.1741771, 0.1806634, 
    0.1603386, 0.1706226, 0.1518782, 0.1572667, 0.1418011, 0.1493923, 
    0.1346702, 0.1286113, 0.1230435, 0.1166953, 0.1757833, 0.1780364, 
    0.1740126, 0.1685168, 0.1634962, 0.1569353, 0.1562719, 0.1550597, 
    0.1519427, 0.1493454, 0.1546767, 0.1486979, 0.1717366, 0.1594611, 
    0.1788911, 0.1729257, 0.1688387, 0.1706266, 0.1614445, 0.1593162, 
    0.1508103, 0.155179, 0.1300928, 0.1409166, 0.1119821, 0.1197205, 
    0.1788267, 0.1757914, 0.1654213, 0.1703176, 0.1565024, 0.1531894, 
    0.1505226, 0.147146, 0.1467843, 0.1448043, 0.1480558, 0.1449323, 
    0.1569214, 0.1515057, 0.1665922, 0.1628551, 0.1645695, 0.1664594, 
    0.1606603, 0.1545918, 0.1544647, 0.1525438, 0.1471923, 0.1564476, 
    0.1287259, 0.1455232, 0.1725099, 0.1667846, 0.1659761, 0.1681774, 
    0.1535199, 0.158755, 0.1448526, 0.1485479, 0.1425179, 0.1454985, 
    0.1459396, 0.1498193, 0.15226, 0.1585128, 0.163692, 0.1678574, 0.1668844, 
    0.1623246, 0.1542247, 0.146751, 0.1483722, 0.1429718, 0.1574848, 
    0.151314, 0.1536842, 0.1475423, 0.1611626, 0.1495229, 0.1642061, 
    0.162892, 0.1588598, 0.1508991, 0.1491669, 0.1473261, 0.1484609, 
    0.1540219, 0.1549432, 0.1589575, 0.1600741, 0.1631777, 0.1657686, 
    0.1634003, 0.1609308, 0.1540201, 0.1479196, 0.1414091, 0.1398387, 
    0.1324589, 0.1384494, 0.1286351, 0.1369531, 0.1227248, 0.1488634, 
    0.1372042, 0.1586779, 0.1562904, 0.1520161, 0.1424368, 0.1475709, 
    0.1415763, 0.1549794, 0.1621677, 0.1640552, 0.1676024, 0.1639745, 
    0.1642682, 0.1608298, 0.1619309, 0.1537932, 0.1581388, 0.1459504, 
    0.1416235, 0.1297616, 0.1227522, 0.1158265, 0.1128355, 0.1119334, 
    0.1115574,
  0.04776575, 0.04543493, 0.0458828, 0.04404155, 0.0450576, 0.04385975, 
    0.04728786, 0.04534366, 0.04657938, 0.04755335, 0.04059398, 0.04396048, 
    0.03726594, 0.03928975, 0.03432754, 0.03757647, 0.0336939, 0.0344191, 
    0.03226544, 0.0328738, 0.03021061, 0.031987, 0.02888454, 0.03062934, 
    0.03035212, 0.03204662, 0.04327058, 0.04100436, 0.04340703, 0.04307887, 
    0.04322601, 0.04503635, 0.04596497, 0.04794696, 0.04758357, 0.04612975, 
    0.04293179, 0.04400246, 0.04133454, 0.04139371, 0.03853657, 0.03980972, 
    0.0351892, 0.03646773, 0.03284827, 0.03373694, 0.03288964, 0.03314522, 
    0.03288632, 0.03419553, 0.03363078, 0.03479691, 0.03956933, 0.03812838, 
    0.04252045, 0.04529829, 0.04720152, 0.04857958, 0.04838336, 0.0480105, 
    0.04612131, 0.04438572, 0.04308916, 0.04223444, 0.04140221, 0.03894195, 
    0.03767676, 0.03493385, 0.0354199, 0.03459908, 0.03382615, 0.03255191, 
    0.03275963, 0.03220546, 0.03462078, 0.03300362, 0.03569851, 0.03494866, 
    0.04117648, 0.04371214, 0.044816, 0.04579646, 0.04823278, 0.04654237, 
    0.04720452, 0.04563844, 0.04465919, 0.04514201, 0.04221121, 0.04333681, 
    0.03760255, 0.04001318, 0.03391576, 0.03531983, 0.03358438, 0.03446337, 
    0.0329656, 0.03431176, 0.03200077, 0.03151042, 0.03184498, 0.03057192, 
    0.03438732, 0.03288954, 0.04515552, 0.04507655, 0.04470984, 0.0463349, 
    0.04643549, 0.04795688, 0.04660186, 0.04603161, 0.0446029, 0.04377003, 
    0.04298692, 0.04129443, 0.03945151, 0.03695856, 0.03522776, 0.03409545, 
    0.03478719, 0.03417604, 0.03485962, 0.03518289, 0.03169354, 0.03362548, 
    0.03075306, 0.03090795, 0.03219231, 0.03089048, 0.04502116, 0.04547636, 
    0.04707724, 0.04582166, 0.0481243, 0.04682712, 0.0460905, 0.04331285, 
    0.04271644, 0.04216739, 0.04109562, 0.03974395, 0.03743757, 0.03549796, 
    0.03378155, 0.03390559, 0.03386188, 0.03348482, 0.03442337, 0.03333226, 
    0.03315113, 0.03362583, 0.03092873, 0.03168524, 0.03091125, 0.03140241, 
    0.04532814, 0.04456526, 0.04497653, 0.04420494, 0.04474761, 0.04236402, 
    0.04166434, 0.03848219, 0.03977023, 0.03773252, 0.03956041, 0.03923268, 
    0.03766666, 0.03946038, 0.03560308, 0.03819177, 0.03347022, 0.03596156, 
    0.03331768, 0.03378887, 0.03301102, 0.0323236, 0.03147149, 0.02993538, 
    0.03028693, 0.0290295, 0.0434422, 0.04247859, 0.04256314, 0.04156736, 
    0.04083983, 0.03928938, 0.03687689, 0.03777341, 0.03613768, 0.03581447, 
    0.03830359, 0.0367632, 0.04184099, 0.04099378, 0.04149713, 0.04336559, 
    0.03756538, 0.04048007, 0.03519954, 0.03670296, 0.03242105, 0.03451012, 
    0.03048149, 0.02885149, 0.02736846, 0.02569561, 0.04195831, 0.04260692, 
    0.04144993, 0.03987982, 0.03845581, 0.03661013, 0.03642448, 0.03608574, 
    0.03521744, 0.03449712, 0.03597884, 0.03431799, 0.04079833, 0.03731861, 
    0.04285346, 0.04113852, 0.03997147, 0.04048119, 0.03787675, 0.03727789, 
    0.03490304, 0.03611906, 0.0292485, 0.03217926, 0.02446634, 0.0264904, 
    0.04283487, 0.04196064, 0.03900067, 0.040393, 0.03648897, 0.03556427, 
    0.03482324, 0.03388936, 0.03378961, 0.03324455, 0.03414052, 0.03327974, 
    0.03660626, 0.03509607, 0.03933274, 0.03827471, 0.03875938, 0.03929505, 
    0.0376559, 0.03595517, 0.03591968, 0.0353846, 0.0339022, 0.03647365, 
    0.02888218, 0.03344232, 0.04101946, 0.03938741, 0.03915794, 0.03978322, 
    0.03565631, 0.03712029, 0.03325782, 0.03427651, 0.03261724, 0.03343548, 
    0.03355688, 0.03462835, 0.03530567, 0.03705232, 0.03851116, 0.03969221, 
    0.03941571, 0.03812495, 0.03585275, 0.03378044, 0.03422796, 0.03274159, 
    0.03676406, 0.03504285, 0.0357021, 0.03399872, 0.03779734, 0.03454631, 
    0.03865653, 0.0382851, 0.03714971, 0.03492769, 0.0344477, 0.03393906, 
    0.03425245, 0.03579622, 0.03605321, 0.03717715, 0.03749096, 0.03836581, 
    0.0390991, 0.03842871, 0.03773206, 0.0357957, 0.03410292, 0.03231383, 
    0.03188505, 0.02988469, 0.03150662, 0.02885787, 0.03110005, 0.02728408, 
    0.03436378, 0.03116817, 0.03709865, 0.03642966, 0.03523786, 0.03259506, 
    0.03400661, 0.03235957, 0.03606332, 0.0380807, 0.03861386, 0.03961973, 
    0.03859104, 0.03867412, 0.03770361, 0.0380139, 0.03573246, 0.0369474, 
    0.03355985, 0.03237246, 0.02915963, 0.02729129, 0.02546818, 0.02468809, 
    0.02445369, 0.0243561,
  0.004169275, 0.003916436, 0.003964748, 0.003766965, 0.003875833, 
    0.003747558, 0.004117152, 0.003906607, 0.004040147, 0.00414609, 
    0.003402713, 0.003758308, 0.003058915, 0.003267038, 0.002762104, 
    0.003090658, 0.00269896, 0.002771252, 0.002557761, 0.002617697, 
    0.002357529, 0.002530428, 0.002230166, 0.00239805, 0.002371206, 
    0.002536275, 0.003684809, 0.003445647, 0.003699321, 0.003664444, 
    0.003680073, 0.00387355, 0.00397363, 0.004189074, 0.004149387, 
    0.003991444, 0.003648835, 0.003762788, 0.003480267, 0.003486481, 
    0.003189238, 0.003320982, 0.002848464, 0.002977645, 0.002615177, 
    0.002703237, 0.002619263, 0.002644533, 0.002618934, 0.002748921, 
    0.002692685, 0.002809075, 0.00329602, 0.003147244, 0.003605258, 
    0.003901726, 0.004107751, 0.004258366, 0.004236847, 0.004196024, 
    0.003990531, 0.003803765, 0.003665535, 0.003575026, 0.003487374, 
    0.003231065, 0.003100923, 0.002822813, 0.002871683, 0.002789258, 
    0.002712112, 0.002585948, 0.002606428, 0.002551869, 0.002791429, 
    0.002630527, 0.002899776, 0.002824299, 0.00346369, 0.003731813, 
    0.003849888, 0.003955425, 0.00422035, 0.004036134, 0.004108078, 
    0.003938372, 0.003833062, 0.003884906, 0.003572573, 0.003691852, 
    0.003093326, 0.003342144, 0.002721032, 0.002861607, 0.002688075, 
    0.002775678, 0.002626768, 0.002760526, 0.002531778, 0.002483789, 
    0.002516511, 0.002392483, 0.002768075, 0.002619254, 0.00388636, 
    0.003877869, 0.003838493, 0.00401365, 0.004024548, 0.004190159, 
    0.004042585, 0.00398083, 0.003827028, 0.003737985, 0.003654683, 
    0.003476057, 0.0032838, 0.003027564, 0.002852343, 0.002738938, 0.0028081, 
    0.002746976, 0.002815364, 0.002847829, 0.002501688, 0.002692159, 
    0.00241005, 0.002425092, 0.002550577, 0.002423394, 0.003871916, 
    0.003920898, 0.004094226, 0.003958145, 0.004208473, 0.004067038, 
    0.003987199, 0.003689305, 0.003626005, 0.003567947, 0.003455203, 
    0.003314148, 0.003076449, 0.00287955, 0.002707674, 0.002720018, 
    0.002715667, 0.002678192, 0.002771678, 0.002663059, 0.002645118, 
    0.002692193, 0.002427111, 0.002500875, 0.002425413, 0.002473242, 
    0.003904933, 0.003822994, 0.00386712, 0.003784425, 0.003842546, 
    0.003588718, 0.003514934, 0.003183638, 0.003316879, 0.003106633, 
    0.003295093, 0.003261128, 0.003099891, 0.003284718, 0.00289015, 
    0.00315376, 0.002676743, 0.00292636, 0.002661614, 0.002708402, 
    0.002631257, 0.002563479, 0.002479986, 0.002330971, 0.002364902, 
    0.002244015, 0.003703062, 0.00360083, 0.003609774, 0.00350473, 
    0.003428413, 0.003266999, 0.003019244, 0.003110822, 0.00294418, 
    0.002911488, 0.003165253, 0.003007674, 0.003533529, 0.003444534, 
    0.003497348, 0.003694912, 0.003089522, 0.003390811, 0.002849504, 
    0.003001546, 0.002573064, 0.002780356, 0.002383725, 0.002227013, 
    0.002086404, 0.001930147, 0.003545891, 0.003614408, 0.003492387, 
    0.003328272, 0.00318092, 0.00299211, 0.002973255, 0.002938922, 
    0.002851304, 0.002779054, 0.002928105, 0.002761147, 0.003424076, 
    0.003064293, 0.003640528, 0.003459704, 0.003337804, 0.003390926, 
    0.003121415, 0.003060132, 0.002819721, 0.002942294, 0.002264977, 
    0.002549296, 0.001816958, 0.002004071, 0.003638556, 0.003546136, 
    0.00323713, 0.003381722, 0.002979802, 0.002886233, 0.002811715, 
    0.002718404, 0.002708476, 0.002654369, 0.002743432, 0.002657855, 
    0.002991716, 0.002839102, 0.00327149, 0.003162284, 0.003212209, 
    0.003267585, 0.003098785, 0.002925711, 0.002922121, 0.002868128, 
    0.002719689, 0.002978246, 0.002229947, 0.00267398, 0.003447222, 
    0.003277157, 0.003253393, 0.003318228, 0.002895519, 0.003044049, 
    0.002655683, 0.002757005, 0.002592385, 0.002673295, 0.002685345, 
    0.002792187, 0.002860181, 0.003037118, 0.00318662, 0.003308773, 
    0.003280087, 0.003146892, 0.002915357, 0.002707564, 0.002752159, 
    0.002604647, 0.00300776, 0.002833757, 0.002900141, 0.002729296, 
    0.003113274, 0.002783982, 0.003201601, 0.003163351, 0.00304705, 
    0.002822196, 0.002774111, 0.002723353, 0.002754602, 0.002909645, 
    0.002935629, 0.003049849, 0.003081907, 0.003171654, 0.003247305, 
    0.003178129, 0.003106586, 0.002909591, 0.002739683, 0.002562518, 
    0.002520435, 0.00232609, 0.00248342, 0.002227626, 0.002443783, 
    0.002078467, 0.002765727, 0.002450412, 0.003041841, 0.002973781, 
    0.00285336, 0.002590202, 0.002730082, 0.002567017, 0.002936652, 
    0.003142348, 0.003197202, 0.003301249, 0.00319485, 0.003203415, 
    0.003103671, 0.003135486, 0.002903205, 0.003026425, 0.00268564, 
    0.002568285, 0.002256465, 0.002079142, 0.001909097, 0.00183727, 
    0.0018158, 0.001806877,
  0.000114897, 0.000106181, 0.0001078352, 0.0001010979, 0.000104795, 
    0.0001004417, 0.0001130883, 0.0001058452, 0.0001104275, 0.0001140917, 
    8.893685e-05, 0.000100805, 7.777032e-05, 8.449257e-05, 6.83921e-05, 
    7.878805e-05, 6.643006e-05, 6.867729e-05, 6.208653e-05, 6.392276e-05, 
    5.603503e-05, 6.125286e-05, 5.225461e-05, 5.724916e-05, 5.644422e-05, 
    6.143101e-05, 9.832645e-05, 9.035307e-05, 9.881479e-05, 9.7642e-05, 
    9.816718e-05, 0.0001047172, 0.0001081399, 0.0001155855, 0.0001142061, 
    0.0001087516, 9.711811e-05, 0.0001009565, 9.149825e-05, 9.170413e-05, 
    8.1966e-05, 8.625379e-05, 7.109458e-05, 7.517746e-05, 6.384531e-05, 
    6.656255e-05, 6.397087e-05, 6.47485e-05, 6.396078e-05, 6.798145e-05, 
    6.623571e-05, 6.985923e-05, 8.543784e-05, 8.060901e-05, 9.565856e-05, 
    0.0001056786, 0.0001127628, 0.0001180023, 0.0001172506, 0.0001158275, 
    0.0001087202, 0.0001023444, 9.76786e-05, 9.464868e-05, 9.173375e-05, 
    8.332247e-05, 7.911772e-05, 7.028961e-05, 7.182488e-05, 6.923944e-05, 
    6.683768e-05, 6.29487e-05, 6.357664e-05, 6.190663e-05, 6.930727e-05, 
    6.431728e-05, 7.271061e-05, 7.033613e-05, 9.094964e-05, 9.991003e-05, 
    0.0001039115, 0.0001075156, 0.0001166751, 0.0001102892, 0.0001127741, 
    0.0001069314, 0.0001033391, 0.0001051044, 9.456686e-05, 9.856335e-05, 
    7.887368e-05, 8.694681e-05, 6.711447e-05, 7.150776e-05, 6.609302e-05, 
    6.881535e-05, 6.420165e-05, 6.834284e-05, 6.129399e-05, 5.983587e-05, 
    6.082932e-05, 5.7082e-05, 6.857818e-05, 6.397061e-05, 0.000105154, 
    0.0001048644, 0.0001035238, 0.0001095151, 0.0001098901, 0.0001156233, 
    0.0001105115, 0.000108387, 0.0001031341, 0.0001001184, 9.731428e-05, 
    9.135883e-05, 8.503905e-05, 7.676791e-05, 7.121645e-05, 6.767081e-05, 
    6.982867e-05, 6.792087e-05, 7.005614e-05, 7.107459e-05, 6.037889e-05, 
    6.621942e-05, 5.760973e-05, 5.80624e-05, 6.186723e-05, 5.801126e-05, 
    0.0001046615, 0.0001063336, 0.0001122948, 0.0001076087, 0.0001162611, 
    0.0001113552, 0.0001086058, 9.847771e-05, 9.635282e-05, 9.441259e-05, 
    9.066873e-05, 8.603025e-05, 7.833209e-05, 7.20727e-05, 6.670006e-05, 
    6.7083e-05, 6.694798e-05, 6.578732e-05, 6.869056e-05, 6.531987e-05, 
    6.476657e-05, 6.622048e-05, 5.812322e-05, 6.035417e-05, 5.807205e-05, 
    5.951637e-05, 0.0001057879, 0.0001029971, 0.0001044981, 0.0001016888, 
    0.0001036616, 9.510584e-05, 9.26483e-05, 8.178482e-05, 8.611958e-05, 
    7.930122e-05, 8.540757e-05, 8.43001e-05, 7.908461e-05, 8.506893e-05, 
    7.240693e-05, 8.081932e-05, 6.574253e-05, 7.355095e-05, 6.527526e-05, 
    6.672261e-05, 6.433971e-05, 6.226123e-05, 5.972062e-05, 5.524218e-05, 
    5.62555e-05, 5.266298e-05, 9.894076e-05, 9.551053e-05, 9.580955e-05, 
    9.230942e-05, 8.978385e-05, 8.449126e-05, 7.650234e-05, 7.943584e-05, 
    7.411517e-05, 7.308053e-05, 8.119032e-05, 7.613337e-05, 9.326632e-05, 
    9.031619e-05, 9.20645e-05, 9.86664e-05, 7.875152e-05, 8.854497e-05, 
    7.112725e-05, 7.593808e-05, 6.255431e-05, 6.89614e-05, 5.681928e-05, 
    5.216175e-05, 4.805496e-05, 4.357558e-05, 9.367769e-05, 9.596458e-05, 
    9.189993e-05, 8.649244e-05, 8.169683e-05, 7.56376e-05, 7.503793e-05, 
    7.394858e-05, 7.118379e-05, 6.892071e-05, 7.360611e-05, 6.836221e-05, 
    8.964092e-05, 7.794252e-05, 9.683947e-05, 9.081766e-05, 8.68046e-05, 
    8.85487e-05, 7.977666e-05, 7.780921e-05, 7.01927e-05, 7.40554e-05, 
    5.328243e-05, 6.182817e-05, 4.038892e-05, 4.568341e-05, 9.677334e-05, 
    9.368582e-05, 8.351941e-05, 8.824596e-05, 7.524603e-05, 7.228335e-05, 
    6.994186e-05, 6.703293e-05, 6.672492e-05, 6.505174e-05, 6.781062e-05, 
    6.515926e-05, 7.562508e-05, 7.080054e-05, 8.463758e-05, 8.109443e-05, 
    8.271029e-05, 8.451035e-05, 7.904894e-05, 7.353036e-05, 7.34167e-05, 
    7.1713e-05, 6.707299e-05, 7.519655e-05, 5.224829e-05, 6.565732e-05, 
    9.040489e-05, 8.482242e-05, 8.404826e-05, 8.616365e-05, 7.257625e-05, 
    7.729462e-05, 6.509225e-05, 6.823314e-05, 6.314592e-05, 6.563597e-05, 
    6.600854e-05, 6.933093e-05, 7.146293e-05, 7.707309e-05, 8.188127e-05, 
    8.585449e-05, 8.491787e-05, 8.059762e-05, 7.320285e-05, 6.669668e-05, 
    6.808227e-05, 6.352199e-05, 7.613609e-05, 7.063281e-05, 7.272215e-05, 
    6.737112e-05, 7.951473e-05, 6.907476e-05, 8.236639e-05, 8.11289e-05, 
    7.739059e-05, 7.027028e-05, 6.876647e-05, 6.718656e-05, 6.81583e-05, 
    7.302232e-05, 7.384427e-05, 7.748009e-05, 7.850715e-05, 8.139718e-05, 
    8.385019e-05, 8.160653e-05, 7.929969e-05, 7.302059e-05, 6.769402e-05, 
    6.223189e-05, 6.094867e-05, 5.50968e-05, 5.982476e-05, 5.217993e-05, 
    5.862611e-05, 4.782535e-05, 6.850507e-05, 5.882615e-05, 7.7224e-05, 
    7.505462e-05, 7.12485e-05, 6.307909e-05, 6.739556e-05, 6.236944e-05, 
    7.387669e-05, 8.045111e-05, 8.222385e-05, 8.560863e-05, 8.214769e-05, 
    8.242516e-05, 7.920592e-05, 8.022983e-05, 7.281887e-05, 7.673149e-05, 
    6.60177e-05, 6.240817e-05, 5.303068e-05, 4.784483e-05, 4.297911e-05, 
    4.095705e-05, 4.035656e-05, 4.010754e-05,
  8.832795e-07, 7.95726e-07, 8.121857e-07, 7.456201e-07, 7.819916e-07, 
    7.392054e-07, 8.649455e-07, 7.923937e-07, 8.381294e-07, 8.751055e-07, 
    6.288043e-07, 7.427559e-07, 5.256611e-07, 5.872552e-07, 4.424229e-07, 
    5.348868e-07, 4.254318e-07, 4.449047e-07, 3.883713e-07, 4.039435e-07, 
    3.380807e-07, 3.813481e-07, 3.075086e-07, 3.480399e-07, 3.414296e-07, 
    3.828465e-07, 7.186105e-07, 6.421767e-07, 7.233536e-07, 7.119747e-07, 
    7.170651e-07, 7.812225e-07, 8.152271e-07, 8.902805e-07, 8.762659e-07, 
    8.213364e-07, 7.069048e-07, 7.442366e-07, 6.530337e-07, 6.549902e-07, 
    5.639245e-07, 6.036433e-07, 4.660714e-07, 5.023229e-07, 4.032839e-07, 
    4.265739e-07, 4.043535e-07, 4.10992e-07, 4.042676e-07, 4.388537e-07, 
    4.237568e-07, 4.55226e-07, 5.960385e-07, 5.514827e-07, 6.928223e-07, 
    7.907419e-07, 8.616549e-07, 9.14952e-07, 9.072628e-07, 8.927443e-07, 
    8.210231e-07, 7.578399e-07, 7.123287e-07, 6.831155e-07, 6.552718e-07, 
    5.764248e-07, 5.378826e-07, 4.589981e-07, 4.7251e-07, 4.498072e-07, 
    4.289488e-07, 3.956655e-07, 4.009976e-07, 3.868534e-07, 4.503992e-07, 
    4.073079e-07, 4.803458e-07, 4.594059e-07, 6.478286e-07, 7.340163e-07, 
    7.732659e-07, 8.089996e-07, 9.01385e-07, 8.367414e-07, 8.617695e-07, 
    8.031828e-07, 7.676232e-07, 7.850524e-07, 6.823303e-07, 7.209105e-07, 
    5.356644e-07, 6.101201e-07, 4.31341e-07, 4.697117e-07, 4.22528e-07, 
    4.461074e-07, 4.063211e-07, 4.419939e-07, 3.816941e-07, 3.694796e-07, 
    3.777917e-07, 3.466645e-07, 4.440416e-07, 4.043515e-07, 7.855435e-07, 
    7.826781e-07, 7.694418e-07, 8.289776e-07, 8.327369e-07, 8.906653e-07, 
    8.389736e-07, 8.176934e-07, 7.656038e-07, 7.360484e-07, 7.088019e-07, 
    6.517097e-07, 5.923296e-07, 5.166099e-07, 4.671444e-07, 4.361583e-07, 
    4.549584e-07, 4.383276e-07, 4.569507e-07, 4.658952e-07, 3.740177e-07, 
    4.236166e-07, 3.510104e-07, 3.547481e-07, 3.865211e-07, 3.543254e-07, 
    7.806715e-07, 7.972401e-07, 8.569286e-07, 8.099277e-07, 8.97162e-07, 
    8.474577e-07, 8.198793e-07, 7.200793e-07, 6.995125e-07, 6.808509e-07, 
    6.45164e-07, 6.015577e-07, 5.307486e-07, 4.746996e-07, 4.277605e-07, 
    4.310688e-07, 4.299015e-07, 4.198988e-07, 4.450202e-07, 4.158855e-07, 
    4.111467e-07, 4.236255e-07, 3.552509e-07, 3.738106e-07, 3.548278e-07, 
    3.668152e-07, 7.91825e-07, 7.642556e-07, 7.790562e-07, 7.514079e-07, 
    7.708008e-07, 6.875063e-07, 6.639806e-07, 5.622601e-07, 6.023911e-07, 
    5.395518e-07, 5.957565e-07, 5.854704e-07, 5.375821e-07, 5.926069e-07, 
    4.776565e-07, 5.534075e-07, 4.195139e-07, 4.878082e-07, 4.15503e-07, 
    4.279551e-07, 4.074991e-07, 3.898468e-07, 3.685178e-07, 3.31613e-07, 
    3.398837e-07, 3.107781e-07, 7.245779e-07, 6.913976e-07, 6.942757e-07, 
    6.607501e-07, 6.367927e-07, 5.872429e-07, 5.142179e-07, 5.407768e-07, 
    4.928316e-07, 4.836273e-07, 5.568045e-07, 5.108992e-07, 6.69879e-07, 
    6.418264e-07, 6.584183e-07, 7.219117e-07, 5.345547e-07, 6.251141e-07, 
    4.66359e-07, 5.091442e-07, 3.923251e-07, 4.473811e-07, 3.445058e-07, 
    3.067665e-07, 2.743633e-07, 2.400246e-07, 6.738118e-07, 6.957692e-07, 
    6.568521e-07, 6.058724e-07, 5.614515e-07, 5.064471e-07, 5.010739e-07, 
    4.91347e-07, 4.668566e-07, 4.470259e-07, 4.882984e-07, 4.421622e-07, 
    6.354442e-07, 5.272192e-07, 7.042112e-07, 6.46576e-07, 6.087898e-07, 
    6.251487e-07, 5.438819e-07, 5.260123e-07, 4.581481e-07, 4.922988e-07, 
    3.157537e-07, 3.861921e-07, 2.162781e-07, 2.56048e-07, 7.03572e-07, 
    6.738895e-07, 5.782438e-07, 6.223021e-07, 5.02937e-07, 4.765624e-07, 
    4.559495e-07, 4.306361e-07, 4.27975e-07, 4.135875e-07, 4.373709e-07, 
    4.145085e-07, 5.063348e-07, 4.634846e-07, 5.886004e-07, 5.55926e-07, 
    5.707748e-07, 5.874198e-07, 5.372565e-07, 4.876247e-07, 4.866135e-07, 
    4.715224e-07, 4.309839e-07, 5.024938e-07, 3.074591e-07, 4.187832e-07, 
    6.426652e-07, 5.903173e-07, 5.831369e-07, 6.028021e-07, 4.791555e-07, 
    5.213609e-07, 4.139344e-07, 4.410401e-07, 3.973383e-07, 4.185983e-07, 
    4.218012e-07, 4.506059e-07, 4.693163e-07, 5.193615e-07, 5.631458e-07, 
    5.999187e-07, 5.91203e-07, 5.513784e-07, 4.847137e-07, 4.277315e-07, 
    4.397294e-07, 4.005328e-07, 5.109231e-07, 4.620107e-07, 4.804485e-07, 
    4.335618e-07, 5.414952e-07, 4.48371e-07, 5.676071e-07, 5.562416e-07, 
    5.222278e-07, 4.588288e-07, 4.456814e-07, 4.319646e-07, 4.403896e-07, 
    4.831108e-07, 4.90418e-07, 5.230363e-07, 5.323361e-07, 5.587012e-07, 
    5.813028e-07, 5.606223e-07, 5.395377e-07, 4.830953e-07, 4.363598e-07, 
    3.895991e-07, 3.787929e-07, 3.304309e-07, 3.693874e-07, 3.069127e-07, 
    3.594172e-07, 2.72578e-07, 4.434061e-07, 3.61076e-07, 5.207232e-07, 
    5.012233e-07, 4.674271e-07, 3.967719e-07, 4.337734e-07, 3.907618e-07, 
    4.907067e-07, 5.500393e-07, 5.662954e-07, 5.976283e-07, 5.655947e-07, 
    5.681482e-07, 5.386842e-07, 5.480169e-07, 4.813057e-07, 5.162814e-07, 
    4.2188e-07, 3.910892e-07, 3.137291e-07, 2.727289e-07, 2.35535e-07, 
    2.204682e-07, 2.160399e-07, 2.142099e-07,
  1.067067e-09, 8.8233e-10, 9.162233e-10, 7.816657e-10, 8.543553e-10, 
    7.690595e-10, 1.027492e-09, 8.755178e-10, 9.704454e-10, 1.049366e-09, 
    5.628623e-10, 7.760288e-10, 3.906317e-10, 4.909234e-10, 2.684904e-10, 
    4.051466e-10, 2.45648e-10, 2.718884e-10, 1.985203e-10, 2.178594e-10, 
    1.40961e-10, 1.90025e-10, 1.09916e-10, 1.517393e-10, 1.445497e-10, 
    1.918255e-10, 7.290314e-10, 5.867045e-10, 7.381892e-10, 7.162822e-10, 
    7.260557e-10, 8.527981e-10, 9.225318e-10, 1.082297e-09, 1.051873e-09, 
    9.352384e-10, 7.0659e-10, 7.7894e-10, 6.062957e-10, 6.098497e-10, 
    4.52011e-10, 5.189008e-10, 3.015066e-10, 3.547519e-10, 2.170263e-10, 
    2.471589e-10, 2.183779e-10, 2.268356e-10, 2.182692e-10, 2.63629e-10, 
    2.434365e-10, 2.861911e-10, 5.05853e-10, 4.31714e-10, 6.79892e-10, 
    8.721489e-10, 1.020439e-09, 1.136492e-09, 1.119516e-09, 1.087674e-09, 
    9.345854e-10, 8.058578e-10, 7.169592e-10, 6.616841e-10, 6.103619e-10, 
    4.727263e-10, 4.098988e-10, 2.914856e-10, 3.107352e-10, 2.78649e-10, 
    2.503133e-10, 2.074939e-10, 2.141486e-10, 1.966725e-10, 2.794688e-10, 
    2.221275e-10, 3.221011e-10, 2.920594e-10, 5.968799e-10, 7.589087e-10, 
    8.367338e-10, 9.096318e-10, 1.106591e-09, 9.67521e-10, 1.020685e-09, 
    8.976344e-10, 8.253953e-10, 8.605643e-10, 6.602184e-10, 7.334672e-10, 
    4.063777e-10, 5.301021e-10, 2.535059e-10, 3.067119e-10, 2.418193e-10, 
    2.735408e-10, 2.208724e-10, 2.679032e-10, 1.904403e-10, 1.75998e-10, 
    1.857783e-10, 1.502313e-10, 2.707043e-10, 2.183756e-10, 8.615624e-10, 
    8.557466e-10, 8.290429e-10, 9.512089e-10, 9.590962e-10, 1.083136e-09, 
    9.722259e-10, 9.276536e-10, 8.213498e-10, 7.628783e-10, 7.102108e-10, 
    6.038951e-10, 4.99531e-10, 3.765723e-10, 3.030376e-10, 2.599798e-10, 
    2.858166e-10, 2.62915e-10, 2.886071e-10, 3.012551e-10, 1.813124e-10, 
    2.432521e-10, 1.550149e-10, 1.591762e-10, 1.962689e-10, 1.587034e-10, 
    8.516815e-10, 8.854297e-10, 1.010333e-09, 9.115493e-10, 1.097333e-09, 
    9.901765e-10, 9.322032e-10, 7.318645e-10, 6.925329e-10, 6.5746e-10, 
    5.920702e-10, 5.153112e-10, 3.98612e-10, 3.138971e-10, 2.487328e-10, 
    2.531415e-10, 2.515828e-10, 2.383729e-10, 2.720468e-10, 2.331478e-10, 
    2.270347e-10, 2.432634e-10, 1.597395e-10, 1.81068e-10, 1.592655e-10, 
    1.729062e-10, 8.743545e-10, 8.186533e-10, 8.484131e-10, 7.930946e-10, 
    8.317732e-10, 6.69902e-10, 6.262703e-10, 4.492785e-10, 5.16745e-10, 
    4.125545e-10, 5.053711e-10, 4.87908e-10, 4.094225e-10, 5.000013e-10, 
    3.181852e-10, 4.348344e-10, 2.378698e-10, 3.330639e-10, 2.326521e-10, 
    2.489915e-10, 2.223702e-10, 2.003235e-10, 1.748792e-10, 1.34132e-10, 
    1.42888e-10, 1.130837e-10, 7.405586e-10, 6.7721e-10, 6.826311e-10, 
    6.203522e-10, 5.770612e-10, 4.909017e-10, 3.728867e-10, 4.145068e-10, 
    3.405132e-10, 3.269049e-10, 4.403556e-10, 3.677954e-10, 6.371182e-10, 
    5.860727e-10, 6.160939e-10, 7.354017e-10, 4.046199e-10, 5.563378e-10, 
    3.019168e-10, 3.651123e-10, 2.033657e-10, 2.752963e-10, 1.478778e-10, 
    1.092027e-10, 7.997167e-11, 5.34024e-11, 6.443853e-10, 6.854501e-10, 
    6.132382e-10, 5.227478e-10, 4.479511e-10, 3.610035e-10, 3.528663e-10, 
    3.383051e-10, 3.026263e-10, 2.748055e-10, 3.337871e-10, 2.68133e-10, 
    5.74659e-10, 3.930692e-10, 7.014572e-10, 5.946166e-10, 5.27795e-10, 
    5.563976e-10, 4.19472e-10, 3.911792e-10, 2.902895e-10, 3.397199e-10, 
    1.179772e-10, 1.958702e-10, 3.79132e-11, 6.520941e-11, 7.002402e-10, 
    6.445285e-10, 4.757644e-10, 5.51384e-10, 3.556802e-10, 3.165953e-10, 
    2.872034e-10, 2.525639e-10, 2.49018e-10, 2.301757e-10, 2.61619e-10, 
    2.31365e-10, 3.608328e-10, 2.978272e-10, 4.931991e-10, 4.389255e-10, 
    4.633218e-10, 4.912009e-10, 4.089021e-10, 3.327916e-10, 3.31298e-10, 
    3.093137e-10, 2.53032e-10, 3.550101e-10, 1.098702e-10, 2.369192e-10, 
    5.875764e-10, 4.961122e-10, 4.839748e-10, 5.174515e-10, 3.203655e-10, 
    3.839286e-10, 2.306234e-10, 2.666022e-10, 2.095728e-10, 2.366749e-10, 
    2.408647e-10, 2.797554e-10, 3.061451e-10, 3.808267e-10, 4.507313e-10, 
    5.124958e-10, 4.976142e-10, 4.31545e-10, 3.285017e-10, 2.486949e-10, 
    2.648189e-10, 2.135652e-10, 3.678314e-10, 2.957387e-10, 3.222521e-10, 
    2.564829e-10, 4.156543e-10, 2.76665e-10, 4.580793e-10, 4.394388e-10, 
    3.852763e-10, 2.912478e-10, 2.72955e-10, 2.543408e-10, 2.657163e-10, 
    3.261478e-10, 3.369259e-10, 3.865345e-10, 4.011136e-10, 4.4345e-10, 
    4.80891e-10, 4.465923e-10, 4.125318e-10, 3.261246e-10, 2.602525e-10, 
    2.000205e-10, 1.869699e-10, 1.329001e-10, 1.758917e-10, 1.093446e-10, 
    1.644391e-10, 7.847639e-11, 2.698358e-10, 1.663222e-10, 3.829377e-10, 
    3.530915e-10, 3.034423e-10, 2.088691e-10, 2.567673e-10, 2.014453e-10, 
    3.373541e-10, 4.293806e-10, 4.559146e-10, 5.085709e-10, 4.547596e-10, 
    4.589734e-10, 4.111718e-10, 4.261163e-10, 3.235041e-10, 3.760643e-10, 
    2.409685e-10, 2.018468e-10, 1.159754e-10, 7.860156e-11, 5.028594e-11, 
    4.046581e-11, 3.777032e-11, 3.668217e-11,
  4.050189e-13, 4.042921e-13, 4.044255e-13, 4.038955e-13, 4.041819e-13, 
    4.038458e-13, 4.048633e-13, 4.042653e-13, 4.046389e-13, 4.049493e-13, 
    4.030321e-13, 4.038733e-13, 4.023507e-13, 4.027477e-13, 4.018664e-13, 
    4.024082e-13, 4.017757e-13, 4.018799e-13, 4.015883e-13, 4.016652e-13, 
    4.013592e-13, 4.015545e-13, 4.012354e-13, 4.014021e-13, 4.013735e-13, 
    4.015617e-13, 4.03688e-13, 4.031263e-13, 4.037241e-13, 4.036377e-13, 
    4.036763e-13, 4.041758e-13, 4.044503e-13, 4.050787e-13, 4.049592e-13, 
    4.045004e-13, 4.035995e-13, 4.038848e-13, 4.032037e-13, 4.032177e-13, 
    4.025938e-13, 4.028583e-13, 4.019974e-13, 4.022085e-13, 4.016619e-13, 
    4.017817e-13, 4.016673e-13, 4.017009e-13, 4.016669e-13, 4.018471e-13, 
    4.017669e-13, 4.019366e-13, 4.028067e-13, 4.025134e-13, 4.034942e-13, 
    4.04252e-13, 4.048355e-13, 4.052917e-13, 4.05225e-13, 4.050999e-13, 
    4.044978e-13, 4.039909e-13, 4.036404e-13, 4.034223e-13, 4.032197e-13, 
    4.026757e-13, 4.02427e-13, 4.019577e-13, 4.02034e-13, 4.019067e-13, 
    4.017942e-13, 4.01624e-13, 4.016505e-13, 4.01581e-13, 4.0191e-13, 
    4.016822e-13, 4.020791e-13, 4.019599e-13, 4.031665e-13, 4.038058e-13, 
    4.041125e-13, 4.043996e-13, 4.051742e-13, 4.046274e-13, 4.048365e-13, 
    4.043523e-13, 4.040678e-13, 4.042064e-13, 4.034166e-13, 4.037055e-13, 
    4.024131e-13, 4.029026e-13, 4.018069e-13, 4.020181e-13, 4.017604e-13, 
    4.018864e-13, 4.016772e-13, 4.01864e-13, 4.015562e-13, 4.014987e-13, 
    4.015376e-13, 4.013961e-13, 4.018752e-13, 4.016673e-13, 4.042103e-13, 
    4.041874e-13, 4.040822e-13, 4.045632e-13, 4.045942e-13, 4.050821e-13, 
    4.046459e-13, 4.044705e-13, 4.040519e-13, 4.038215e-13, 4.036138e-13, 
    4.031942e-13, 4.027818e-13, 4.02295e-13, 4.020035e-13, 4.018326e-13, 
    4.019352e-13, 4.018442e-13, 4.019462e-13, 4.019964e-13, 4.015199e-13, 
    4.017661e-13, 4.014152e-13, 4.014318e-13, 4.015794e-13, 4.014299e-13, 
    4.041714e-13, 4.043043e-13, 4.047958e-13, 4.044071e-13, 4.051378e-13, 
    4.047165e-13, 4.044884e-13, 4.036992e-13, 4.035441e-13, 4.034057e-13, 
    4.031475e-13, 4.028442e-13, 4.023823e-13, 4.020466e-13, 4.017879e-13, 
    4.018054e-13, 4.017992e-13, 4.017468e-13, 4.018805e-13, 4.01726e-13, 
    4.017017e-13, 4.017662e-13, 4.01434e-13, 4.015189e-13, 4.014321e-13, 
    4.014864e-13, 4.042607e-13, 4.040413e-13, 4.041585e-13, 4.039406e-13, 
    4.04093e-13, 4.034548e-13, 4.032826e-13, 4.025829e-13, 4.028498e-13, 
    4.024376e-13, 4.028049e-13, 4.027358e-13, 4.024251e-13, 4.027836e-13, 
    4.020636e-13, 4.025258e-13, 4.017447e-13, 4.021226e-13, 4.01724e-13, 
    4.017889e-13, 4.016832e-13, 4.015955e-13, 4.014943e-13, 4.01332e-13, 
    4.013669e-13, 4.012481e-13, 4.037335e-13, 4.034836e-13, 4.03505e-13, 
    4.032592e-13, 4.030882e-13, 4.027476e-13, 4.022804e-13, 4.024453e-13, 
    4.021521e-13, 4.020981e-13, 4.025476e-13, 4.022602e-13, 4.033254e-13, 
    4.031238e-13, 4.032424e-13, 4.037131e-13, 4.024061e-13, 4.030063e-13, 
    4.01999e-13, 4.022496e-13, 4.016076e-13, 4.018934e-13, 4.013868e-13, 
    4.012326e-13, 4.011159e-13, 4.010098e-13, 4.033541e-13, 4.035161e-13, 
    4.032311e-13, 4.028736e-13, 4.025777e-13, 4.022333e-13, 4.022011e-13, 
    4.021434e-13, 4.020019e-13, 4.018914e-13, 4.021254e-13, 4.01865e-13, 
    4.030787e-13, 4.023604e-13, 4.035793e-13, 4.031575e-13, 4.028935e-13, 
    4.030066e-13, 4.02465e-13, 4.023529e-13, 4.019529e-13, 4.02149e-13, 
    4.012676e-13, 4.015778e-13, 4.009479e-13, 4.01057e-13, 4.035745e-13, 
    4.033546e-13, 4.026877e-13, 4.029868e-13, 4.022122e-13, 4.020573e-13, 
    4.019407e-13, 4.018031e-13, 4.01789e-13, 4.017142e-13, 4.018391e-13, 
    4.017189e-13, 4.022326e-13, 4.019828e-13, 4.027567e-13, 4.02542e-13, 
    4.026385e-13, 4.027488e-13, 4.024231e-13, 4.021215e-13, 4.021156e-13, 
    4.020284e-13, 4.01805e-13, 4.022096e-13, 4.012353e-13, 4.01741e-13, 
    4.031297e-13, 4.027682e-13, 4.027202e-13, 4.028526e-13, 4.020722e-13, 
    4.023242e-13, 4.01716e-13, 4.018589e-13, 4.016323e-13, 4.0174e-13, 
    4.017566e-13, 4.019111e-13, 4.020158e-13, 4.023119e-13, 4.025887e-13, 
    4.02833e-13, 4.027742e-13, 4.025127e-13, 4.021045e-13, 4.017878e-13, 
    4.018518e-13, 4.016482e-13, 4.022604e-13, 4.019745e-13, 4.020797e-13, 
    4.018187e-13, 4.024498e-13, 4.018988e-13, 4.026178e-13, 4.02544e-13, 
    4.023295e-13, 4.019567e-13, 4.018841e-13, 4.018102e-13, 4.018554e-13, 
    4.020952e-13, 4.021379e-13, 4.023345e-13, 4.023922e-13, 4.025599e-13, 
    4.02708e-13, 4.025723e-13, 4.024375e-13, 4.020951e-13, 4.018337e-13, 
    4.015943e-13, 4.015424e-13, 4.013271e-13, 4.014983e-13, 4.012332e-13, 
    4.014527e-13, 4.0111e-13, 4.018717e-13, 4.014602e-13, 4.023202e-13, 
    4.02202e-13, 4.020051e-13, 4.016295e-13, 4.018198e-13, 4.016e-13, 
    4.021396e-13, 4.025042e-13, 4.026092e-13, 4.028175e-13, 4.026046e-13, 
    4.026213e-13, 4.024321e-13, 4.024912e-13, 4.020847e-13, 4.02293e-13, 
    4.017571e-13, 4.016016e-13, 4.012596e-13, 4.011105e-13, 4.009973e-13, 
    4.009581e-13, 4.009473e-13, 4.009429e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949657e-07, 8.949656e-07, 8.949657e-07, 8.949657e-07, 
    8.949655e-07, 8.949656e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949657e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949656e-07, 
    8.949656e-07, 8.949657e-07, 8.949657e-07, 8.949657e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949654e-07, 
    8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949657e-07, 8.949657e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949653e-07, 8.949652e-07, 8.949654e-07, 8.949653e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949657e-07, 8.949657e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949656e-07, 8.949656e-07, 8.949657e-07, 8.949656e-07, 8.949657e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949653e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949655e-07, 8.949654e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949652e-07, 8.949653e-07, 8.94965e-07, 8.949651e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 
    8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949654e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949654e-07, 8.949652e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.94965e-07, 8.94965e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.760409e-16, 6.778689e-16, 6.775138e-16, 6.789867e-16, 6.7817e-16, 
    6.791341e-16, 6.764119e-16, 6.779412e-16, 6.769652e-16, 6.762059e-16, 
    6.818409e-16, 6.790525e-16, 6.847346e-16, 6.829595e-16, 6.874156e-16, 
    6.844582e-16, 6.880114e-16, 6.873309e-16, 6.893794e-16, 6.887928e-16, 
    6.914089e-16, 6.8965e-16, 6.927641e-16, 6.909893e-16, 6.912668e-16, 
    6.895919e-16, 6.796146e-16, 6.814938e-16, 6.79503e-16, 6.797712e-16, 
    6.79651e-16, 6.781867e-16, 6.77448e-16, 6.759015e-16, 6.761824e-16, 
    6.773185e-16, 6.798917e-16, 6.79019e-16, 6.812187e-16, 6.81169e-16, 
    6.836142e-16, 6.825121e-16, 6.866168e-16, 6.854514e-16, 6.888173e-16, 
    6.879714e-16, 6.887775e-16, 6.885332e-16, 6.887807e-16, 6.875399e-16, 
    6.880716e-16, 6.869796e-16, 6.827185e-16, 6.839718e-16, 6.802308e-16, 
    6.779766e-16, 6.764789e-16, 6.75415e-16, 6.755654e-16, 6.758521e-16, 
    6.773251e-16, 6.787093e-16, 6.797633e-16, 6.804679e-16, 6.811619e-16, 
    6.832594e-16, 6.843697e-16, 6.868521e-16, 6.864049e-16, 6.871628e-16, 
    6.878873e-16, 6.891021e-16, 6.889023e-16, 6.894372e-16, 6.871432e-16, 
    6.88668e-16, 6.861499e-16, 6.86839e-16, 6.813487e-16, 6.792546e-16, 
    6.783622e-16, 6.77582e-16, 6.75681e-16, 6.769939e-16, 6.764765e-16, 
    6.777077e-16, 6.784893e-16, 6.781028e-16, 6.804872e-16, 6.795605e-16, 
    6.844355e-16, 6.823374e-16, 6.878028e-16, 6.864968e-16, 6.881157e-16, 
    6.872899e-16, 6.887045e-16, 6.874315e-16, 6.896364e-16, 6.901159e-16, 
    6.897882e-16, 6.910472e-16, 6.873608e-16, 6.887773e-16, 6.780919e-16, 
    6.781549e-16, 6.784487e-16, 6.771569e-16, 6.770779e-16, 6.758937e-16, 
    6.769476e-16, 6.773961e-16, 6.785347e-16, 6.792075e-16, 6.79847e-16, 
    6.812521e-16, 6.828196e-16, 6.850096e-16, 6.865814e-16, 6.876341e-16, 
    6.869888e-16, 6.875585e-16, 6.869215e-16, 6.86623e-16, 6.899361e-16, 
    6.880765e-16, 6.908662e-16, 6.907121e-16, 6.894499e-16, 6.907294e-16, 
    6.781992e-16, 6.778365e-16, 6.765758e-16, 6.775625e-16, 6.757647e-16, 
    6.76771e-16, 6.773492e-16, 6.795795e-16, 6.800695e-16, 6.805233e-16, 
    6.814194e-16, 6.825686e-16, 6.845824e-16, 6.863329e-16, 6.879295e-16, 
    6.878126e-16, 6.878537e-16, 6.8821e-16, 6.873271e-16, 6.883549e-16, 
    6.885272e-16, 6.880765e-16, 6.906914e-16, 6.899448e-16, 6.907088e-16, 
    6.902227e-16, 6.779544e-16, 6.785648e-16, 6.78235e-16, 6.78855e-16, 
    6.784181e-16, 6.803597e-16, 6.809414e-16, 6.83661e-16, 6.825459e-16, 
    6.843208e-16, 6.827264e-16, 6.830089e-16, 6.843779e-16, 6.828127e-16, 
    6.862361e-16, 6.839153e-16, 6.882239e-16, 6.859084e-16, 6.883688e-16, 
    6.879226e-16, 6.886615e-16, 6.893228e-16, 6.901546e-16, 6.916878e-16, 
    6.91333e-16, 6.926146e-16, 6.794745e-16, 6.802653e-16, 6.80196e-16, 
    6.810234e-16, 6.81635e-16, 6.829602e-16, 6.850831e-16, 6.842853e-16, 
    6.8575e-16, 6.860439e-16, 6.838185e-16, 6.851849e-16, 6.807945e-16, 
    6.815043e-16, 6.81082e-16, 6.795367e-16, 6.844687e-16, 6.819392e-16, 
    6.866073e-16, 6.852394e-16, 6.892284e-16, 6.872455e-16, 6.911375e-16, 
    6.927975e-16, 6.943598e-16, 6.961815e-16, 6.806971e-16, 6.801599e-16, 
    6.811219e-16, 6.824513e-16, 6.836849e-16, 6.853228e-16, 6.854905e-16, 
    6.85797e-16, 6.865911e-16, 6.872584e-16, 6.858936e-16, 6.874256e-16, 
    6.816682e-16, 6.846882e-16, 6.799564e-16, 6.813823e-16, 6.823731e-16, 
    6.819389e-16, 6.841941e-16, 6.847251e-16, 6.868808e-16, 6.85767e-16, 
    6.923877e-16, 6.894619e-16, 6.975682e-16, 6.95307e-16, 6.799721e-16, 
    6.806954e-16, 6.832097e-16, 6.820139e-16, 6.854322e-16, 6.862724e-16, 
    6.869554e-16, 6.878274e-16, 6.879218e-16, 6.884383e-16, 6.875918e-16, 
    6.88405e-16, 6.853263e-16, 6.867028e-16, 6.829229e-16, 6.838435e-16, 
    6.834202e-16, 6.829555e-16, 6.843893e-16, 6.85915e-16, 6.859481e-16, 
    6.864369e-16, 6.878125e-16, 6.854461e-16, 6.927638e-16, 6.882477e-16, 
    6.814837e-16, 6.828746e-16, 6.830738e-16, 6.825351e-16, 6.861882e-16, 
    6.848654e-16, 6.884258e-16, 6.874644e-16, 6.890394e-16, 6.882569e-16, 
    6.881417e-16, 6.871362e-16, 6.865097e-16, 6.84926e-16, 6.836364e-16, 
    6.826133e-16, 6.828513e-16, 6.839749e-16, 6.860084e-16, 6.879301e-16, 
    6.875092e-16, 6.889197e-16, 6.851846e-16, 6.867516e-16, 6.86146e-16, 
    6.877248e-16, 6.842639e-16, 6.872098e-16, 6.835098e-16, 6.838347e-16, 
    6.848392e-16, 6.868575e-16, 6.873045e-16, 6.877806e-16, 6.874869e-16, 
    6.860601e-16, 6.858264e-16, 6.848149e-16, 6.845352e-16, 6.83764e-16, 
    6.83125e-16, 6.837087e-16, 6.843214e-16, 6.860609e-16, 6.876266e-16, 
    6.893321e-16, 6.897494e-16, 6.917378e-16, 6.901186e-16, 6.927889e-16, 
    6.905178e-16, 6.944476e-16, 6.873812e-16, 6.90452e-16, 6.84885e-16, 
    6.854858e-16, 6.865714e-16, 6.890596e-16, 6.877174e-16, 6.892872e-16, 
    6.858173e-16, 6.840134e-16, 6.83547e-16, 6.826754e-16, 6.83567e-16, 
    6.834945e-16, 6.843471e-16, 6.840732e-16, 6.861187e-16, 6.850203e-16, 
    6.881387e-16, 6.89275e-16, 6.924801e-16, 6.944413e-16, 6.96436e-16, 
    6.973155e-16, 6.975831e-16, 6.97695e-16 ;

 CWDC_TO_LITR2C =
  5.137911e-16, 5.151804e-16, 5.149105e-16, 5.160299e-16, 5.154092e-16, 
    5.16142e-16, 5.14073e-16, 5.152353e-16, 5.144936e-16, 5.139165e-16, 
    5.181991e-16, 5.160799e-16, 5.203983e-16, 5.190492e-16, 5.224358e-16, 
    5.201882e-16, 5.228886e-16, 5.223715e-16, 5.239283e-16, 5.234826e-16, 
    5.254707e-16, 5.24134e-16, 5.265007e-16, 5.251519e-16, 5.253628e-16, 
    5.240898e-16, 5.16507e-16, 5.179353e-16, 5.164223e-16, 5.166261e-16, 
    5.165347e-16, 5.154219e-16, 5.148605e-16, 5.136851e-16, 5.138986e-16, 
    5.14762e-16, 5.167177e-16, 5.160545e-16, 5.177262e-16, 5.176885e-16, 
    5.195468e-16, 5.187092e-16, 5.218288e-16, 5.209431e-16, 5.235011e-16, 
    5.228583e-16, 5.234709e-16, 5.232852e-16, 5.234733e-16, 5.225303e-16, 
    5.229344e-16, 5.221044e-16, 5.188661e-16, 5.198186e-16, 5.169754e-16, 
    5.152622e-16, 5.14124e-16, 5.133154e-16, 5.134297e-16, 5.136476e-16, 
    5.147671e-16, 5.158191e-16, 5.166201e-16, 5.171556e-16, 5.17683e-16, 
    5.192772e-16, 5.20121e-16, 5.220076e-16, 5.216677e-16, 5.222438e-16, 
    5.227943e-16, 5.237176e-16, 5.235657e-16, 5.239723e-16, 5.222288e-16, 
    5.233877e-16, 5.21474e-16, 5.219977e-16, 5.17825e-16, 5.162335e-16, 
    5.155552e-16, 5.149623e-16, 5.135176e-16, 5.145154e-16, 5.141221e-16, 
    5.150578e-16, 5.156518e-16, 5.153581e-16, 5.171702e-16, 5.16466e-16, 
    5.20171e-16, 5.185765e-16, 5.227301e-16, 5.217375e-16, 5.229679e-16, 
    5.223403e-16, 5.234154e-16, 5.224479e-16, 5.241237e-16, 5.244881e-16, 
    5.24239e-16, 5.251959e-16, 5.223942e-16, 5.234708e-16, 5.153498e-16, 
    5.153977e-16, 5.15621e-16, 5.146392e-16, 5.145792e-16, 5.136792e-16, 
    5.144802e-16, 5.14821e-16, 5.156864e-16, 5.161977e-16, 5.166837e-16, 
    5.177516e-16, 5.189429e-16, 5.206073e-16, 5.218019e-16, 5.226019e-16, 
    5.221115e-16, 5.225445e-16, 5.220604e-16, 5.218335e-16, 5.243515e-16, 
    5.229381e-16, 5.250583e-16, 5.249412e-16, 5.239819e-16, 5.249543e-16, 
    5.154314e-16, 5.151557e-16, 5.141977e-16, 5.149475e-16, 5.135812e-16, 
    5.14346e-16, 5.147854e-16, 5.164804e-16, 5.168528e-16, 5.171977e-16, 
    5.178787e-16, 5.187521e-16, 5.202826e-16, 5.21613e-16, 5.228264e-16, 
    5.227375e-16, 5.227688e-16, 5.230396e-16, 5.223686e-16, 5.231497e-16, 
    5.232806e-16, 5.229381e-16, 5.249254e-16, 5.24358e-16, 5.249387e-16, 
    5.245693e-16, 5.152454e-16, 5.157092e-16, 5.154586e-16, 5.159298e-16, 
    5.155977e-16, 5.170734e-16, 5.175154e-16, 5.195823e-16, 5.187348e-16, 
    5.200838e-16, 5.188721e-16, 5.190868e-16, 5.201272e-16, 5.189376e-16, 
    5.215394e-16, 5.197756e-16, 5.230501e-16, 5.212904e-16, 5.231603e-16, 
    5.228211e-16, 5.233827e-16, 5.238853e-16, 5.245175e-16, 5.256827e-16, 
    5.254131e-16, 5.263871e-16, 5.164006e-16, 5.170016e-16, 5.16949e-16, 
    5.175778e-16, 5.180426e-16, 5.190498e-16, 5.206632e-16, 5.200568e-16, 
    5.211701e-16, 5.213933e-16, 5.197021e-16, 5.207405e-16, 5.174039e-16, 
    5.179433e-16, 5.176223e-16, 5.164479e-16, 5.201962e-16, 5.182738e-16, 
    5.218215e-16, 5.207819e-16, 5.238136e-16, 5.223066e-16, 5.252646e-16, 
    5.265261e-16, 5.277134e-16, 5.290979e-16, 5.173298e-16, 5.169215e-16, 
    5.176526e-16, 5.18663e-16, 5.196005e-16, 5.208453e-16, 5.209727e-16, 
    5.212057e-16, 5.218092e-16, 5.223164e-16, 5.212791e-16, 5.224435e-16, 
    5.180678e-16, 5.20363e-16, 5.167669e-16, 5.178505e-16, 5.186036e-16, 
    5.182736e-16, 5.199875e-16, 5.20391e-16, 5.220294e-16, 5.211829e-16, 
    5.262146e-16, 5.23991e-16, 5.301518e-16, 5.284333e-16, 5.167788e-16, 
    5.173285e-16, 5.192394e-16, 5.183306e-16, 5.209285e-16, 5.21567e-16, 
    5.220861e-16, 5.227488e-16, 5.228206e-16, 5.23213e-16, 5.225698e-16, 
    5.231878e-16, 5.20848e-16, 5.218942e-16, 5.190214e-16, 5.197211e-16, 
    5.193993e-16, 5.190462e-16, 5.201359e-16, 5.212954e-16, 5.213206e-16, 
    5.21692e-16, 5.227375e-16, 5.20939e-16, 5.265005e-16, 5.230682e-16, 
    5.179276e-16, 5.189847e-16, 5.191361e-16, 5.187267e-16, 5.21503e-16, 
    5.204977e-16, 5.232036e-16, 5.22473e-16, 5.236699e-16, 5.230752e-16, 
    5.229877e-16, 5.222236e-16, 5.217474e-16, 5.205437e-16, 5.195637e-16, 
    5.187861e-16, 5.18967e-16, 5.198209e-16, 5.213664e-16, 5.228269e-16, 
    5.22507e-16, 5.23579e-16, 5.207403e-16, 5.219312e-16, 5.214709e-16, 
    5.226708e-16, 5.200406e-16, 5.222795e-16, 5.194675e-16, 5.197144e-16, 
    5.204778e-16, 5.220117e-16, 5.223514e-16, 5.227133e-16, 5.224901e-16, 
    5.214056e-16, 5.212281e-16, 5.204593e-16, 5.202467e-16, 5.196606e-16, 
    5.19175e-16, 5.196187e-16, 5.200843e-16, 5.214063e-16, 5.225962e-16, 
    5.238924e-16, 5.242095e-16, 5.257207e-16, 5.244901e-16, 5.265195e-16, 
    5.247935e-16, 5.277802e-16, 5.224097e-16, 5.247435e-16, 5.205126e-16, 
    5.209693e-16, 5.217943e-16, 5.236853e-16, 5.226652e-16, 5.238583e-16, 
    5.212211e-16, 5.198502e-16, 5.194957e-16, 5.188333e-16, 5.195109e-16, 
    5.194558e-16, 5.201038e-16, 5.198956e-16, 5.214502e-16, 5.206154e-16, 
    5.229854e-16, 5.23849e-16, 5.262849e-16, 5.277754e-16, 5.292914e-16, 
    5.299598e-16, 5.301632e-16, 5.302482e-16 ;

 CWDC_TO_LITR3C =
  1.622498e-16, 1.626885e-16, 1.626033e-16, 1.629568e-16, 1.627608e-16, 
    1.629922e-16, 1.623389e-16, 1.627059e-16, 1.624717e-16, 1.622894e-16, 
    1.636418e-16, 1.629726e-16, 1.643363e-16, 1.639103e-16, 1.649797e-16, 
    1.6427e-16, 1.651227e-16, 1.649594e-16, 1.654511e-16, 1.653103e-16, 
    1.659381e-16, 1.65516e-16, 1.662634e-16, 1.658374e-16, 1.65904e-16, 
    1.65502e-16, 1.631075e-16, 1.635585e-16, 1.630807e-16, 1.631451e-16, 
    1.631162e-16, 1.627648e-16, 1.625875e-16, 1.622164e-16, 1.622838e-16, 
    1.625564e-16, 1.63174e-16, 1.629646e-16, 1.634925e-16, 1.634806e-16, 
    1.640674e-16, 1.638029e-16, 1.64788e-16, 1.645083e-16, 1.653162e-16, 
    1.651131e-16, 1.653066e-16, 1.65248e-16, 1.653074e-16, 1.650096e-16, 
    1.651372e-16, 1.648751e-16, 1.638524e-16, 1.641532e-16, 1.632554e-16, 
    1.627144e-16, 1.623549e-16, 1.620996e-16, 1.621357e-16, 1.622045e-16, 
    1.62558e-16, 1.628902e-16, 1.631432e-16, 1.633123e-16, 1.634789e-16, 
    1.639823e-16, 1.642487e-16, 1.648445e-16, 1.647372e-16, 1.649191e-16, 
    1.650929e-16, 1.653845e-16, 1.653366e-16, 1.654649e-16, 1.649144e-16, 
    1.652803e-16, 1.64676e-16, 1.648414e-16, 1.635237e-16, 1.630211e-16, 
    1.628069e-16, 1.626197e-16, 1.621635e-16, 1.624785e-16, 1.623544e-16, 
    1.626498e-16, 1.628374e-16, 1.627447e-16, 1.633169e-16, 1.630945e-16, 
    1.642645e-16, 1.63761e-16, 1.650727e-16, 1.647592e-16, 1.651478e-16, 
    1.649496e-16, 1.652891e-16, 1.649835e-16, 1.655127e-16, 1.656278e-16, 
    1.655492e-16, 1.658513e-16, 1.649666e-16, 1.653066e-16, 1.627421e-16, 
    1.627572e-16, 1.628277e-16, 1.625176e-16, 1.624987e-16, 1.622145e-16, 
    1.624674e-16, 1.625751e-16, 1.628483e-16, 1.630098e-16, 1.631633e-16, 
    1.635005e-16, 1.638767e-16, 1.644023e-16, 1.647795e-16, 1.650322e-16, 
    1.648773e-16, 1.65014e-16, 1.648612e-16, 1.647895e-16, 1.655847e-16, 
    1.651384e-16, 1.658079e-16, 1.657709e-16, 1.65468e-16, 1.657751e-16, 
    1.627678e-16, 1.626808e-16, 1.623782e-16, 1.62615e-16, 1.621835e-16, 
    1.62425e-16, 1.625638e-16, 1.630991e-16, 1.632167e-16, 1.633256e-16, 
    1.635407e-16, 1.638164e-16, 1.642998e-16, 1.647199e-16, 1.651031e-16, 
    1.65075e-16, 1.650849e-16, 1.651704e-16, 1.649585e-16, 1.652052e-16, 
    1.652465e-16, 1.651384e-16, 1.657659e-16, 1.655867e-16, 1.657701e-16, 
    1.656535e-16, 1.627091e-16, 1.628556e-16, 1.627764e-16, 1.629252e-16, 
    1.628203e-16, 1.632863e-16, 1.634259e-16, 1.640786e-16, 1.63811e-16, 
    1.64237e-16, 1.638543e-16, 1.639221e-16, 1.642507e-16, 1.638751e-16, 
    1.646967e-16, 1.641397e-16, 1.651737e-16, 1.64618e-16, 1.652085e-16, 
    1.651014e-16, 1.652787e-16, 1.654375e-16, 1.656371e-16, 1.660051e-16, 
    1.659199e-16, 1.662275e-16, 1.630739e-16, 1.632637e-16, 1.63247e-16, 
    1.634456e-16, 1.635924e-16, 1.639105e-16, 1.644199e-16, 1.642285e-16, 
    1.6458e-16, 1.646505e-16, 1.641164e-16, 1.644444e-16, 1.633907e-16, 
    1.63561e-16, 1.634597e-16, 1.630888e-16, 1.642725e-16, 1.636654e-16, 
    1.647857e-16, 1.644575e-16, 1.654148e-16, 1.649389e-16, 1.65873e-16, 
    1.662714e-16, 1.666463e-16, 1.670835e-16, 1.633673e-16, 1.632384e-16, 
    1.634693e-16, 1.637883e-16, 1.640844e-16, 1.644775e-16, 1.645177e-16, 
    1.645913e-16, 1.647819e-16, 1.64942e-16, 1.646145e-16, 1.649822e-16, 
    1.636004e-16, 1.643252e-16, 1.631896e-16, 1.635317e-16, 1.637696e-16, 
    1.636653e-16, 1.642066e-16, 1.64334e-16, 1.648514e-16, 1.645841e-16, 
    1.66173e-16, 1.654709e-16, 1.674164e-16, 1.668737e-16, 1.631933e-16, 
    1.633669e-16, 1.639703e-16, 1.636833e-16, 1.645037e-16, 1.647054e-16, 
    1.648693e-16, 1.650786e-16, 1.651012e-16, 1.652252e-16, 1.65022e-16, 
    1.652172e-16, 1.644783e-16, 1.648087e-16, 1.639015e-16, 1.641225e-16, 
    1.640208e-16, 1.639093e-16, 1.642534e-16, 1.646196e-16, 1.646276e-16, 
    1.647449e-16, 1.65075e-16, 1.645071e-16, 1.662633e-16, 1.651794e-16, 
    1.635561e-16, 1.638899e-16, 1.639377e-16, 1.638084e-16, 1.646852e-16, 
    1.643677e-16, 1.652222e-16, 1.649915e-16, 1.653694e-16, 1.651817e-16, 
    1.65154e-16, 1.649127e-16, 1.647623e-16, 1.643822e-16, 1.640727e-16, 
    1.638272e-16, 1.638843e-16, 1.64154e-16, 1.64642e-16, 1.651032e-16, 
    1.650022e-16, 1.653407e-16, 1.644443e-16, 1.648204e-16, 1.64675e-16, 
    1.650539e-16, 1.642233e-16, 1.649304e-16, 1.640424e-16, 1.641203e-16, 
    1.643614e-16, 1.648458e-16, 1.649531e-16, 1.650673e-16, 1.649969e-16, 
    1.646544e-16, 1.645983e-16, 1.643556e-16, 1.642884e-16, 1.641034e-16, 
    1.6395e-16, 1.640901e-16, 1.642371e-16, 1.646546e-16, 1.650304e-16, 
    1.654397e-16, 1.655398e-16, 1.660171e-16, 1.656285e-16, 1.662693e-16, 
    1.657243e-16, 1.666674e-16, 1.649715e-16, 1.657085e-16, 1.643724e-16, 
    1.645166e-16, 1.647771e-16, 1.653743e-16, 1.650522e-16, 1.654289e-16, 
    1.645962e-16, 1.641632e-16, 1.640513e-16, 1.638421e-16, 1.640561e-16, 
    1.640387e-16, 1.642433e-16, 1.641776e-16, 1.646685e-16, 1.644049e-16, 
    1.651533e-16, 1.65426e-16, 1.661952e-16, 1.666659e-16, 1.671446e-16, 
    1.673557e-16, 1.6742e-16, 1.674468e-16 ;

 CWDC_vr =
  5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110347e-05, 5.110346e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110346e-05, 5.110346e-05, 5.110347e-05, 5.110346e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  1.027582e-18, 1.030361e-18, 1.029821e-18, 1.03206e-18, 1.030818e-18, 
    1.032284e-18, 1.028146e-18, 1.030471e-18, 1.028987e-18, 1.027833e-18, 
    1.036398e-18, 1.03216e-18, 1.040797e-18, 1.038099e-18, 1.044872e-18, 
    1.040376e-18, 1.045777e-18, 1.044743e-18, 1.047857e-18, 1.046965e-18, 
    1.050941e-18, 1.048268e-18, 1.053001e-18, 1.050304e-18, 1.050726e-18, 
    1.04818e-18, 1.033014e-18, 1.035871e-18, 1.032845e-18, 1.033252e-18, 
    1.033069e-18, 1.030844e-18, 1.029721e-18, 1.02737e-18, 1.027797e-18, 
    1.029524e-18, 1.033435e-18, 1.032109e-18, 1.035452e-18, 1.035377e-18, 
    1.039094e-18, 1.037418e-18, 1.043658e-18, 1.041886e-18, 1.047002e-18, 
    1.045717e-18, 1.046942e-18, 1.04657e-18, 1.046947e-18, 1.045061e-18, 
    1.045869e-18, 1.044209e-18, 1.037732e-18, 1.039637e-18, 1.033951e-18, 
    1.030524e-18, 1.028248e-18, 1.026631e-18, 1.026859e-18, 1.027295e-18, 
    1.029534e-18, 1.031638e-18, 1.03324e-18, 1.034311e-18, 1.035366e-18, 
    1.038554e-18, 1.040242e-18, 1.044015e-18, 1.043335e-18, 1.044487e-18, 
    1.045589e-18, 1.047435e-18, 1.047132e-18, 1.047945e-18, 1.044458e-18, 
    1.046775e-18, 1.042948e-18, 1.043995e-18, 1.03565e-18, 1.032467e-18, 
    1.031111e-18, 1.029925e-18, 1.027035e-18, 1.029031e-18, 1.028244e-18, 
    1.030116e-18, 1.031304e-18, 1.030716e-18, 1.03434e-18, 1.032932e-18, 
    1.040342e-18, 1.037153e-18, 1.04546e-18, 1.043475e-18, 1.045936e-18, 
    1.044681e-18, 1.046831e-18, 1.044896e-18, 1.048247e-18, 1.048976e-18, 
    1.048478e-18, 1.050392e-18, 1.044788e-18, 1.046942e-18, 1.0307e-18, 
    1.030795e-18, 1.031242e-18, 1.029278e-18, 1.029158e-18, 1.027358e-18, 
    1.02896e-18, 1.029642e-18, 1.031373e-18, 1.032395e-18, 1.033367e-18, 
    1.035503e-18, 1.037886e-18, 1.041215e-18, 1.043604e-18, 1.045204e-18, 
    1.044223e-18, 1.045089e-18, 1.044121e-18, 1.043667e-18, 1.048703e-18, 
    1.045876e-18, 1.050117e-18, 1.049882e-18, 1.047964e-18, 1.049909e-18, 
    1.030863e-18, 1.030311e-18, 1.028395e-18, 1.029895e-18, 1.027162e-18, 
    1.028692e-18, 1.029571e-18, 1.032961e-18, 1.033706e-18, 1.034395e-18, 
    1.035758e-18, 1.037504e-18, 1.040565e-18, 1.043226e-18, 1.045653e-18, 
    1.045475e-18, 1.045538e-18, 1.046079e-18, 1.044737e-18, 1.046299e-18, 
    1.046561e-18, 1.045876e-18, 1.049851e-18, 1.048716e-18, 1.049877e-18, 
    1.049139e-18, 1.030491e-18, 1.031419e-18, 1.030917e-18, 1.03186e-18, 
    1.031196e-18, 1.034147e-18, 1.035031e-18, 1.039165e-18, 1.03747e-18, 
    1.040168e-18, 1.037744e-18, 1.038174e-18, 1.040254e-18, 1.037875e-18, 
    1.043079e-18, 1.039551e-18, 1.0461e-18, 1.042581e-18, 1.046321e-18, 
    1.045642e-18, 1.046765e-18, 1.047771e-18, 1.049035e-18, 1.051365e-18, 
    1.050826e-18, 1.052774e-18, 1.032801e-18, 1.034003e-18, 1.033898e-18, 
    1.035156e-18, 1.036085e-18, 1.0381e-18, 1.041326e-18, 1.040114e-18, 
    1.04234e-18, 1.042787e-18, 1.039404e-18, 1.041481e-18, 1.034808e-18, 
    1.035887e-18, 1.035245e-18, 1.032896e-18, 1.040392e-18, 1.036548e-18, 
    1.043643e-18, 1.041564e-18, 1.047627e-18, 1.044613e-18, 1.050529e-18, 
    1.053052e-18, 1.055427e-18, 1.058196e-18, 1.03466e-18, 1.033843e-18, 
    1.035305e-18, 1.037326e-18, 1.039201e-18, 1.041691e-18, 1.041945e-18, 
    1.042411e-18, 1.043619e-18, 1.044633e-18, 1.042558e-18, 1.044887e-18, 
    1.036136e-18, 1.040726e-18, 1.033534e-18, 1.035701e-18, 1.037207e-18, 
    1.036547e-18, 1.039975e-18, 1.040782e-18, 1.044059e-18, 1.042366e-18, 
    1.052429e-18, 1.047982e-18, 1.060304e-18, 1.056867e-18, 1.033558e-18, 
    1.034657e-18, 1.038479e-18, 1.036661e-18, 1.041857e-18, 1.043134e-18, 
    1.044172e-18, 1.045498e-18, 1.045641e-18, 1.046426e-18, 1.045139e-18, 
    1.046376e-18, 1.041696e-18, 1.043788e-18, 1.038043e-18, 1.039442e-18, 
    1.038799e-18, 1.038092e-18, 1.040272e-18, 1.042591e-18, 1.042641e-18, 
    1.043384e-18, 1.045475e-18, 1.041878e-18, 1.053001e-18, 1.046136e-18, 
    1.035855e-18, 1.037969e-18, 1.038272e-18, 1.037453e-18, 1.043006e-18, 
    1.040995e-18, 1.046407e-18, 1.044946e-18, 1.04734e-18, 1.046151e-18, 
    1.045975e-18, 1.044447e-18, 1.043495e-18, 1.041087e-18, 1.039127e-18, 
    1.037572e-18, 1.037934e-18, 1.039642e-18, 1.042733e-18, 1.045654e-18, 
    1.045014e-18, 1.047158e-18, 1.041481e-18, 1.043862e-18, 1.042942e-18, 
    1.045342e-18, 1.040081e-18, 1.044559e-18, 1.038935e-18, 1.039429e-18, 
    1.040956e-18, 1.044023e-18, 1.044703e-18, 1.045427e-18, 1.04498e-18, 
    1.042811e-18, 1.042456e-18, 1.040919e-18, 1.040494e-18, 1.039321e-18, 
    1.03835e-18, 1.039237e-18, 1.040168e-18, 1.042813e-18, 1.045192e-18, 
    1.047785e-18, 1.048419e-18, 1.051441e-18, 1.04898e-18, 1.053039e-18, 
    1.049587e-18, 1.05556e-18, 1.044819e-18, 1.049487e-18, 1.041025e-18, 
    1.041939e-18, 1.043589e-18, 1.047371e-18, 1.04533e-18, 1.047717e-18, 
    1.042442e-18, 1.0397e-18, 1.038991e-18, 1.037667e-18, 1.039022e-18, 
    1.038912e-18, 1.040208e-18, 1.039791e-18, 1.0429e-18, 1.041231e-18, 
    1.045971e-18, 1.047698e-18, 1.05257e-18, 1.055551e-18, 1.058583e-18, 
    1.05992e-18, 1.060326e-18, 1.060496e-18 ;

 CWDN_TO_LITR3N =
  3.244996e-19, 3.253771e-19, 3.252066e-19, 3.259136e-19, 3.255216e-19, 
    3.259844e-19, 3.246777e-19, 3.254118e-19, 3.249433e-19, 3.245788e-19, 
    3.272836e-19, 3.259452e-19, 3.286726e-19, 3.278206e-19, 3.299595e-19, 
    3.285399e-19, 3.302454e-19, 3.299188e-19, 3.309021e-19, 3.306205e-19, 
    3.318762e-19, 3.31032e-19, 3.325267e-19, 3.316748e-19, 3.318081e-19, 
    3.310041e-19, 3.26215e-19, 3.27117e-19, 3.261615e-19, 3.262902e-19, 
    3.262325e-19, 3.255296e-19, 3.25175e-19, 3.244327e-19, 3.245676e-19, 
    3.251129e-19, 3.26348e-19, 3.259291e-19, 3.26985e-19, 3.269611e-19, 
    3.281348e-19, 3.276058e-19, 3.295761e-19, 3.290167e-19, 3.306323e-19, 
    3.302263e-19, 3.306132e-19, 3.304959e-19, 3.306147e-19, 3.300192e-19, 
    3.302744e-19, 3.297502e-19, 3.277049e-19, 3.283065e-19, 3.265108e-19, 
    3.254288e-19, 3.247099e-19, 3.241992e-19, 3.242714e-19, 3.24409e-19, 
    3.251161e-19, 3.257805e-19, 3.262864e-19, 3.266246e-19, 3.269577e-19, 
    3.279645e-19, 3.284975e-19, 3.29689e-19, 3.294743e-19, 3.298382e-19, 
    3.301859e-19, 3.30769e-19, 3.306731e-19, 3.309299e-19, 3.298287e-19, 
    3.305606e-19, 3.29352e-19, 3.296827e-19, 3.270474e-19, 3.260422e-19, 
    3.256138e-19, 3.252394e-19, 3.243269e-19, 3.249571e-19, 3.247087e-19, 
    3.252997e-19, 3.256749e-19, 3.254894e-19, 3.266338e-19, 3.261891e-19, 
    3.28529e-19, 3.27522e-19, 3.301453e-19, 3.295184e-19, 3.302955e-19, 
    3.298991e-19, 3.305782e-19, 3.299671e-19, 3.310255e-19, 3.312556e-19, 
    3.310983e-19, 3.317027e-19, 3.299332e-19, 3.306131e-19, 3.254841e-19, 
    3.255144e-19, 3.256554e-19, 3.250353e-19, 3.249974e-19, 3.24429e-19, 
    3.249348e-19, 3.251501e-19, 3.256967e-19, 3.260196e-19, 3.263266e-19, 
    3.27001e-19, 3.277534e-19, 3.288046e-19, 3.295591e-19, 3.300643e-19, 
    3.297546e-19, 3.300281e-19, 3.297223e-19, 3.295791e-19, 3.311693e-19, 
    3.302767e-19, 3.316158e-19, 3.315418e-19, 3.309359e-19, 3.315501e-19, 
    3.255356e-19, 3.253615e-19, 3.247564e-19, 3.2523e-19, 3.243671e-19, 
    3.248501e-19, 3.251276e-19, 3.261982e-19, 3.264334e-19, 3.266512e-19, 
    3.270813e-19, 3.276329e-19, 3.285996e-19, 3.294398e-19, 3.302062e-19, 
    3.3015e-19, 3.301698e-19, 3.303408e-19, 3.29917e-19, 3.304104e-19, 
    3.30493e-19, 3.302767e-19, 3.315319e-19, 3.311735e-19, 3.315402e-19, 
    3.313069e-19, 3.254181e-19, 3.257111e-19, 3.255528e-19, 3.258504e-19, 
    3.256407e-19, 3.265726e-19, 3.268519e-19, 3.281573e-19, 3.27622e-19, 
    3.28474e-19, 3.277087e-19, 3.278443e-19, 3.285014e-19, 3.277501e-19, 
    3.293933e-19, 3.282793e-19, 3.303475e-19, 3.29236e-19, 3.30417e-19, 
    3.302028e-19, 3.305575e-19, 3.308749e-19, 3.312742e-19, 3.320102e-19, 
    3.318398e-19, 3.32455e-19, 3.261478e-19, 3.265273e-19, 3.264941e-19, 
    3.268912e-19, 3.271848e-19, 3.278209e-19, 3.288399e-19, 3.284569e-19, 
    3.2916e-19, 3.29301e-19, 3.282329e-19, 3.288887e-19, 3.267814e-19, 
    3.271221e-19, 3.269194e-19, 3.261776e-19, 3.28545e-19, 3.273308e-19, 
    3.295715e-19, 3.289149e-19, 3.308296e-19, 3.298778e-19, 3.31746e-19, 
    3.325428e-19, 3.332927e-19, 3.341671e-19, 3.267346e-19, 3.264767e-19, 
    3.269385e-19, 3.275766e-19, 3.281687e-19, 3.289549e-19, 3.290354e-19, 
    3.291825e-19, 3.295637e-19, 3.29884e-19, 3.292289e-19, 3.299643e-19, 
    3.272007e-19, 3.286503e-19, 3.263791e-19, 3.270635e-19, 3.275391e-19, 
    3.273307e-19, 3.284132e-19, 3.28668e-19, 3.297028e-19, 3.291681e-19, 
    3.323461e-19, 3.309417e-19, 3.348327e-19, 3.337474e-19, 3.263866e-19, 
    3.267338e-19, 3.279407e-19, 3.273667e-19, 3.290075e-19, 3.294107e-19, 
    3.297386e-19, 3.301571e-19, 3.302025e-19, 3.304504e-19, 3.300441e-19, 
    3.304344e-19, 3.289566e-19, 3.296174e-19, 3.27803e-19, 3.282449e-19, 
    3.280417e-19, 3.278186e-19, 3.285069e-19, 3.292392e-19, 3.292551e-19, 
    3.294897e-19, 3.3015e-19, 3.290141e-19, 3.325267e-19, 3.303589e-19, 
    3.271122e-19, 3.277798e-19, 3.278754e-19, 3.276168e-19, 3.293703e-19, 
    3.287354e-19, 3.304444e-19, 3.299829e-19, 3.307389e-19, 3.303633e-19, 
    3.30308e-19, 3.298254e-19, 3.295247e-19, 3.287645e-19, 3.281455e-19, 
    3.276544e-19, 3.277686e-19, 3.28308e-19, 3.29284e-19, 3.302064e-19, 
    3.300044e-19, 3.306815e-19, 3.288886e-19, 3.296408e-19, 3.293501e-19, 
    3.301079e-19, 3.284467e-19, 3.298607e-19, 3.280847e-19, 3.282407e-19, 
    3.287228e-19, 3.296916e-19, 3.299061e-19, 3.301347e-19, 3.299937e-19, 
    3.293088e-19, 3.291967e-19, 3.287111e-19, 3.285769e-19, 3.282067e-19, 
    3.279e-19, 3.281802e-19, 3.284743e-19, 3.293092e-19, 3.300608e-19, 
    3.308794e-19, 3.310797e-19, 3.320341e-19, 3.312569e-19, 3.325387e-19, 
    3.314485e-19, 3.333349e-19, 3.29943e-19, 3.31417e-19, 3.287448e-19, 
    3.290332e-19, 3.295543e-19, 3.307486e-19, 3.301043e-19, 3.308579e-19, 
    3.291923e-19, 3.283264e-19, 3.281026e-19, 3.276842e-19, 3.281122e-19, 
    3.280774e-19, 3.284866e-19, 3.283551e-19, 3.293369e-19, 3.288097e-19, 
    3.303066e-19, 3.30852e-19, 3.323905e-19, 3.333319e-19, 3.342893e-19, 
    3.347114e-19, 3.348399e-19, 3.348936e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.904545e-44, 0, 3.640714e-41, 
    2.382207e-44, 1.485699e-40, 2.970192e-41, 3.462017e-39, 9.090784e-40, 
    3.043702e-37, 6.372947e-39, 5.297037e-36, 1.228662e-37, 2.240759e-37, 
    5.592868e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 
    5.327737e-42, 3.012792e-43, 9.616453e-40, 1.350768e-40, 8.778827e-40, 
    4.997395e-40, 8.843286e-40, 4.883105e-41, 1.708729e-40, 1.279946e-41, 0, 
    7.006492e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    1.961818e-44, 9.427936e-42, 3.179546e-42, 1.989283e-41, 1.108483e-40, 
    1.845646e-39, 1.168838e-39, 3.948533e-39, 1.895536e-41, 6.828597e-40, 
    1.702578e-42, 9.121052e-42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.242078e-44, 0, 9.087421e-41, 3.976885e-42, 1.893603e-40, 2.691614e-41, 
    7.425691e-40, 3.771455e-41, 6.183549e-39, 1.806158e-38, 8.695494e-39, 
    1.391768e-37, 3.187954e-41, 8.78027e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9.949219e-44, 4.887729e-42, 6.099011e-41, 1.308112e-41, 
    5.099465e-41, 1.112771e-41, 5.404808e-42, 1.210799e-38, 1.728852e-40, 
    9.393621e-38, 6.709526e-38, 4.063952e-39, 6.969254e-38, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3.363116e-44, 2.668072e-42, 1.22367e-40, 9.295093e-41, 
    1.024097e-40, 2.360095e-40, 2.942166e-41, 3.306658e-40, 4.932346e-40, 
    1.727591e-40, 6.41323e-38, 1.233066e-38, 6.661603e-38, 2.286338e-38, 0, 
    0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 1.681558e-44, 0, 0, 1.961818e-44, 0, 
    2.107553e-42, 5.605194e-45, 2.437545e-40, 9.416726e-43, 3.41488e-40, 
    1.20401e-40, 6.718792e-40, 3.047178e-39, 1.966447e-38, 5.518767e-37, 
    2.580681e-37, 3.881303e-36, 0, 0, 0, 0, 0, 0, 1.191104e-43, 1.541428e-44, 
    6.347882e-43, 1.311615e-42, 4.203895e-45, 1.541428e-43, 0, 0, 0, 0, 
    2.522337e-44, 0, 5.205824e-42, 1.765636e-43, 2.460338e-39, 2.425227e-41, 
    1.693173e-37, 5.68547e-36, 1.346246e-34, 4.604947e-33, 0, 0, 0, 0, 
    2.802597e-45, 2.186026e-43, 3.321077e-43, 7.132609e-43, 5.002636e-42, 
    2.496693e-41, 9.066401e-43, 3.719607e-41, 0, 4.344025e-44, 0, 0, 0, 0, 
    1.261169e-44, 4.764415e-44, 1.009916e-41, 6.614129e-43, 2.424143e-36, 
    4.18154e-39, 6.026268e-32, 8.63849e-34, 0, 0, 1.401298e-45, 0, 
    2.872662e-43, 2.299531e-42, 1.206938e-41, 9.634768e-41, 1.20202e-40, 
    4.013333e-40, 5.518173e-41, 3.713385e-40, 2.200039e-43, 6.562281e-42, 0, 
    5.605194e-45, 1.401298e-45, 0, 2.101948e-44, 9.556856e-43, 1.03556e-42, 
    3.440188e-42, 9.359973e-41, 2.970753e-43, 5.321813e-36, 2.591547e-40, 0, 
    0, 0, 0, 1.870733e-42, 6.866362e-44, 3.897558e-40, 4.0789e-41, 
    1.598796e-39, 2.632255e-40, 2.012363e-40, 1.863867e-41, 4.105805e-42, 
    7.987401e-44, 2.802597e-45, 0, 0, 7.006492e-45, 1.203715e-42, 
    1.226613e-40, 4.54329e-41, 1.216202e-39, 1.541428e-43, 7.390448e-42, 
    1.688565e-42, 7.559725e-41, 1.541428e-44, 2.236612e-41, 1.401298e-45, 
    4.203895e-45, 6.445973e-44, 9.556856e-42, 2.787043e-41, 8.629336e-41, 
    4.303107e-41, 1.366266e-42, 7.665103e-43, 6.025583e-44, 2.942727e-44, 
    4.203895e-45, 1.401298e-45, 4.203895e-45, 1.681558e-44, 1.367667e-42, 
    5.998398e-41, 3.113122e-39, 7.966207e-39, 6.155813e-37, 1.82089e-38, 
    5.606511e-36, 4.415561e-38, 1.609795e-34, 3.358352e-41, 3.807932e-38, 
    7.286752e-44, 3.279038e-43, 4.778428e-42, 1.678356e-39, 7.428563e-41, 
    2.815552e-39, 7.496947e-43, 8.407791e-45, 2.802597e-45, 0, 2.802597e-45, 
    1.401298e-45, 1.821688e-44, 8.407791e-45, 1.576461e-42, 1.022948e-43, 
    1.99912e-40, 2.737107e-39, 2.934797e-36, 1.585659e-34, 7.423095e-33, 
    3.795473e-32, 6.187504e-32, 7.582037e-32 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  23.77457, 23.83677, 23.82469, 23.87484, 23.84705, 23.87987, 23.78721, 
    23.8392, 23.80603, 23.78022, 23.97214, 23.87709, 24.07142, 24.01063, 
    24.16357, 24.0619, 24.1841, 24.16073, 24.23133, 24.21111, 24.30128, 
    24.24067, 24.34822, 24.28685, 24.29641, 24.23866, 23.8963, 23.96027, 
    23.89249, 23.90161, 23.89754, 23.84759, 23.82237, 23.76989, 23.77943, 
    23.81802, 23.90572, 23.876, 23.95111, 23.94942, 24.03307, 23.99534, 
    24.13616, 24.09613, 24.21195, 24.18279, 24.21056, 24.20215, 24.21067, 
    24.16792, 24.18623, 24.14865, 24.00238, 24.04531, 23.91731, 23.84033, 
    23.78948, 23.75335, 23.75846, 23.76817, 23.81824, 23.86544, 23.9014, 
    23.92545, 23.94917, 24.02077, 24.0589, 24.14421, 24.12889, 24.15491, 
    24.1799, 24.22175, 24.21487, 24.2333, 24.15428, 24.20676, 24.12015, 
    24.14381, 23.95529, 23.88403, 23.85348, 23.827, 23.76238, 23.80698, 
    23.78938, 23.83132, 23.85793, 23.84478, 23.92611, 23.89447, 24.06116, 
    23.98932, 24.17698, 24.13204, 24.18777, 24.15934, 24.20803, 24.16421, 
    24.24018, 24.2567, 24.2454, 24.28891, 24.16177, 24.21053, 23.8444, 
    23.84654, 23.85656, 23.81252, 23.80984, 23.76961, 23.80544, 23.82067, 
    23.8595, 23.88242, 23.90423, 23.95223, 24.00581, 24.0809, 24.13495, 
    24.17119, 24.14899, 24.16858, 24.14667, 24.13641, 24.25049, 24.18638, 
    24.28265, 24.27733, 24.23372, 24.27793, 23.84805, 23.83571, 23.79278, 
    23.82638, 23.76523, 23.79941, 23.81904, 23.89506, 23.91185, 23.92732, 
    23.95796, 23.99727, 24.06625, 24.12638, 24.18136, 24.17734, 24.17875, 
    24.19101, 24.16061, 24.196, 24.20191, 24.18641, 24.27661, 24.25084, 
    24.27721, 24.26044, 23.83973, 23.86051, 23.84928, 23.87039, 23.85549, 
    23.92167, 23.94153, 24.03461, 23.99647, 24.05726, 24.00267, 24.01232, 
    24.05911, 24.00564, 24.123, 24.04329, 24.19148, 24.11168, 24.19648, 
    24.18112, 24.20658, 24.22935, 24.25808, 24.311, 24.29875, 24.34309, 
    23.89154, 23.91848, 23.91617, 23.94443, 23.96531, 24.01069, 24.08346, 
    24.0561, 24.10639, 24.11647, 24.04011, 24.08693, 23.93657, 23.96078, 
    23.94641, 23.89363, 24.06232, 23.97566, 24.13583, 24.08883, 24.2261, 
    24.15774, 24.292, 24.34931, 24.40357, 24.4667, 23.93326, 23.91494, 
    23.9478, 23.99319, 24.0355, 24.09169, 24.09747, 24.10799, 24.13531, 
    24.15825, 24.11125, 24.16401, 23.96627, 24.06988, 23.90796, 23.95659, 
    23.99054, 23.97571, 24.05299, 24.0712, 24.14521, 24.10698, 24.3351, 
    24.23408, 24.515, 24.43635, 23.90852, 23.93323, 24.01918, 23.97828, 
    24.09547, 24.12432, 24.14784, 24.17781, 24.18109, 24.19886, 24.16973, 
    24.19773, 24.09181, 24.13913, 24.00943, 24.04094, 24.02646, 24.01054, 
    24.05968, 24.11198, 24.1132, 24.12995, 24.17702, 24.09595, 24.34797, 
    24.19205, 23.96017, 24.00766, 24.01457, 23.99614, 24.12143, 24.07599, 
    24.19844, 24.16535, 24.2196, 24.19263, 24.18866, 24.15405, 24.13249, 
    24.07806, 24.03383, 23.99883, 24.00697, 24.04543, 24.1152, 24.18134, 
    24.16683, 24.21548, 24.08697, 24.14077, 24.11994, 24.1743, 24.05536, 
    24.15633, 24.02953, 24.04066, 24.07509, 24.14436, 24.15984, 24.1762, 
    24.16612, 24.11699, 24.10899, 24.07428, 24.06465, 24.03825, 24.01635, 
    24.03633, 24.0573, 24.11705, 24.17089, 24.22966, 24.24409, 24.31259, 
    24.25669, 24.34882, 24.27028, 24.40639, 24.16233, 24.26817, 24.07669, 
    24.09732, 24.13454, 24.22019, 24.17404, 24.22806, 24.10868, 24.04671, 
    24.0308, 24.00094, 24.03148, 24.029, 24.05824, 24.04885, 24.11904, 
    24.08133, 24.18853, 24.22766, 24.33841, 24.40631, 24.47566, 24.50624, 
    24.51556, 24.51945 ;

 EFLX_LH_TOT_R =
  23.77457, 23.83677, 23.82469, 23.87484, 23.84705, 23.87987, 23.78721, 
    23.8392, 23.80603, 23.78022, 23.97214, 23.87709, 24.07142, 24.01063, 
    24.16357, 24.0619, 24.1841, 24.16073, 24.23133, 24.21111, 24.30128, 
    24.24067, 24.34822, 24.28685, 24.29641, 24.23866, 23.8963, 23.96027, 
    23.89249, 23.90161, 23.89754, 23.84759, 23.82237, 23.76989, 23.77943, 
    23.81802, 23.90572, 23.876, 23.95111, 23.94942, 24.03307, 23.99534, 
    24.13616, 24.09613, 24.21195, 24.18279, 24.21056, 24.20215, 24.21067, 
    24.16792, 24.18623, 24.14865, 24.00238, 24.04531, 23.91731, 23.84033, 
    23.78948, 23.75335, 23.75846, 23.76817, 23.81824, 23.86544, 23.9014, 
    23.92545, 23.94917, 24.02077, 24.0589, 24.14421, 24.12889, 24.15491, 
    24.1799, 24.22175, 24.21487, 24.2333, 24.15428, 24.20676, 24.12015, 
    24.14381, 23.95529, 23.88403, 23.85348, 23.827, 23.76238, 23.80698, 
    23.78938, 23.83132, 23.85793, 23.84478, 23.92611, 23.89447, 24.06116, 
    23.98932, 24.17698, 24.13204, 24.18777, 24.15934, 24.20803, 24.16421, 
    24.24018, 24.2567, 24.2454, 24.28891, 24.16177, 24.21053, 23.8444, 
    23.84654, 23.85656, 23.81252, 23.80984, 23.76961, 23.80544, 23.82067, 
    23.8595, 23.88242, 23.90423, 23.95223, 24.00581, 24.0809, 24.13495, 
    24.17119, 24.14899, 24.16858, 24.14667, 24.13641, 24.25049, 24.18638, 
    24.28265, 24.27733, 24.23372, 24.27793, 23.84805, 23.83571, 23.79278, 
    23.82638, 23.76523, 23.79941, 23.81904, 23.89506, 23.91185, 23.92732, 
    23.95796, 23.99727, 24.06625, 24.12638, 24.18136, 24.17734, 24.17875, 
    24.19101, 24.16061, 24.196, 24.20191, 24.18641, 24.27661, 24.25084, 
    24.27721, 24.26044, 23.83973, 23.86051, 23.84928, 23.87039, 23.85549, 
    23.92167, 23.94153, 24.03461, 23.99647, 24.05726, 24.00267, 24.01232, 
    24.05911, 24.00564, 24.123, 24.04329, 24.19148, 24.11168, 24.19648, 
    24.18112, 24.20658, 24.22935, 24.25808, 24.311, 24.29875, 24.34309, 
    23.89154, 23.91848, 23.91617, 23.94443, 23.96531, 24.01069, 24.08346, 
    24.0561, 24.10639, 24.11647, 24.04011, 24.08693, 23.93657, 23.96078, 
    23.94641, 23.89363, 24.06232, 23.97566, 24.13583, 24.08883, 24.2261, 
    24.15774, 24.292, 24.34931, 24.40357, 24.4667, 23.93326, 23.91494, 
    23.9478, 23.99319, 24.0355, 24.09169, 24.09747, 24.10799, 24.13531, 
    24.15825, 24.11125, 24.16401, 23.96627, 24.06988, 23.90796, 23.95659, 
    23.99054, 23.97571, 24.05299, 24.0712, 24.14521, 24.10698, 24.3351, 
    24.23408, 24.515, 24.43635, 23.90852, 23.93323, 24.01918, 23.97828, 
    24.09547, 24.12432, 24.14784, 24.17781, 24.18109, 24.19886, 24.16973, 
    24.19773, 24.09181, 24.13913, 24.00943, 24.04094, 24.02646, 24.01054, 
    24.05968, 24.11198, 24.1132, 24.12995, 24.17702, 24.09595, 24.34797, 
    24.19205, 23.96017, 24.00766, 24.01457, 23.99614, 24.12143, 24.07599, 
    24.19844, 24.16535, 24.2196, 24.19263, 24.18866, 24.15405, 24.13249, 
    24.07806, 24.03383, 23.99883, 24.00697, 24.04543, 24.1152, 24.18134, 
    24.16683, 24.21548, 24.08697, 24.14077, 24.11994, 24.1743, 24.05536, 
    24.15633, 24.02953, 24.04066, 24.07509, 24.14436, 24.15984, 24.1762, 
    24.16612, 24.11699, 24.10899, 24.07428, 24.06465, 24.03825, 24.01635, 
    24.03633, 24.0573, 24.11705, 24.17089, 24.22966, 24.24409, 24.31259, 
    24.25669, 24.34882, 24.27028, 24.40639, 24.16233, 24.26817, 24.07669, 
    24.09732, 24.13454, 24.22019, 24.17404, 24.22806, 24.10868, 24.04671, 
    24.0308, 24.00094, 24.03148, 24.029, 24.05824, 24.04885, 24.11904, 
    24.08133, 24.18853, 24.22766, 24.33841, 24.40631, 24.47566, 24.50624, 
    24.51556, 24.51945 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 ERRH2O =
  -22918.68, -22953.21, -22946.44, -22974.69, -22958.97, -22977.54, 
    -22925.62, -22954.6, -22936.04, -22921.76, -23030.73, -22975.96, 
    -23089.37, -23053.11, -23144.9, -23083.67, -23157.47, -23143.1, 
    -23186.74, -23174.12, -23231.19, -23192.59, -23261.58, -23221.88, 
    -23228.03, -23191.33, -22986.87, -23023.84, -22984.7, -22989.93, 
    -22987.58, -22959.29, -22945.21, -22916.05, -22921.32, -22942.74, 
    -22992.28, -22975.31, -23018.36, -23017.38, -23066.38, -23044.11, 
    -23128.17, -23104.11, -23174.64, -23156.61, -23173.79, -23168.56, 
    -23173.86, -23147.5, -23158.74, -23135.74, -23048.25, -23073.68, 
    -22998.92, -22955.29, -22926.88, -22906.97, -22909.78, -22915.14, 
    -22942.86, -22969.33, -22989.76, -23003.57, -23017.24, -23059.2, 
    -23081.85, -23133.08, -23123.77, -23139.58, -23154.83, -23180.77, 
    -23176.47, -23188, -23139.16, -23171.46, -23118.48, -23132.8, -23020.97, 
    -22979.87, -22962.67, -22947.74, -22911.94, -22936.59, -22926.84, 
    -22950.13, -22965.09, -22957.68, -23003.95, -22985.81, -23083.2, 
    -23040.61, -23153.04, -23125.68, -23159.67, -23142.23, -23172.23, 
    -23145.21, -23192.3, -23202.73, -23195.6, -23223.15, -23143.72, 
    -23173.79, -22957.47, -22958.68, -22964.31, -22939.68, -22938.18, 
    -22915.91, -22935.71, -22944.21, -22965.96, -22978.96, -22991.4, 
    -23019.02, -23050.3, -23095.05, -23127.44, -23149.48, -23135.92, 
    -23147.88, -23134.52, -23128.29, -23198.82, -23158.85, -23219.16, 
    -23215.77, -23188.27, -23216.15, -22959.53, -22952.58, -22928.71, 
    -22947.36, -22913.5, -22932.38, -22943.32, -22986.19, -22995.75, 
    -23004.67, -23022.33, -23045.24, -23086.21, -23122.28, -23155.72, 
    -23153.25, -23154.12, -23161.68, -23143.02, -23164.76, -23168.44, 
    -23158.84, -23215.31, -23198.99, -23215.7, -23205.05, -22954.84, 
    -22966.54, -22960.21, -22972.14, -22963.73, -23001.46, -23012.91, 
    -23067.35, -23044.79, -23080.83, -23048.41, -23054.11, -23082.03, 
    -23050.14, -23120.29, -23072.54, -23161.97, -23113.53, -23165.06, 
    -23155.58, -23171.3, -23185.52, -23203.56, -23237.38, -23229.49, 
    -23258.19, -22984.14, -22999.6, -22998.23, -23014.51, -23026.6, 
    -23053.12, -23096.57, -23080.09, -23110.24, -23116.3, -23070.54, 
    -23098.68, -23010.01, -23024.02, -23015.67, -22985.35, -23083.88, 
    -23032.66, -23127.98, -23099.78, -23183.49, -23141.32, -23225.16, 
    -23262.36, -23298.18, -23340.73, -23008.09, -22997.52, -23016.45, 
    -23042.9, -23067.82, -23101.49, -23104.91, -23111.21, -23127.63, 
    -23141.57, -23113.21, -23145.09, -23027.29, -23088.4, -22993.54, 
    -23021.61, -23041.33, -23032.64, -23078.22, -23089.15, -23133.68, 
    -23110.59, -23253.1, -23188.54, -23373.44, -23320.33, -22993.84, 
    -23008.05, -23058.17, -23034.14, -23103.72, -23121.02, -23135.23, 
    -23153.57, -23155.56, -23166.54, -23148.59, -23165.83, -23101.56, 
    -23129.96, -23052.37, -23071.05, -23062.43, -23053.02, -23082.23, 
    -23113.65, -23114.32, -23124.44, -23153.31, -23104.01, -23261.63, 
    -23162.53, -23023.6, -23051.41, -23055.42, -23044.56, -23119.28, 
    -23092.05, -23166.27, -23145.9, -23179.41, -23162.67, -23160.23, 
    -23139.01, -23125.95, -23093.31, -23066.83, -23046.13, -23050.92, 
    -23073.74, -23115.58, -23155.74, -23146.86, -23176.84, -23098.66, 
    -23130.98, -23118.42, -23151.39, -23079.66, -23140.61, -23064.25, 
    -23070.87, -23091.51, -23133.2, -23142.54, -23152.58, -23146.38, 
    -23116.64, -23111.82, -23091, -23085.24, -23069.42, -23056.45, -23068.3, 
    -23080.84, -23116.65, -23149.33, -23185.73, -23194.75, -23238.53, 
    -23202.81, -23262.2, -23211.57, -23300.28, -23144.18, -23210.1, 
    -23092.46, -23104.82, -23127.24, -23179.87, -23151.24, -23184.77, 
    -23111.63, -23074.54, -23065.01, -23047.38, -23065.41, -23063.94, 
    -23081.36, -23075.74, -23117.84, -23095.26, -23160.17, -23184.5, 
    -23255.16, -23300.1, -23346.67, -23367.43, -23373.78, -23376.45 ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -1.350608e-14, -1.156243e-14, -6.650601e-15, -1.670047e-14, -1.83785e-14, 
    -2.504105e-14, -1.61773e-14, -4.35947e-15, -1.735697e-14, -1.197693e-14, 
    -1.615249e-14, -4.201965e-15, -1.487777e-14, -2.383231e-14, 
    -1.307129e-14, -1.594587e-14, -1.172673e-14, -1.635951e-14, 
    -5.258168e-15, -9.227459e-15, -1.169335e-14, -1.219595e-14, 
    -1.637282e-14, -1.755731e-14, -8.189196e-15, -9.399165e-15, 
    -6.631955e-15, -7.550463e-15, -1.12933e-14, -2.546021e-14, -1.39384e-14, 
    -1.467608e-14, -6.567065e-15, -1.184686e-14, -1.643275e-14, 
    -1.637466e-14, -8.118534e-15, -1.443269e-14, -8.316461e-15, 
    -1.371641e-14, -1.962525e-15, -2.00728e-14, -2.344144e-14, -2.21421e-14, 
    -1.610667e-14, -1.504466e-14, -1.305255e-14, -1.160459e-14, 
    -1.478157e-14, -1.70523e-14, -1.448308e-14, -1.727593e-14, -4.033055e-15, 
    -1.235181e-14, -1.993116e-14, -1.400814e-14, -8.329989e-15, 
    -1.270911e-14, -9.016129e-15, -1.167585e-14, -2.410661e-14, 
    -1.204484e-14, -1.447033e-14, -1.488882e-14, -2.25621e-14, -1.40694e-14, 
    -6.332509e-15, -1.215066e-14, -1.966954e-14, -7.183703e-15, 
    -1.506224e-14, -5.313774e-15, -1.765622e-14, -7.895271e-15, 
    -1.372735e-14, -1.433026e-14, -1.226677e-14, -2.007271e-14, 
    -2.162009e-14, -1.642662e-14, -5.49624e-15, -1.299438e-14, -1.749103e-14, 
    -1.121292e-14, -1.376483e-14, -1.561913e-14, -1.274483e-14, -1.09565e-14, 
    -1.162882e-14, -6.817703e-15, -1.263829e-14, -4.487106e-15, 
    -1.836996e-14, -1.362619e-14, -1.446422e-14, -6.755466e-15, 
    -1.022536e-14, -2.335367e-14, -9.853401e-15, -1.76207e-14, -1.610233e-14, 
    -6.95854e-15, -1.23714e-14, -2.268839e-14, -1.292773e-14, -1.814044e-14, 
    -1.68639e-14, -1.601625e-14, -1.852653e-14, -1.088853e-14, -1.576847e-14, 
    -1.134139e-14, -2.087519e-14, -1.871688e-14, -3.474242e-15, 
    -1.438201e-14, -1.104671e-14, -2.609646e-14, -1.19462e-14, -1.569307e-14, 
    -1.033372e-14, -1.161857e-14, -1.357566e-14, -1.186285e-14, 
    -1.706687e-14, -1.354355e-14, -1.535045e-14, -1.270974e-14, 
    -6.262219e-15, -1.21562e-14, -1.592315e-14, -1.429938e-14, -1.051323e-14, 
    -1.023053e-14, -1.959165e-14, -5.772926e-15, -2.577438e-14, 
    -1.616016e-14, -1.661222e-14, -9.835942e-15, -1.566263e-14, 
    -7.526681e-15, -1.682889e-14, -2.367842e-14, -7.043925e-15, 
    -1.262215e-14, -1.993505e-14, -1.163688e-14, -1.806022e-14, 
    -1.268745e-14, -1.928179e-14, -2.012736e-14, -1.964656e-14, 
    -5.080493e-15, -5.467643e-15, -1.672225e-14, -1.339783e-14, 
    -1.172458e-14, -9.679425e-15, -1.306686e-14, -1.448128e-14, 
    -1.549237e-14, -1.365668e-14, -7.368283e-15, -8.938197e-15, 
    -8.354683e-15, -1.464643e-14, -1.199508e-14, -1.702493e-14, 
    -1.423939e-14, -1.849828e-14, -1.585521e-14, -4.634186e-15, -9.91457e-15, 
    -1.414342e-14, -1.608452e-14, -1.509293e-14, -1.924072e-14, 
    -2.026222e-14, -1.161819e-14, -1.527722e-14, -1.607438e-14, 
    -1.021613e-14, -1.246885e-14, -7.031029e-15, -8.069868e-15, 
    -1.423019e-14, -6.352333e-15, -1.158637e-14, -1.548893e-14, 
    -1.280142e-14, -3.132848e-15, -9.82224e-15, -1.503771e-14, -8.678556e-15, 
    -1.799875e-14, -7.59897e-15, -1.211594e-14, -1.601215e-14, -1.208239e-14, 
    -6.44776e-15, -8.664055e-15, -1.257149e-14, -1.479615e-14, -9.364859e-15, 
    -1.674433e-14, -2.393323e-14, -6.460655e-15, -9.938682e-15, -9.83873e-15, 
    -1.250787e-14, -1.21317e-14, -1.001311e-14, -4.189343e-15, -1.27979e-14, 
    -1.376826e-14, -2.518157e-14, -1.480849e-14, -6.256081e-15, 
    -1.851933e-14, -1.011767e-14, -1.360335e-14, -7.534211e-15, 
    -1.438116e-14, -1.943114e-14, -8.905268e-15, -9.622656e-15, 
    -8.512967e-15, -7.327104e-16, -8.45307e-15, -1.403814e-14, -1.603479e-14, 
    -2.23026e-14, -1.596875e-14, -1.355606e-14, -1.327863e-14, -1.538694e-14, 
    -4.262757e-15, -1.033418e-14, -1.581461e-14, -5.114715e-15, 
    -8.440787e-15, -2.763371e-14, -2.309445e-14, -6.252664e-15, 
    -1.104798e-14, -1.336699e-14, -2.181876e-14, -5.800311e-15, 
    -1.203703e-14, -4.137943e-15, -8.528241e-15, -1.421621e-14, 
    -1.294809e-14, -1.13539e-14, -1.322957e-14, -1.172355e-14, -5.134428e-15, 
    -1.174636e-14, -7.770769e-15, -1.96013e-14, -1.34465e-14, -1.601443e-14, 
    -1.738559e-14, -1.531285e-14, -1.00234e-14, -1.695297e-14, -1.348923e-14, 
    -8.200628e-15, -1.155416e-14, -6.881518e-15, -1.377802e-14, 
    -8.063187e-15, -1.492782e-14, -1.99862e-14, -2.074638e-14, -8.471722e-15, 
    -1.676662e-14, -2.324246e-14, -1.574076e-14, -8.85916e-15, 2.731787e-16, 
    -1.551246e-14, -3.975589e-15, -2.15708e-14, -2.695193e-14, -8.187341e-15, 
    -3.876666e-15, -1.971292e-14, -1.751515e-14, -9.723228e-15, 
    -1.397164e-14, -1.093385e-14, -1.47359e-14, -1.970822e-14, -1.508498e-14, 
    -1.00471e-14, -3.963401e-15, -1.759893e-14, -1.325693e-14, -1.175693e-14, 
    -1.242106e-14, -1.422721e-14, -1.451393e-14, -7.581672e-15, 
    -2.357592e-14, -1.375516e-14, -1.740398e-14, -8.258171e-15, 
    -1.279306e-14, -1.152855e-14, -2.071323e-14, -1.380216e-14, 
    -1.841574e-14, -1.543548e-14, -1.174562e-14, -1.036164e-14, 
    -1.338821e-14, -1.214372e-14, -5.338177e-15, -9.850072e-15, 
    -8.652206e-15, -1.095896e-14, -1.279129e-14, -1.939448e-14, 
    -1.254443e-14, -1.02092e-14, -1.352248e-14, -1.471459e-14, -1.510893e-14, 
    -9.694047e-15, -1.292222e-14, -2.113545e-14, -1.870657e-14, -1.02525e-14, 
    -9.823969e-15, -1.496084e-14, -2.005968e-14 ;

 ERRSOI =
  -2.283608e-10, -2.267257e-10, -2.613371e-10, -3.844841e-10, -4.593186e-10, 
    -3.167814e-10, -2.717674e-10, -2.89482e-10, -2.751878e-10, -2.652795e-10, 
    -1.971304e-10, -4.041057e-10, -4.189091e-10, -3.455408e-10, 
    -4.879056e-10, -3.994058e-10, -2.386126e-10, -3.117926e-10, -2.64551e-10, 
    -3.647553e-10, -3.766673e-10, -3.319402e-10, -1.629919e-10, 
    -4.471607e-10, -3.039053e-10, -3.34989e-10, -4.176939e-10, -2.679035e-10, 
    -4.388909e-10, -3.01036e-10, -3.277318e-10, -4.840625e-10, -3.089353e-10, 
    -4.920772e-10, -3.594809e-10, -1.705783e-10, -2.786916e-10, -3.9423e-10, 
    -5.285824e-10, -4.030772e-10, -3.040123e-10, -4.452867e-10, 
    -4.841705e-10, -3.517722e-10, -4.220249e-10, -2.968484e-10, 
    -2.569937e-10, -2.97208e-10, -2.906811e-10, -4.073169e-10, -3.012541e-10, 
    -3.260568e-10, -2.890274e-10, -3.794558e-10, -5.055662e-10, 
    -4.034449e-10, -6.150147e-10, -2.654779e-10, -5.070632e-10, 
    -1.223149e-10, -2.948535e-10, -2.388147e-10, -3.24829e-10, -3.271353e-10, 
    -2.12872e-10, -3.137987e-10, -3.947619e-10, -4.0395e-10, -4.370341e-10, 
    -3.236777e-10, -1.694705e-10, -5.958211e-10, -3.792306e-10, 
    -3.599356e-10, -2.484705e-10, -4.14524e-10, -4.352962e-10, -7.72906e-11, 
    -3.919149e-10, -2.961912e-10, -3.578778e-10, -2.818608e-10, 
    -4.190274e-10, -3.405955e-10, -2.905112e-10, -3.871472e-10, 
    -3.321896e-10, -4.060523e-10, -3.608381e-10, -3.045551e-10, -2.92659e-10, 
    -1.740444e-10, -1.916034e-10, -3.400422e-10, -4.043388e-10, 
    -2.182565e-10, -2.458318e-10, -2.597959e-10, -2.150482e-10, 
    -4.742593e-10, -4.197426e-10, -4.94022e-10, -2.91753e-10, -4.42108e-10, 
    -2.935658e-10, -4.373806e-10, -2.678176e-10, -3.036661e-10, 
    -3.641725e-10, -2.241613e-10, -3.832972e-10, -5.799685e-10, 
    -5.561179e-10, -3.788896e-10, -2.886606e-10, -3.355443e-10, 
    -3.909751e-10, -3.105106e-10, -4.763883e-10, -2.70141e-10, -5.080887e-10, 
    -2.53337e-10, -3.734715e-10, -3.576199e-10, -2.483131e-10, -4.611163e-12, 
    -5.420188e-10, -4.148019e-10, -2.348874e-10, -2.786516e-10, -3.55597e-10, 
    -3.391041e-10, -2.185533e-10, -3.845581e-10, -3.899031e-10, -3.68974e-10, 
    -3.304263e-10, -4.67414e-10, -5.541618e-10, -3.716039e-10, -3.434283e-10, 
    -4.345349e-10, -3.022753e-10, -2.292647e-10, -3.840682e-10, 
    -3.948523e-10, -2.562603e-10, -4.58842e-10, -3.227136e-10, -2.238253e-10, 
    -2.135419e-10, -3.130202e-10, -2.148004e-10, -4.374842e-10, 
    -3.949222e-10, -4.935485e-10, -2.378133e-10, -4.23257e-10, -4.875033e-10, 
    -3.870134e-10, -2.59634e-10, -3.80474e-10, -2.416657e-10, -4.065205e-10, 
    -5.16128e-10, -2.924153e-10, -3.977235e-10, -2.368487e-10, -3.455491e-10, 
    -2.550714e-10, -2.754892e-10, -3.613049e-10, -4.29135e-10, -4.697379e-10, 
    -2.984601e-10, -2.104381e-10, -4.296942e-10, -4.585785e-10, 
    -3.509796e-10, -3.224803e-10, -3.306221e-10, -4.495858e-10, 
    -2.204472e-10, -3.51534e-10, -2.657551e-10, -4.908466e-10, -3.642708e-10, 
    -4.01027e-10, -2.670122e-10, -2.835996e-10, -4.290405e-10, -2.849405e-10, 
    -3.033806e-10, -4.57282e-10, -3.151757e-10, -4.427884e-10, -1.741964e-10, 
    -3.205186e-10, -1.648007e-10, -3.894026e-10, -4.064729e-10, 
    -2.022366e-10, -5.663067e-10, -4.489087e-10, -3.120159e-10, 
    -2.474468e-10, -4.505247e-10, -1.99471e-10, -3.694678e-10, -3.124928e-10, 
    -2.639618e-10, -3.372211e-10, -5.458449e-10, -3.375708e-10, 
    -3.174676e-10, -2.299224e-11, -3.537439e-10, -5.411139e-10, 
    -3.033127e-10, -3.646105e-10, -4.163891e-10, -4.571961e-10, 
    -2.121076e-10, -3.065479e-10, -4.490462e-10, -3.743237e-10, 
    -4.065689e-10, -3.660225e-10, -4.146902e-10, -1.812421e-10, 
    -3.284778e-10, -2.794893e-10, -3.74453e-10, -3.30778e-10, -2.904435e-10, 
    -1.856916e-10, -3.371493e-10, -2.210167e-10, -1.822225e-10, 
    -4.264411e-10, -2.926654e-10, -5.631945e-10, -3.091984e-10, 
    -4.019327e-10, -3.261711e-10, -2.755086e-10, -4.286783e-10, 
    -4.425242e-10, -4.749056e-10, -2.876712e-10, -6.52889e-10, -2.126241e-10, 
    -2.351572e-10, -3.219992e-10, -4.575022e-10, -3.782026e-10, 
    -3.802088e-10, -3.803763e-10, -2.122894e-10, -1.118816e-10, 
    -2.288519e-10, -3.480252e-10, -3.884555e-10, -4.328327e-10, 
    -3.785934e-10, -4.239593e-10, -3.063371e-10, -2.166833e-10, 
    -4.040799e-10, -4.185449e-10, -5.875569e-10, -2.614627e-10, 
    -3.749715e-10, -3.421216e-10, -4.000628e-10, -5.713375e-10, 
    -4.648006e-10, -3.285297e-10, -3.588651e-10, -1.751427e-10, -2.53991e-10, 
    -2.721442e-10, -4.076381e-10, -4.890651e-10, -2.309285e-10, 
    -4.225242e-10, -4.930542e-10, -3.803947e-10, -2.497877e-10, 
    -2.965433e-10, -3.482137e-10, -1.745281e-10, -2.697196e-10, 
    -3.310807e-10, -4.180049e-10, -2.557678e-10, -2.95706e-10, -4.180837e-10, 
    -3.410396e-10, -4.074304e-10, -3.024466e-10, -3.87134e-10, -4.707005e-10, 
    -3.301617e-10, -4.141402e-10, -4.637613e-10, -4.614204e-10, 
    -2.633691e-10, -4.021618e-10, -2.9928e-10, -3.202962e-10, -2.389348e-10, 
    -3.281123e-10, -4.562007e-10, -4.582403e-10, -3.44903e-10, -3.732066e-10, 
    -3.617128e-10, -5.442603e-10, -4.790813e-10, -2.580196e-10, 
    -3.204771e-10, -2.283606e-10, -3.516383e-10, -4.126847e-10, 
    -3.096118e-10, -3.48382e-10, -3.534796e-10, -2.118515e-10, -4.416491e-10, 
    -3.914978e-10, -3.100582e-10, -6.514694e-11, -3.689852e-10, 
    -1.304833e-10, -4.898537e-10, -1.892348e-10, -2.871083e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4 =
  1.863407e-16, 1.812636e-16, 1.822508e-16, 1.781551e-16, 1.804273e-16, 
    1.777453e-16, 1.853117e-16, 1.810617e-16, 1.83775e-16, 1.85884e-16, 
    1.70205e-16, 1.779725e-16, 1.621374e-16, 1.670922e-16, 1.546446e-16, 
    1.629081e-16, 1.529781e-16, 1.548837e-16, 1.491493e-16, 1.507923e-16, 
    1.434546e-16, 1.48391e-16, 1.39651e-16, 1.44634e-16, 1.438543e-16, 
    1.485537e-16, 1.7641e-16, 1.711719e-16, 1.767202e-16, 1.759733e-16, 
    1.763086e-16, 1.803802e-16, 1.824314e-16, 1.867291e-16, 1.85949e-16, 
    1.827927e-16, 1.756375e-16, 1.780669e-16, 1.719452e-16, 1.720835e-16, 
    1.652665e-16, 1.683403e-16, 1.568808e-16, 1.601384e-16, 1.507238e-16, 
    1.530917e-16, 1.508349e-16, 1.515193e-16, 1.50826e-16, 1.542988e-16, 
    1.528109e-16, 1.558668e-16, 1.677645e-16, 1.642682e-16, 1.746945e-16, 
    1.809615e-16, 1.851252e-16, 1.880791e-16, 1.876615e-16, 1.868653e-16, 
    1.827743e-16, 1.789282e-16, 1.759967e-16, 1.740356e-16, 1.721033e-16, 
    1.662521e-16, 1.631561e-16, 1.562217e-16, 1.574738e-16, 1.553529e-16, 
    1.533273e-16, 1.499254e-16, 1.504854e-16, 1.489864e-16, 1.554093e-16, 
    1.511406e-16, 1.581869e-16, 1.562599e-16, 1.715757e-16, 1.774117e-16, 
    1.7989e-16, 1.820609e-16, 1.873404e-16, 1.836944e-16, 1.851317e-16, 
    1.817128e-16, 1.795399e-16, 1.806147e-16, 1.73982e-16, 1.765607e-16, 
    1.629726e-16, 1.688261e-16, 1.535636e-16, 1.572169e-16, 1.526879e-16, 
    1.549992e-16, 1.510387e-16, 1.546032e-16, 1.484286e-16, 1.470836e-16, 
    1.480027e-16, 1.444727e-16, 1.548007e-16, 1.508347e-16, 1.806447e-16, 
    1.804694e-16, 1.79653e-16, 1.832416e-16, 1.834613e-16, 1.867504e-16, 
    1.83824e-16, 1.825775e-16, 1.794142e-16, 1.775425e-16, 1.757634e-16, 
    1.718514e-16, 1.674816e-16, 1.613707e-16, 1.569801e-16, 1.540362e-16, 
    1.558416e-16, 1.542477e-16, 1.560294e-16, 1.568645e-16, 1.475874e-16, 
    1.527969e-16, 1.449805e-16, 1.454132e-16, 1.489506e-16, 1.453644e-16, 
    1.803464e-16, 1.81355e-16, 1.848563e-16, 1.821163e-16, 1.871086e-16, 
    1.843139e-16, 1.827068e-16, 1.765063e-16, 1.751444e-16, 1.738808e-16, 
    1.713857e-16, 1.68183e-16, 1.625638e-16, 1.576741e-16, 1.532096e-16, 
    1.535368e-16, 1.534216e-16, 1.524239e-16, 1.548948e-16, 1.520182e-16, 
    1.515352e-16, 1.527978e-16, 1.454711e-16, 1.475645e-16, 1.454223e-16, 
    1.467855e-16, 1.810272e-16, 1.793301e-16, 1.802471e-16, 1.785225e-16, 
    1.797373e-16, 1.743346e-16, 1.727146e-16, 1.65134e-16, 1.682459e-16, 
    1.632938e-16, 1.677431e-16, 1.669546e-16, 1.631313e-16, 1.675028e-16, 
    1.579432e-16, 1.644238e-16, 1.523851e-16, 1.588574e-16, 1.519794e-16, 
    1.532289e-16, 1.511603e-16, 1.493073e-16, 1.469762e-16, 1.426737e-16, 
    1.436702e-16, 1.400719e-16, 1.768e-16, 1.745983e-16, 1.747926e-16, 
    1.724886e-16, 1.707845e-16, 1.670913e-16, 1.611663e-16, 1.633946e-16, 
    1.593042e-16, 1.584828e-16, 1.646974e-16, 1.608815e-16, 1.73125e-16, 
    1.711468e-16, 1.723249e-16, 1.766261e-16, 1.628806e-16, 1.699352e-16, 
    1.569074e-16, 1.607302e-16, 1.495714e-16, 1.551212e-16, 1.442186e-16, 
    1.395549e-16, 1.351667e-16, 1.300347e-16, 1.733971e-16, 1.748931e-16, 
    1.722147e-16, 1.68508e-16, 1.650695e-16, 1.60497e-16, 1.600294e-16, 
    1.591725e-16, 1.569535e-16, 1.550872e-16, 1.589012e-16, 1.546194e-16, 
    1.706871e-16, 1.622684e-16, 1.754583e-16, 1.714865e-16, 1.687267e-16, 
    1.699378e-16, 1.636494e-16, 1.62167e-16, 1.561419e-16, 1.59257e-16, 
    1.407057e-16, 1.489152e-16, 1.261276e-16, 1.324984e-16, 1.754157e-16, 
    1.734024e-16, 1.66394e-16, 1.697289e-16, 1.60192e-16, 1.578438e-16, 
    1.559351e-16, 1.534941e-16, 1.532309e-16, 1.517845e-16, 1.541545e-16, 
    1.518783e-16, 1.604873e-16, 1.566407e-16, 1.671957e-16, 1.646268e-16, 
    1.658088e-16, 1.671049e-16, 1.631044e-16, 1.58841e-16, 1.587506e-16, 
    1.573833e-16, 1.535284e-16, 1.601533e-16, 1.396446e-16, 1.523114e-16, 
    1.712069e-16, 1.673275e-16, 1.667742e-16, 1.682769e-16, 1.580792e-16, 
    1.617745e-16, 1.518199e-16, 1.545109e-16, 1.501017e-16, 1.522928e-16, 
    1.526151e-16, 1.55429e-16, 1.571805e-16, 1.61605e-16, 1.652046e-16, 
    1.68059e-16, 1.673954e-16, 1.642598e-16, 1.585804e-16, 1.532067e-16, 
    1.543839e-16, 1.504368e-16, 1.608835e-16, 1.565034e-16, 1.581962e-16, 
    1.53782e-16, 1.634537e-16, 1.552159e-16, 1.655587e-16, 1.646522e-16, 
    1.618479e-16, 1.562058e-16, 1.549583e-16, 1.53625e-16, 1.544479e-16, 
    1.584363e-16, 1.5909e-16, 1.619162e-16, 1.626961e-16, 1.648496e-16, 
    1.66632e-16, 1.650033e-16, 1.632926e-16, 1.584349e-16, 1.540559e-16, 
    1.492808e-16, 1.481123e-16, 1.425297e-16, 1.470733e-16, 1.395739e-16, 
    1.459485e-16, 1.34913e-16, 1.547394e-16, 1.461374e-16, 1.617205e-16, 
    1.600424e-16, 1.570062e-16, 1.500421e-16, 1.538028e-16, 1.494049e-16, 
    1.591156e-16, 1.641512e-16, 1.654548e-16, 1.678854e-16, 1.653992e-16, 
    1.656015e-16, 1.632223e-16, 1.639869e-16, 1.582736e-16, 1.613427e-16, 
    1.52623e-16, 1.494398e-16, 1.404488e-16, 1.349345e-16, 1.293207e-16, 
    1.268414e-16, 1.260867e-16, 1.257712e-16 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  23.77457, 23.83677, 23.82469, 23.87484, 23.84705, 23.87987, 23.78721, 
    23.8392, 23.80603, 23.78022, 23.97214, 23.87709, 24.07142, 24.01063, 
    24.16357, 24.0619, 24.1841, 24.16073, 24.23133, 24.21111, 24.30128, 
    24.24067, 24.34822, 24.28685, 24.29641, 24.23866, 23.8963, 23.96027, 
    23.89249, 23.90161, 23.89754, 23.84759, 23.82237, 23.76989, 23.77943, 
    23.81802, 23.90572, 23.876, 23.95111, 23.94942, 24.03307, 23.99534, 
    24.13616, 24.09613, 24.21195, 24.18279, 24.21056, 24.20215, 24.21067, 
    24.16792, 24.18623, 24.14865, 24.00238, 24.04531, 23.91731, 23.84033, 
    23.78948, 23.75335, 23.75846, 23.76817, 23.81824, 23.86544, 23.9014, 
    23.92545, 23.94917, 24.02077, 24.0589, 24.14421, 24.12889, 24.15491, 
    24.1799, 24.22175, 24.21487, 24.2333, 24.15428, 24.20676, 24.12015, 
    24.14381, 23.95529, 23.88403, 23.85348, 23.827, 23.76238, 23.80698, 
    23.78938, 23.83132, 23.85793, 23.84478, 23.92611, 23.89447, 24.06116, 
    23.98932, 24.17698, 24.13204, 24.18777, 24.15934, 24.20803, 24.16421, 
    24.24018, 24.2567, 24.2454, 24.28891, 24.16177, 24.21053, 23.8444, 
    23.84654, 23.85656, 23.81252, 23.80984, 23.76961, 23.80544, 23.82067, 
    23.8595, 23.88242, 23.90423, 23.95223, 24.00581, 24.0809, 24.13495, 
    24.17119, 24.14899, 24.16858, 24.14667, 24.13641, 24.25049, 24.18638, 
    24.28265, 24.27733, 24.23372, 24.27793, 23.84805, 23.83571, 23.79278, 
    23.82638, 23.76523, 23.79941, 23.81904, 23.89506, 23.91185, 23.92732, 
    23.95796, 23.99727, 24.06625, 24.12638, 24.18136, 24.17734, 24.17875, 
    24.19101, 24.16061, 24.196, 24.20191, 24.18641, 24.27661, 24.25084, 
    24.27721, 24.26044, 23.83973, 23.86051, 23.84928, 23.87039, 23.85549, 
    23.92167, 23.94153, 24.03461, 23.99647, 24.05726, 24.00267, 24.01232, 
    24.05911, 24.00564, 24.123, 24.04329, 24.19148, 24.11168, 24.19648, 
    24.18112, 24.20658, 24.22935, 24.25808, 24.311, 24.29875, 24.34309, 
    23.89154, 23.91848, 23.91617, 23.94443, 23.96531, 24.01069, 24.08346, 
    24.0561, 24.10639, 24.11647, 24.04011, 24.08693, 23.93657, 23.96078, 
    23.94641, 23.89363, 24.06232, 23.97566, 24.13583, 24.08883, 24.2261, 
    24.15774, 24.292, 24.34931, 24.40357, 24.4667, 23.93326, 23.91494, 
    23.9478, 23.99319, 24.0355, 24.09169, 24.09747, 24.10799, 24.13531, 
    24.15825, 24.11125, 24.16401, 23.96627, 24.06988, 23.90796, 23.95659, 
    23.99054, 23.97571, 24.05299, 24.0712, 24.14521, 24.10698, 24.3351, 
    24.23408, 24.515, 24.43635, 23.90852, 23.93323, 24.01918, 23.97828, 
    24.09547, 24.12432, 24.14784, 24.17781, 24.18109, 24.19886, 24.16973, 
    24.19773, 24.09181, 24.13913, 24.00943, 24.04094, 24.02646, 24.01054, 
    24.05968, 24.11198, 24.1132, 24.12995, 24.17702, 24.09595, 24.34797, 
    24.19205, 23.96017, 24.00766, 24.01457, 23.99614, 24.12143, 24.07599, 
    24.19844, 24.16535, 24.2196, 24.19263, 24.18866, 24.15405, 24.13249, 
    24.07806, 24.03383, 23.99883, 24.00697, 24.04543, 24.1152, 24.18134, 
    24.16683, 24.21548, 24.08697, 24.14077, 24.11994, 24.1743, 24.05536, 
    24.15633, 24.02953, 24.04066, 24.07509, 24.14436, 24.15984, 24.1762, 
    24.16612, 24.11699, 24.10899, 24.07428, 24.06465, 24.03825, 24.01635, 
    24.03633, 24.0573, 24.11705, 24.17089, 24.22966, 24.24409, 24.31259, 
    24.25669, 24.34882, 24.27028, 24.40639, 24.16233, 24.26817, 24.07669, 
    24.09732, 24.13454, 24.22019, 24.17404, 24.22806, 24.10868, 24.04671, 
    24.0308, 24.00094, 24.03148, 24.029, 24.05824, 24.04885, 24.11904, 
    24.08133, 24.18853, 24.22766, 24.33841, 24.40631, 24.47566, 24.50624, 
    24.51556, 24.51945 ;

 FGR =
  -426.9097, -427.9266, -427.7291, -428.5489, -428.0944, -428.631, -427.1161, 
    -427.9667, -427.4239, -427.0016, -430.1389, -428.5856, -431.7549, 
    -430.764, -433.2536, -431.6003, -433.587, -433.2066, -434.3532, 
    -434.0248, -435.4895, -434.5048, -436.2497, -435.2548, -435.4102, 
    -434.4722, -428.8988, -429.9453, -428.8367, -428.986, -428.9191, 
    -428.1035, -427.6921, -426.8324, -426.9886, -427.6203, -429.0531, 
    -428.5672, -429.7931, -429.7654, -431.1295, -430.5145, -432.8072, 
    -432.1558, -434.0385, -433.565, -434.0161, -433.8794, -434.0179, 
    -433.3235, -433.621, -433.0101, -430.6295, -431.329, -429.2421, 
    -427.9861, -427.1533, -426.5619, -426.6455, -426.8047, -427.624, 
    -428.3947, -428.9818, -429.3745, -429.7614, -430.9308, -431.5511, 
    -432.9386, -432.6888, -433.1124, -433.5179, -434.1978, -434.086, 
    -434.3854, -433.1017, -433.9547, -432.5464, -432.9315, -429.8643, 
    -428.6984, -428.2008, -427.767, -426.7097, -427.4397, -427.1519, 
    -427.8371, -428.2722, -428.0571, -429.3852, -428.8688, -431.5878, 
    -430.4168, -433.4706, -432.7401, -433.6458, -433.1838, -433.9752, 
    -433.2629, -434.497, -434.7654, -434.582, -435.2875, -433.2234, 
    -434.0159, -428.051, -428.086, -428.2496, -427.5304, -427.4865, -426.828, 
    -427.4141, -427.6635, -428.2975, -428.6721, -429.0284, -429.8116, 
    -430.6858, -431.9087, -432.7874, -433.3763, -433.0154, -433.334, 
    -432.9777, -432.8108, -434.6647, -433.6236, -435.186, -435.0997, 
    -434.3925, -435.1094, -428.1107, -427.9088, -427.2073, -427.7563, 
    -426.7563, -427.3158, -427.6373, -428.8791, -429.1525, -429.4052, 
    -429.9049, -430.5459, -431.6701, -432.6483, -433.5416, -433.4762, 
    -433.4992, -433.6985, -433.2045, -433.7796, -433.8759, -433.6238, 
    -435.0881, -434.6698, -435.0978, -434.8256, -427.9745, -428.3142, 
    -428.1306, -428.4758, -428.2324, -429.3138, -429.6379, -431.1553, 
    -430.5332, -431.5239, -430.634, -430.7916, -431.5552, -430.6823, 
    -432.594, -431.2971, -433.7062, -432.4105, -433.7874, -433.5377, 
    -433.9513, -434.3214, -434.7874, -435.6463, -435.4475, -436.1661, 
    -428.8209, -429.2613, -429.223, -429.6841, -430.0251, -430.7646, 
    -431.9499, -431.5043, -432.3228, -432.4869, -431.2437, -432.0066, 
    -429.5564, -429.9519, -429.7167, -428.8554, -431.6064, -430.1945, 
    -432.8019, -432.0373, -434.2685, -433.1586, -435.338, -436.2682, 
    -437.1454, -438.168, -429.5021, -429.2029, -429.7391, -430.4802, 
    -431.1689, -432.0838, -432.1776, -432.3489, -432.793, -433.1661, 
    -432.4026, -433.2597, -430.0428, -431.7291, -429.0893, -429.8837, 
    -430.4367, -430.1946, -431.4535, -431.75, -432.9547, -432.3322, 
    -436.0382, -434.3989, -438.9479, -437.6769, -429.0982, -429.5013, 
    -430.9036, -430.2365, -432.1451, -432.6147, -432.9967, -433.4843, 
    -433.5372, -433.8262, -433.3527, -433.8076, -432.0858, -432.8554, 
    -430.7438, -431.2576, -431.0214, -430.762, -431.5625, -432.4146, 
    -432.4334, -432.7065, -433.4747, -432.1529, -436.2484, -433.7184, 
    -429.9408, -430.7163, -430.8279, -430.5273, -432.5675, -431.8283, 
    -433.8192, -433.2814, -434.1628, -433.7248, -433.6603, -433.0978, 
    -432.7474, -431.8621, -431.1418, -430.571, -430.7038, -431.3308, 
    -432.4668, -433.5417, -433.3062, -434.0958, -432.0067, -432.8825, 
    -432.5438, -433.427, -431.4923, -433.1377, -431.0714, -431.2528, 
    -431.8136, -432.9414, -433.1919, -433.4581, -433.294, -432.4958, 
    -432.3653, -431.8002, -431.6438, -431.2133, -430.8566, -431.1824, 
    -431.5243, -432.4964, -433.3719, -434.3265, -434.5604, -435.6736, 
    -434.7665, -436.2624, -434.9892, -437.1937, -433.2341, -434.9531, 
    -431.8394, -432.1751, -432.7815, -434.1736, -433.4228, -434.3011, 
    -432.3603, -431.3521, -431.0921, -430.6056, -431.1033, -431.0628, 
    -431.5389, -431.386, -432.5287, -431.9149, -433.6585, -434.2944, 
    -436.0906, -437.1908, -438.3116, -438.8059, -438.9564, -439.0193 ;

 FGR12 =
  -127.4534, -127.5083, -127.4977, -127.5421, -127.5175, -127.5466, 
    -127.4646, -127.5105, -127.4812, -127.4584, -127.6288, -127.5441, 
    -127.7183, -127.6636, -127.8017, -127.7097, -127.8204, -127.7993, 
    -127.8636, -127.8451, -127.9274, -127.8721, -127.9705, -127.9143, 
    -127.923, -127.8703, -127.5613, -127.6182, -127.5579, -127.566, 
    -127.5623, -127.518, -127.4955, -127.4493, -127.4577, -127.4917, 
    -127.5696, -127.5432, -127.6102, -127.6087, -127.6838, -127.6499, 
    -127.7769, -127.7407, -127.8459, -127.8193, -127.8446, -127.837, 
    -127.8447, -127.8058, -127.8224, -127.7883, -127.6562, -127.6947, 
    -127.58, -127.5114, -127.4665, -127.4347, -127.4392, -127.4478, -127.492, 
    -127.5338, -127.5658, -127.5873, -127.6085, -127.6725, -127.707, 
    -127.7842, -127.7704, -127.7939, -127.8167, -127.8548, -127.8486, 
    -127.8653, -127.7934, -127.8411, -127.7625, -127.7839, -127.6137, 
    -127.5503, -127.5231, -127.4997, -127.4427, -127.482, -127.4665, 
    -127.5036, -127.5271, -127.5155, -127.5879, -127.5596, -127.709, 
    -127.6444, -127.814, -127.7732, -127.8239, -127.798, -127.8423, 
    -127.8025, -127.8717, -127.8867, -127.8764, -127.9162, -127.8002, 
    -127.8446, -127.5152, -127.5171, -127.5259, -127.4869, -127.4845, 
    -127.4491, -127.4807, -127.4941, -127.5285, -127.5489, -127.5683, 
    -127.6112, -127.6592, -127.7269, -127.7759, -127.8088, -127.7886, 
    -127.8064, -127.7865, -127.7772, -127.881, -127.8226, -127.9105, 
    -127.9056, -127.8658, -127.9062, -127.5184, -127.5075, -127.4695, 
    -127.4992, -127.4452, -127.4753, -127.4927, -127.5601, -127.5752, 
    -127.5889, -127.6164, -127.6516, -127.7137, -127.768, -127.818, 
    -127.8144, -127.8157, -127.8268, -127.7992, -127.8313, -127.8367, 
    -127.8226, -127.905, -127.8814, -127.9055, -127.8902, -127.511, 
    -127.5294, -127.5195, -127.5382, -127.525, -127.5838, -127.6016, 
    -127.6851, -127.6509, -127.7055, -127.6565, -127.6651, -127.7071, 
    -127.6591, -127.7649, -127.6929, -127.8272, -127.7547, -127.8318, 
    -127.8178, -127.841, -127.8618, -127.888, -127.9364, -127.9252, 
    -127.9659, -127.557, -127.581, -127.579, -127.6042, -127.6229, -127.6637, 
    -127.7292, -127.7046, -127.75, -127.7591, -127.6902, -127.7323, 
    -127.5972, -127.6188, -127.606, -127.5589, -127.7101, -127.6322, 
    -127.7766, -127.7341, -127.8588, -127.7965, -127.919, -127.9715, 
    -128.0216, -128.0799, -127.5942, -127.5779, -127.6073, -127.6479, 
    -127.686, -127.7367, -127.7419, -127.7514, -127.7762, -127.797, 
    -127.7543, -127.8022, -127.6236, -127.7169, -127.5717, -127.615, 
    -127.6455, -127.6322, -127.7018, -127.7182, -127.7851, -127.7505, 
    -127.9584, -127.866, -128.1248, -128.0518, -127.5722, -127.5943, 
    -127.6712, -127.6346, -127.7401, -127.7662, -127.7876, -127.8148, 
    -127.8178, -127.8339, -127.8075, -127.8329, -127.7368, -127.7796, 
    -127.6626, -127.6909, -127.6779, -127.6636, -127.7078, -127.755, 
    -127.7562, -127.7713, -127.8138, -127.7406, -127.9701, -127.8276, 
    -127.6184, -127.6608, -127.6671, -127.6506, -127.7636, -127.7225, 
    -127.8336, -127.8035, -127.8529, -127.8283, -127.8247, -127.7932, 
    -127.7736, -127.7244, -127.6845, -127.653, -127.6604, -127.6949, 
    -127.7579, -127.818, -127.8048, -127.8491, -127.7325, -127.7811, 
    -127.7622, -127.8116, -127.7039, -127.795, -127.6806, -127.6907, 
    -127.7217, -127.7843, -127.7985, -127.8133, -127.8042, -127.7596, 
    -127.7523, -127.721, -127.7122, -127.6885, -127.6688, -127.6867, 
    -127.7056, -127.7596, -127.8085, -127.862, -127.8753, -127.9377, 
    -127.8866, -127.9708, -127.8989, -128.024, -127.8006, -127.897, 
    -127.7232, -127.7418, -127.7754, -127.8533, -127.8114, -127.8605, 
    -127.7521, -127.696, -127.6818, -127.6549, -127.6824, -127.6802, 
    -127.7065, -127.698, -127.7614, -127.7274, -127.8245, -127.8602, 
    -127.9616, -128.024, -128.0883, -128.1167, -128.1254, -128.129 ;

 FGR_R =
  -426.9097, -427.9266, -427.7291, -428.5489, -428.0944, -428.631, -427.1161, 
    -427.9667, -427.4239, -427.0016, -430.1389, -428.5856, -431.7549, 
    -430.764, -433.2536, -431.6003, -433.587, -433.2066, -434.3532, 
    -434.0248, -435.4895, -434.5048, -436.2497, -435.2548, -435.4102, 
    -434.4722, -428.8988, -429.9453, -428.8367, -428.986, -428.9191, 
    -428.1035, -427.6921, -426.8324, -426.9886, -427.6203, -429.0531, 
    -428.5672, -429.7931, -429.7654, -431.1295, -430.5145, -432.8072, 
    -432.1558, -434.0385, -433.565, -434.0161, -433.8794, -434.0179, 
    -433.3235, -433.621, -433.0101, -430.6295, -431.329, -429.2421, 
    -427.9861, -427.1533, -426.5619, -426.6455, -426.8047, -427.624, 
    -428.3947, -428.9818, -429.3745, -429.7614, -430.9308, -431.5511, 
    -432.9386, -432.6888, -433.1124, -433.5179, -434.1978, -434.086, 
    -434.3854, -433.1017, -433.9547, -432.5464, -432.9315, -429.8643, 
    -428.6984, -428.2008, -427.767, -426.7097, -427.4397, -427.1519, 
    -427.8371, -428.2722, -428.0571, -429.3852, -428.8688, -431.5878, 
    -430.4168, -433.4706, -432.7401, -433.6458, -433.1838, -433.9752, 
    -433.2629, -434.497, -434.7654, -434.582, -435.2875, -433.2234, 
    -434.0159, -428.051, -428.086, -428.2496, -427.5304, -427.4865, -426.828, 
    -427.4141, -427.6635, -428.2975, -428.6721, -429.0284, -429.8116, 
    -430.6858, -431.9087, -432.7874, -433.3763, -433.0154, -433.334, 
    -432.9777, -432.8108, -434.6647, -433.6236, -435.186, -435.0997, 
    -434.3925, -435.1094, -428.1107, -427.9088, -427.2073, -427.7563, 
    -426.7563, -427.3158, -427.6373, -428.8791, -429.1525, -429.4052, 
    -429.9049, -430.5459, -431.6701, -432.6483, -433.5416, -433.4762, 
    -433.4992, -433.6985, -433.2045, -433.7796, -433.8759, -433.6238, 
    -435.0881, -434.6698, -435.0978, -434.8256, -427.9745, -428.3142, 
    -428.1306, -428.4758, -428.2324, -429.3138, -429.6379, -431.1553, 
    -430.5332, -431.5239, -430.634, -430.7916, -431.5552, -430.6823, 
    -432.594, -431.2971, -433.7062, -432.4105, -433.7874, -433.5377, 
    -433.9513, -434.3214, -434.7874, -435.6463, -435.4475, -436.1661, 
    -428.8209, -429.2613, -429.223, -429.6841, -430.0251, -430.7646, 
    -431.9499, -431.5043, -432.3228, -432.4869, -431.2437, -432.0066, 
    -429.5564, -429.9519, -429.7167, -428.8554, -431.6064, -430.1945, 
    -432.8019, -432.0373, -434.2685, -433.1586, -435.338, -436.2682, 
    -437.1454, -438.168, -429.5021, -429.2029, -429.7391, -430.4802, 
    -431.1689, -432.0838, -432.1776, -432.3489, -432.793, -433.1661, 
    -432.4026, -433.2597, -430.0428, -431.7291, -429.0893, -429.8837, 
    -430.4367, -430.1946, -431.4535, -431.75, -432.9547, -432.3322, 
    -436.0382, -434.3989, -438.9479, -437.6769, -429.0982, -429.5013, 
    -430.9036, -430.2365, -432.1451, -432.6147, -432.9967, -433.4843, 
    -433.5372, -433.8262, -433.3527, -433.8076, -432.0858, -432.8554, 
    -430.7438, -431.2576, -431.0214, -430.762, -431.5625, -432.4146, 
    -432.4334, -432.7065, -433.4747, -432.1529, -436.2484, -433.7184, 
    -429.9408, -430.7163, -430.8279, -430.5273, -432.5675, -431.8283, 
    -433.8192, -433.2814, -434.1628, -433.7248, -433.6603, -433.0978, 
    -432.7474, -431.8621, -431.1418, -430.571, -430.7038, -431.3308, 
    -432.4668, -433.5417, -433.3062, -434.0958, -432.0067, -432.8825, 
    -432.5438, -433.427, -431.4923, -433.1377, -431.0714, -431.2528, 
    -431.8136, -432.9414, -433.1919, -433.4581, -433.294, -432.4958, 
    -432.3653, -431.8002, -431.6438, -431.2133, -430.8566, -431.1824, 
    -431.5243, -432.4964, -433.3719, -434.3265, -434.5604, -435.6736, 
    -434.7665, -436.2624, -434.9892, -437.1937, -433.2341, -434.9531, 
    -431.8394, -432.1751, -432.7815, -434.1736, -433.4228, -434.3011, 
    -432.3603, -431.3521, -431.0921, -430.6056, -431.1033, -431.0628, 
    -431.5389, -431.386, -432.5287, -431.9149, -433.6585, -434.2944, 
    -436.0906, -437.1908, -438.3116, -438.8059, -438.9564, -439.0193 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  49.00589, 49.07697, 49.06317, 49.12046, 49.0887, 49.1262, 49.02033, 
    49.07978, 49.04184, 49.01233, 49.23157, 49.12303, 49.3445, 49.27526, 
    49.44923, 49.3337, 49.47253, 49.44595, 49.52608, 49.50313, 49.60547, 
    49.53667, 49.6586, 49.58907, 49.59993, 49.53439, 49.14492, 49.21804, 
    49.14058, 49.151, 49.14634, 49.08934, 49.06058, 49.0005, 49.01141, 
    49.05556, 49.1557, 49.12174, 49.20741, 49.20548, 49.3008, 49.25783, 
    49.41805, 49.37253, 49.50409, 49.471, 49.50252, 49.49297, 49.50265, 
    49.45412, 49.47491, 49.43222, 49.26587, 49.31475, 49.16891, 49.08112, 
    49.02293, 48.98159, 48.98743, 48.99856, 49.05582, 49.10969, 49.15072, 
    49.17816, 49.2052, 49.28691, 49.33026, 49.42722, 49.40977, 49.43937, 
    49.46771, 49.51522, 49.50741, 49.52833, 49.43862, 49.49823, 49.39982, 
    49.42673, 49.21238, 49.13091, 49.09613, 49.06582, 48.99192, 49.04294, 
    49.02283, 49.07072, 49.10112, 49.0861, 49.17891, 49.14282, 49.33282, 
    49.251, 49.4644, 49.41336, 49.47664, 49.44436, 49.49966, 49.44989, 
    49.53613, 49.55488, 49.54206, 49.59136, 49.44713, 49.50251, 49.08567, 
    49.08812, 49.09955, 49.04928, 49.04621, 49.00019, 49.04116, 49.05859, 
    49.1029, 49.12908, 49.15397, 49.20871, 49.26979, 49.35525, 49.41666, 
    49.45781, 49.43259, 49.45486, 49.42996, 49.4183, 49.54784, 49.47509, 
    49.58427, 49.57824, 49.52882, 49.57892, 49.08984, 49.07573, 49.0267, 
    49.06507, 48.99517, 49.03428, 49.05675, 49.14354, 49.16265, 49.18031, 
    49.21523, 49.26003, 49.33858, 49.40694, 49.46936, 49.46479, 49.4664, 
    49.48033, 49.44581, 49.48599, 49.49272, 49.47511, 49.57743, 49.5482, 
    49.57811, 49.55909, 49.08033, 49.10406, 49.09124, 49.11535, 49.09835, 
    49.17391, 49.19657, 49.3026, 49.25913, 49.32836, 49.26618, 49.27719, 
    49.33054, 49.26955, 49.40314, 49.31251, 49.48087, 49.39032, 49.48654, 
    49.46909, 49.49799, 49.52385, 49.55641, 49.61643, 49.60254, 49.65276, 
    49.13948, 49.17025, 49.16757, 49.1998, 49.22363, 49.2753, 49.35814, 
    49.327, 49.38419, 49.39566, 49.30879, 49.3621, 49.19087, 49.21851, 
    49.20208, 49.14188, 49.33413, 49.23546, 49.41767, 49.36424, 49.52016, 
    49.44259, 49.59489, 49.65988, 49.72118, 49.79263, 49.18708, 49.16617, 
    49.20364, 49.25542, 49.30356, 49.36749, 49.37405, 49.38602, 49.41705, 
    49.44313, 49.38977, 49.44967, 49.22485, 49.3427, 49.15823, 49.21375, 
    49.25239, 49.23547, 49.32345, 49.34417, 49.42835, 49.38485, 49.64381, 
    49.52927, 49.84713, 49.75832, 49.15885, 49.18702, 49.28502, 49.2384, 
    49.37178, 49.40459, 49.43129, 49.46535, 49.46906, 49.48925, 49.45616, 
    49.48795, 49.36763, 49.42141, 49.27385, 49.30975, 49.29325, 49.27512, 
    49.33107, 49.3906, 49.39193, 49.41101, 49.46467, 49.37232, 49.65849, 
    49.4817, 49.21774, 49.27192, 49.27973, 49.25873, 49.4013, 49.34964, 
    49.48877, 49.45118, 49.51277, 49.48216, 49.47766, 49.43835, 49.41386, 
    49.352, 49.30167, 49.26178, 49.27106, 49.31488, 49.39426, 49.46937, 
    49.45291, 49.50809, 49.36211, 49.4233, 49.39964, 49.46135, 49.32616, 
    49.44112, 49.29675, 49.30942, 49.34861, 49.42741, 49.44493, 49.46353, 
    49.45206, 49.39628, 49.38717, 49.34768, 49.33674, 49.30667, 49.28174, 
    49.3045, 49.32839, 49.39632, 49.4575, 49.52421, 49.54055, 49.61833, 
    49.55495, 49.65947, 49.5705, 49.72454, 49.44787, 49.56799, 49.35041, 
    49.37387, 49.41624, 49.51352, 49.46106, 49.52243, 49.38681, 49.31636, 
    49.29819, 49.26419, 49.29897, 49.29615, 49.32942, 49.31873, 49.39858, 
    49.35569, 49.47753, 49.52197, 49.64747, 49.72435, 49.80267, 49.83721, 
    49.84772, 49.85212 ;

 FIRA_R =
  49.00589, 49.07697, 49.06317, 49.12046, 49.0887, 49.1262, 49.02033, 
    49.07978, 49.04184, 49.01233, 49.23157, 49.12303, 49.3445, 49.27526, 
    49.44923, 49.3337, 49.47253, 49.44595, 49.52608, 49.50313, 49.60547, 
    49.53667, 49.6586, 49.58907, 49.59993, 49.53439, 49.14492, 49.21804, 
    49.14058, 49.151, 49.14634, 49.08934, 49.06058, 49.0005, 49.01141, 
    49.05556, 49.1557, 49.12174, 49.20741, 49.20548, 49.3008, 49.25783, 
    49.41805, 49.37253, 49.50409, 49.471, 49.50252, 49.49297, 49.50265, 
    49.45412, 49.47491, 49.43222, 49.26587, 49.31475, 49.16891, 49.08112, 
    49.02293, 48.98159, 48.98743, 48.99856, 49.05582, 49.10969, 49.15072, 
    49.17816, 49.2052, 49.28691, 49.33026, 49.42722, 49.40977, 49.43937, 
    49.46771, 49.51522, 49.50741, 49.52833, 49.43862, 49.49823, 49.39982, 
    49.42673, 49.21238, 49.13091, 49.09613, 49.06582, 48.99192, 49.04294, 
    49.02283, 49.07072, 49.10112, 49.0861, 49.17891, 49.14282, 49.33282, 
    49.251, 49.4644, 49.41336, 49.47664, 49.44436, 49.49966, 49.44989, 
    49.53613, 49.55488, 49.54206, 49.59136, 49.44713, 49.50251, 49.08567, 
    49.08812, 49.09955, 49.04928, 49.04621, 49.00019, 49.04116, 49.05859, 
    49.1029, 49.12908, 49.15397, 49.20871, 49.26979, 49.35525, 49.41666, 
    49.45781, 49.43259, 49.45486, 49.42996, 49.4183, 49.54784, 49.47509, 
    49.58427, 49.57824, 49.52882, 49.57892, 49.08984, 49.07573, 49.0267, 
    49.06507, 48.99517, 49.03428, 49.05675, 49.14354, 49.16265, 49.18031, 
    49.21523, 49.26003, 49.33858, 49.40694, 49.46936, 49.46479, 49.4664, 
    49.48033, 49.44581, 49.48599, 49.49272, 49.47511, 49.57743, 49.5482, 
    49.57811, 49.55909, 49.08033, 49.10406, 49.09124, 49.11535, 49.09835, 
    49.17391, 49.19657, 49.3026, 49.25913, 49.32836, 49.26618, 49.27719, 
    49.33054, 49.26955, 49.40314, 49.31251, 49.48087, 49.39032, 49.48654, 
    49.46909, 49.49799, 49.52385, 49.55641, 49.61643, 49.60254, 49.65276, 
    49.13948, 49.17025, 49.16757, 49.1998, 49.22363, 49.2753, 49.35814, 
    49.327, 49.38419, 49.39566, 49.30879, 49.3621, 49.19087, 49.21851, 
    49.20208, 49.14188, 49.33413, 49.23546, 49.41767, 49.36424, 49.52016, 
    49.44259, 49.59489, 49.65988, 49.72118, 49.79263, 49.18708, 49.16617, 
    49.20364, 49.25542, 49.30356, 49.36749, 49.37405, 49.38602, 49.41705, 
    49.44313, 49.38977, 49.44967, 49.22485, 49.3427, 49.15823, 49.21375, 
    49.25239, 49.23547, 49.32345, 49.34417, 49.42835, 49.38485, 49.64381, 
    49.52927, 49.84713, 49.75832, 49.15885, 49.18702, 49.28502, 49.2384, 
    49.37178, 49.40459, 49.43129, 49.46535, 49.46906, 49.48925, 49.45616, 
    49.48795, 49.36763, 49.42141, 49.27385, 49.30975, 49.29325, 49.27512, 
    49.33107, 49.3906, 49.39193, 49.41101, 49.46467, 49.37232, 49.65849, 
    49.4817, 49.21774, 49.27192, 49.27973, 49.25873, 49.4013, 49.34964, 
    49.48877, 49.45118, 49.51277, 49.48216, 49.47766, 49.43835, 49.41386, 
    49.352, 49.30167, 49.26178, 49.27106, 49.31488, 49.39426, 49.46937, 
    49.45291, 49.50809, 49.36211, 49.4233, 49.39964, 49.46135, 49.32616, 
    49.44112, 49.29675, 49.30942, 49.34861, 49.42741, 49.44493, 49.46353, 
    49.45206, 49.39628, 49.38717, 49.34768, 49.33674, 49.30667, 49.28174, 
    49.3045, 49.32839, 49.39632, 49.4575, 49.52421, 49.54055, 49.61833, 
    49.55495, 49.65947, 49.5705, 49.72454, 49.44787, 49.56799, 49.35041, 
    49.37387, 49.41624, 49.51352, 49.46106, 49.52243, 49.38681, 49.31636, 
    49.29819, 49.26419, 49.29897, 49.29615, 49.32942, 49.31873, 49.39858, 
    49.35569, 49.47753, 49.52197, 49.64747, 49.72435, 49.80267, 49.83721, 
    49.84772, 49.85212 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  263.3521, 263.4231, 263.4093, 263.4666, 263.4348, 263.4724, 263.3665, 
    263.4259, 263.388, 263.3585, 263.5777, 263.4692, 263.6906, 263.6214, 
    263.7954, 263.6798, 263.8187, 263.7921, 263.8722, 263.8493, 263.9516, 
    263.8828, 264.0047, 263.9352, 263.9461, 263.8805, 263.4911, 263.5642, 
    263.4867, 263.4972, 263.4925, 263.4355, 263.4067, 263.3466, 263.3575, 
    263.4017, 263.5018, 263.4679, 263.5536, 263.5516, 263.6469, 263.604, 
    263.7642, 263.7187, 263.8502, 263.8171, 263.8487, 263.8391, 263.8488, 
    263.8003, 263.821, 263.7784, 263.612, 263.6609, 263.515, 263.4273, 
    263.3691, 263.3277, 263.3336, 263.3447, 263.402, 263.4558, 263.4969, 
    263.5243, 263.5514, 263.6331, 263.6764, 263.7734, 263.7559, 263.7855, 
    263.8138, 263.8614, 263.8535, 263.8745, 263.7848, 263.8444, 263.746, 
    263.7729, 263.5585, 263.4771, 263.4423, 263.412, 263.3381, 263.3891, 
    263.369, 263.4169, 263.4473, 263.4323, 263.5251, 263.489, 263.679, 
    263.5971, 263.8105, 263.7595, 263.8228, 263.7905, 263.8458, 263.796, 
    263.8823, 263.901, 263.8882, 263.9375, 263.7933, 263.8487, 263.4318, 
    263.4343, 263.4457, 263.3954, 263.3924, 263.3463, 263.3873, 263.4047, 
    263.449, 263.4752, 263.5001, 263.5548, 263.6159, 263.7014, 263.7628, 
    263.804, 263.7787, 263.801, 263.7761, 263.7644, 263.894, 263.8212, 
    263.9304, 263.9244, 263.875, 263.925, 263.436, 263.4219, 263.3728, 
    263.4112, 263.3413, 263.3804, 263.4029, 263.4897, 263.5088, 263.5265, 
    263.5614, 263.6062, 263.6847, 263.7531, 263.8155, 263.8109, 263.8125, 
    263.8265, 263.792, 263.8321, 263.8389, 263.8213, 263.9236, 263.8943, 
    263.9243, 263.9052, 263.4265, 263.4502, 263.4374, 263.4615, 263.4445, 
    263.5201, 263.5427, 263.6487, 263.6053, 263.6745, 263.6123, 263.6233, 
    263.6767, 263.6157, 263.7493, 263.6587, 263.827, 263.7365, 263.8327, 
    263.8152, 263.8441, 263.87, 263.9026, 263.9626, 263.9487, 263.9989, 
    263.4856, 263.5164, 263.5137, 263.546, 263.5698, 263.6215, 263.7043, 
    263.6732, 263.7303, 263.7418, 263.6549, 263.7083, 263.537, 263.5646, 
    263.5482, 263.488, 263.6803, 263.5816, 263.7638, 263.7104, 263.8663, 
    263.7887, 263.941, 264.006, 264.0673, 264.1388, 263.5332, 263.5123, 
    263.5498, 263.6016, 263.6497, 263.7136, 263.7202, 263.7321, 263.7632, 
    263.7893, 263.7359, 263.7958, 263.571, 263.6888, 263.5044, 263.5599, 
    263.5985, 263.5816, 263.6696, 263.6903, 263.7745, 263.731, 263.99, 
    263.8754, 264.1933, 264.1045, 263.505, 263.5332, 263.6312, 263.5845, 
    263.7179, 263.7507, 263.7774, 263.8115, 263.8152, 263.8354, 263.8023, 
    263.8341, 263.7138, 263.7675, 263.62, 263.6559, 263.6394, 263.6213, 
    263.6772, 263.7368, 263.7381, 263.7571, 263.8108, 263.7185, 264.0046, 
    263.8279, 263.5639, 263.6181, 263.6259, 263.6049, 263.7474, 263.6958, 
    263.8349, 263.7973, 263.8589, 263.8283, 263.8238, 263.7845, 263.76, 
    263.6982, 263.6478, 263.6079, 263.6172, 263.661, 263.7404, 263.8155, 
    263.799, 263.8542, 263.7083, 263.7694, 263.7458, 263.8075, 263.6723, 
    263.7873, 263.6429, 263.6556, 263.6948, 263.7736, 263.7911, 263.8097, 
    263.7982, 263.7424, 263.7333, 263.6938, 263.6829, 263.6528, 263.6279, 
    263.6506, 263.6745, 263.7425, 263.8036, 263.8704, 263.8867, 263.9645, 
    263.9011, 264.0056, 263.9166, 264.0707, 263.794, 263.9141, 263.6966, 
    263.72, 263.7624, 263.8596, 263.8072, 263.8686, 263.7329, 263.6625, 
    263.6443, 263.6104, 263.6451, 263.6423, 263.6756, 263.6649, 263.7447, 
    263.7018, 263.8237, 263.8681, 263.9936, 264.0705, 264.1488, 264.1833, 
    264.1939, 264.1983 ;

 FIRE_R =
  263.3521, 263.4231, 263.4093, 263.4666, 263.4348, 263.4724, 263.3665, 
    263.4259, 263.388, 263.3585, 263.5777, 263.4692, 263.6906, 263.6214, 
    263.7954, 263.6798, 263.8187, 263.7921, 263.8722, 263.8493, 263.9516, 
    263.8828, 264.0047, 263.9352, 263.9461, 263.8805, 263.4911, 263.5642, 
    263.4867, 263.4972, 263.4925, 263.4355, 263.4067, 263.3466, 263.3575, 
    263.4017, 263.5018, 263.4679, 263.5536, 263.5516, 263.6469, 263.604, 
    263.7642, 263.7187, 263.8502, 263.8171, 263.8487, 263.8391, 263.8488, 
    263.8003, 263.821, 263.7784, 263.612, 263.6609, 263.515, 263.4273, 
    263.3691, 263.3277, 263.3336, 263.3447, 263.402, 263.4558, 263.4969, 
    263.5243, 263.5514, 263.6331, 263.6764, 263.7734, 263.7559, 263.7855, 
    263.8138, 263.8614, 263.8535, 263.8745, 263.7848, 263.8444, 263.746, 
    263.7729, 263.5585, 263.4771, 263.4423, 263.412, 263.3381, 263.3891, 
    263.369, 263.4169, 263.4473, 263.4323, 263.5251, 263.489, 263.679, 
    263.5971, 263.8105, 263.7595, 263.8228, 263.7905, 263.8458, 263.796, 
    263.8823, 263.901, 263.8882, 263.9375, 263.7933, 263.8487, 263.4318, 
    263.4343, 263.4457, 263.3954, 263.3924, 263.3463, 263.3873, 263.4047, 
    263.449, 263.4752, 263.5001, 263.5548, 263.6159, 263.7014, 263.7628, 
    263.804, 263.7787, 263.801, 263.7761, 263.7644, 263.894, 263.8212, 
    263.9304, 263.9244, 263.875, 263.925, 263.436, 263.4219, 263.3728, 
    263.4112, 263.3413, 263.3804, 263.4029, 263.4897, 263.5088, 263.5265, 
    263.5614, 263.6062, 263.6847, 263.7531, 263.8155, 263.8109, 263.8125, 
    263.8265, 263.792, 263.8321, 263.8389, 263.8213, 263.9236, 263.8943, 
    263.9243, 263.9052, 263.4265, 263.4502, 263.4374, 263.4615, 263.4445, 
    263.5201, 263.5427, 263.6487, 263.6053, 263.6745, 263.6123, 263.6233, 
    263.6767, 263.6157, 263.7493, 263.6587, 263.827, 263.7365, 263.8327, 
    263.8152, 263.8441, 263.87, 263.9026, 263.9626, 263.9487, 263.9989, 
    263.4856, 263.5164, 263.5137, 263.546, 263.5698, 263.6215, 263.7043, 
    263.6732, 263.7303, 263.7418, 263.6549, 263.7083, 263.537, 263.5646, 
    263.5482, 263.488, 263.6803, 263.5816, 263.7638, 263.7104, 263.8663, 
    263.7887, 263.941, 264.006, 264.0673, 264.1388, 263.5332, 263.5123, 
    263.5498, 263.6016, 263.6497, 263.7136, 263.7202, 263.7321, 263.7632, 
    263.7893, 263.7359, 263.7958, 263.571, 263.6888, 263.5044, 263.5599, 
    263.5985, 263.5816, 263.6696, 263.6903, 263.7745, 263.731, 263.99, 
    263.8754, 264.1933, 264.1045, 263.505, 263.5332, 263.6312, 263.5845, 
    263.7179, 263.7507, 263.7774, 263.8115, 263.8152, 263.8354, 263.8023, 
    263.8341, 263.7138, 263.7675, 263.62, 263.6559, 263.6394, 263.6213, 
    263.6772, 263.7368, 263.7381, 263.7571, 263.8108, 263.7185, 264.0046, 
    263.8279, 263.5639, 263.6181, 263.6259, 263.6049, 263.7474, 263.6958, 
    263.8349, 263.7973, 263.8589, 263.8283, 263.8238, 263.7845, 263.76, 
    263.6982, 263.6478, 263.6079, 263.6172, 263.661, 263.7404, 263.8155, 
    263.799, 263.8542, 263.7083, 263.7694, 263.7458, 263.8075, 263.6723, 
    263.7873, 263.6429, 263.6556, 263.6948, 263.7736, 263.7911, 263.8097, 
    263.7982, 263.7424, 263.7333, 263.6938, 263.6829, 263.6528, 263.6279, 
    263.6506, 263.6745, 263.7425, 263.8036, 263.8704, 263.8867, 263.9645, 
    263.9011, 264.0056, 263.9166, 264.0707, 263.794, 263.9141, 263.6966, 
    263.72, 263.7624, 263.8596, 263.8072, 263.8686, 263.7329, 263.6625, 
    263.6443, 263.6104, 263.6451, 263.6423, 263.6756, 263.6649, 263.7447, 
    263.7018, 263.8237, 263.8681, 263.9936, 264.0705, 264.1488, 264.1833, 
    264.1939, 264.1983 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSA_R =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347 ;

 FSDSND =
  0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532 ;

 FSDSNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSDSNI =
  0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819 ;

 FSDSVD =
  0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128 ;

 FSDSVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSDSVI =
  0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223 ;

 FSDSVILN =
  0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376 ;

 FSH =
  354.1815, 355.0652, 354.8935, 355.6059, 355.2109, 355.6772, 354.3609, 
    355.1, 354.6283, 354.2614, 356.9875, 355.6378, 358.3912, 357.5304, 
    359.6931, 358.257, 359.9827, 359.6522, 360.6481, 360.3628, 361.6351, 
    360.7797, 362.2952, 361.4311, 361.5661, 360.7514, 355.9099, 356.8193, 
    355.8559, 355.9856, 355.9275, 355.2189, 354.8615, 354.1143, 354.25, 
    354.799, 356.044, 355.6217, 356.6868, 356.6628, 357.8479, 357.3136, 
    359.3053, 358.7394, 360.3748, 359.9635, 360.3553, 360.2366, 360.3569, 
    359.7538, 360.0121, 359.4815, 357.4135, 358.0213, 356.2082, 355.1169, 
    354.3932, 353.8792, 353.9519, 354.0903, 354.8022, 355.4719, 355.982, 
    356.3232, 356.6593, 357.6754, 358.2142, 359.4194, 359.2024, 359.5704, 
    359.9226, 360.5132, 360.416, 360.6761, 359.561, 360.302, 359.0787, 
    359.4132, 356.7489, 355.7357, 355.3035, 354.9265, 354.0077, 354.6421, 
    354.392, 354.9874, 355.3654, 355.1785, 356.3325, 355.8838, 358.2461, 
    357.2288, 359.8815, 359.247, 360.0337, 359.6324, 360.3198, 359.7011, 
    360.773, 361.0062, 360.8468, 361.4595, 359.6668, 360.3552, 355.1732, 
    355.2036, 355.3458, 354.7209, 354.6827, 354.1105, 354.6198, 354.8365, 
    355.3874, 355.7129, 356.0224, 356.7029, 357.4625, 358.5248, 359.2881, 
    359.7996, 359.4861, 359.7628, 359.4534, 359.3084, 360.9187, 360.0145, 
    361.3714, 361.2964, 360.6822, 361.3048, 355.2251, 355.0497, 354.4401, 
    354.9171, 354.0482, 354.5344, 354.8138, 355.8928, 356.1302, 356.3499, 
    356.784, 357.3409, 358.3175, 359.1673, 359.9431, 359.8864, 359.9063, 
    360.0794, 359.6504, 360.1499, 360.2336, 360.0146, 361.2863, 360.9231, 
    361.2948, 361.0583, 355.1067, 355.4019, 355.2424, 355.5423, 355.3309, 
    356.2705, 356.5522, 357.8704, 357.3299, 358.1906, 357.4174, 357.5544, 
    358.2179, 357.4594, 359.1201, 357.9936, 360.0862, 358.9608, 360.1566, 
    359.9398, 360.299, 360.6205, 361.0251, 361.7711, 361.5985, 362.2226, 
    355.8422, 356.2249, 356.1915, 356.5922, 356.8884, 357.5309, 358.5606, 
    358.1735, 358.8845, 359.027, 357.9471, 358.6099, 356.4812, 356.8249, 
    356.6205, 355.8722, 358.2622, 357.0356, 359.3007, 358.6365, 360.5746, 
    359.6105, 361.5034, 362.3112, 363.073, 363.961, 356.4341, 356.174, 
    356.64, 357.2839, 357.8822, 358.6769, 358.7584, 358.9072, 359.2929, 
    359.617, 358.9539, 359.6983, 356.9039, 358.3688, 356.0754, 356.7657, 
    357.2461, 357.0357, 358.1293, 358.3869, 359.4334, 358.8927, 362.1116, 
    360.6879, 364.638, 363.5345, 356.0831, 356.4333, 357.6516, 357.0721, 
    358.7302, 359.138, 359.4698, 359.8934, 359.9394, 360.1904, 359.7791, 
    360.1743, 358.6786, 359.3471, 357.5128, 357.9592, 357.7539, 357.5286, 
    358.224, 358.9643, 358.9806, 359.2178, 359.8853, 358.7369, 362.2943, 
    360.0969, 356.8152, 357.489, 357.5859, 357.3248, 359.0971, 358.455, 
    360.1843, 359.7171, 360.4827, 360.1023, 360.0463, 359.5577, 359.2533, 
    358.4843, 357.8586, 357.3627, 357.4781, 358.0228, 359.0097, 359.9433, 
    359.7387, 360.4245, 358.61, 359.3707, 359.0765, 359.8436, 358.1631, 
    359.5926, 357.7974, 357.955, 358.4422, 359.4219, 359.6394, 359.8707, 
    359.7281, 359.0348, 358.9214, 358.4305, 358.2947, 357.9207, 357.6108, 
    357.8938, 358.1909, 359.0353, 359.7958, 360.6249, 360.828, 361.795, 
    361.0071, 362.3064, 361.2007, 363.1151, 359.6762, 361.1693, 358.4646, 
    358.7562, 359.283, 360.4922, 359.84, 360.6029, 358.9171, 358.0414, 
    357.8154, 357.3928, 357.8251, 357.7899, 358.2036, 358.0707, 359.0634, 
    358.5302, 360.0447, 360.5971, 362.157, 363.1125, 364.0856, 364.5148, 
    364.6454, 364.7 ;

 FSH_G =
  360.841, 361.7252, 361.5534, 362.2663, 361.8711, 362.3376, 361.0205, 
    361.7601, 361.2881, 360.9209, 363.6487, 362.2981, 365.0533, 364.192, 
    366.356, 364.919, 366.6458, 366.3151, 367.3116, 367.0262, 368.2992, 
    367.4433, 368.9597, 368.0951, 368.2302, 367.415, 362.5705, 363.4804, 
    362.5164, 362.6462, 362.5881, 361.879, 361.5213, 360.7737, 360.9095, 
    361.4588, 362.7046, 362.2821, 363.3479, 363.3238, 364.5096, 363.975, 
    365.968, 365.4018, 367.0381, 366.6266, 367.0187, 366.8998, 367.0202, 
    366.4167, 366.6752, 366.1443, 364.075, 364.6831, 362.8689, 361.7769, 
    361.0528, 360.5385, 360.6112, 360.7497, 361.4621, 362.1321, 362.6426, 
    362.9839, 363.3203, 364.337, 364.8762, 366.0822, 365.865, 366.2332, 
    366.5857, 367.1766, 367.0794, 367.3396, 366.2239, 366.9653, 365.7412, 
    366.076, 363.41, 362.3962, 361.9637, 361.5864, 360.6671, 361.3018, 
    361.0516, 361.6473, 362.0256, 361.8386, 362.9933, 362.5443, 364.9081, 
    363.8901, 366.5446, 365.9096, 366.6968, 366.2952, 366.9831, 366.364, 
    367.4366, 367.6699, 367.5104, 368.1235, 366.3297, 367.0185, 361.8333, 
    361.8638, 362.006, 361.3807, 361.3425, 360.7699, 361.2796, 361.4965, 
    362.0477, 362.3734, 362.6831, 363.364, 364.124, 365.187, 365.9508, 
    366.4626, 366.1489, 366.4258, 366.1161, 365.9711, 367.5824, 366.6776, 
    368.0353, 367.9603, 367.3457, 367.9688, 361.8852, 361.7097, 361.0997, 
    361.5771, 360.7076, 361.1941, 361.4737, 362.5533, 362.791, 363.0107, 
    363.4451, 364.0023, 364.9796, 365.8299, 366.6062, 366.5494, 366.5694, 
    366.7426, 366.3133, 366.8131, 366.8968, 366.6777, 367.9502, 367.5868, 
    367.9587, 367.7221, 361.7668, 362.0622, 361.9026, 362.2026, 361.9911, 
    362.9312, 363.2131, 364.5321, 363.9913, 364.8525, 364.0789, 364.2159, 
    364.8798, 364.1208, 365.7827, 364.6554, 366.7493, 365.6232, 366.8198, 
    366.6029, 366.9623, 367.2839, 367.6889, 368.4354, 368.2626, 368.8871, 
    362.5027, 362.8856, 362.8522, 363.2532, 363.5496, 364.1924, 365.2228, 
    364.8355, 365.5469, 365.6895, 364.6089, 365.2721, 363.1421, 363.486, 
    363.2815, 362.5327, 364.9243, 363.6969, 365.9633, 365.2987, 367.238, 
    366.2734, 368.1674, 368.9758, 369.738, 370.6266, 363.0949, 362.8347, 
    363.301, 363.9453, 364.5439, 365.3392, 365.4207, 365.5696, 365.9556, 
    366.2799, 365.6163, 366.3612, 363.5651, 365.0309, 362.7361, 363.4268, 
    363.9074, 363.6969, 364.7913, 365.049, 366.0962, 365.5551, 368.776, 
    367.3514, 371.304, 370.1998, 362.7437, 363.0942, 364.3133, 363.7334, 
    365.3925, 365.8006, 366.1326, 366.5565, 366.6024, 366.8536, 366.442, 
    366.8375, 365.3409, 366.0098, 364.1743, 364.621, 364.4156, 364.1902, 
    364.886, 365.6267, 365.6431, 365.8804, 366.5482, 365.3992, 368.9588, 
    366.7601, 363.4763, 364.1505, 364.2475, 363.9862, 365.7596, 365.1171, 
    366.8475, 366.3801, 367.1461, 366.7654, 366.7094, 366.2205, 365.9159, 
    365.1465, 364.5204, 364.0242, 364.1396, 364.6847, 365.6721, 366.6064, 
    366.4017, 367.0879, 365.2722, 366.0334, 365.739, 366.5066, 364.8251, 
    366.2554, 364.4592, 364.6168, 365.1043, 366.0846, 366.3023, 366.5337, 
    366.391, 365.6973, 365.5839, 365.0926, 364.9567, 364.5825, 364.2724, 
    364.5556, 364.8529, 365.6978, 366.4588, 367.2884, 367.4916, 368.4592, 
    367.6709, 368.9709, 367.8645, 369.7801, 366.3391, 367.8331, 365.1267, 
    365.4185, 365.9457, 367.1555, 366.503, 367.2664, 365.5795, 364.7032, 
    364.4772, 364.0542, 364.4868, 364.4517, 364.8656, 364.7326, 365.7259, 
    365.1924, 366.7079, 367.2605, 368.8214, 369.7775, 370.7512, 371.1807, 
    371.3115, 371.3661 ;

 FSH_NODYNLNDUSE =
  354.1815, 355.0652, 354.8935, 355.6059, 355.2109, 355.6772, 354.3609, 
    355.1, 354.6283, 354.2614, 356.9875, 355.6378, 358.3912, 357.5304, 
    359.6931, 358.257, 359.9827, 359.6522, 360.6481, 360.3628, 361.6351, 
    360.7797, 362.2952, 361.4311, 361.5661, 360.7514, 355.9099, 356.8193, 
    355.8559, 355.9856, 355.9275, 355.2189, 354.8615, 354.1143, 354.25, 
    354.799, 356.044, 355.6217, 356.6868, 356.6628, 357.8479, 357.3136, 
    359.3053, 358.7394, 360.3748, 359.9635, 360.3553, 360.2366, 360.3569, 
    359.7538, 360.0121, 359.4815, 357.4135, 358.0213, 356.2082, 355.1169, 
    354.3932, 353.8792, 353.9519, 354.0903, 354.8022, 355.4719, 355.982, 
    356.3232, 356.6593, 357.6754, 358.2142, 359.4194, 359.2024, 359.5704, 
    359.9226, 360.5132, 360.416, 360.6761, 359.561, 360.302, 359.0787, 
    359.4132, 356.7489, 355.7357, 355.3035, 354.9265, 354.0077, 354.6421, 
    354.392, 354.9874, 355.3654, 355.1785, 356.3325, 355.8838, 358.2461, 
    357.2288, 359.8815, 359.247, 360.0337, 359.6324, 360.3198, 359.7011, 
    360.773, 361.0062, 360.8468, 361.4595, 359.6668, 360.3552, 355.1732, 
    355.2036, 355.3458, 354.7209, 354.6827, 354.1105, 354.6198, 354.8365, 
    355.3874, 355.7129, 356.0224, 356.7029, 357.4625, 358.5248, 359.2881, 
    359.7996, 359.4861, 359.7628, 359.4534, 359.3084, 360.9187, 360.0145, 
    361.3714, 361.2964, 360.6822, 361.3048, 355.2251, 355.0497, 354.4401, 
    354.9171, 354.0482, 354.5344, 354.8138, 355.8928, 356.1302, 356.3499, 
    356.784, 357.3409, 358.3175, 359.1673, 359.9431, 359.8864, 359.9063, 
    360.0794, 359.6504, 360.1499, 360.2336, 360.0146, 361.2863, 360.9231, 
    361.2948, 361.0583, 355.1067, 355.4019, 355.2424, 355.5423, 355.3309, 
    356.2705, 356.5522, 357.8704, 357.3299, 358.1906, 357.4174, 357.5544, 
    358.2179, 357.4594, 359.1201, 357.9936, 360.0862, 358.9608, 360.1566, 
    359.9398, 360.299, 360.6205, 361.0251, 361.7711, 361.5985, 362.2226, 
    355.8422, 356.2249, 356.1915, 356.5922, 356.8884, 357.5309, 358.5606, 
    358.1735, 358.8845, 359.027, 357.9471, 358.6099, 356.4812, 356.8249, 
    356.6205, 355.8722, 358.2622, 357.0356, 359.3007, 358.6365, 360.5746, 
    359.6105, 361.5034, 362.3112, 363.073, 363.961, 356.4341, 356.174, 
    356.64, 357.2839, 357.8822, 358.6769, 358.7584, 358.9072, 359.2929, 
    359.617, 358.9539, 359.6983, 356.9039, 358.3688, 356.0754, 356.7657, 
    357.2461, 357.0357, 358.1293, 358.3869, 359.4334, 358.8927, 362.1116, 
    360.6879, 364.638, 363.5345, 356.0831, 356.4333, 357.6516, 357.0721, 
    358.7302, 359.138, 359.4698, 359.8934, 359.9394, 360.1904, 359.7791, 
    360.1743, 358.6786, 359.3471, 357.5128, 357.9592, 357.7539, 357.5286, 
    358.224, 358.9643, 358.9806, 359.2178, 359.8853, 358.7369, 362.2943, 
    360.0969, 356.8152, 357.489, 357.5859, 357.3248, 359.0971, 358.455, 
    360.1843, 359.7171, 360.4827, 360.1023, 360.0463, 359.5577, 359.2533, 
    358.4843, 357.8586, 357.3627, 357.4781, 358.0228, 359.0097, 359.9433, 
    359.7387, 360.4245, 358.61, 359.3707, 359.0765, 359.8436, 358.1631, 
    359.5926, 357.7974, 357.955, 358.4422, 359.4219, 359.6394, 359.8707, 
    359.7281, 359.0348, 358.9214, 358.4305, 358.2947, 357.9207, 357.6108, 
    357.8938, 358.1909, 359.0353, 359.7958, 360.6249, 360.828, 361.795, 
    361.0071, 362.3064, 361.2007, 363.1151, 359.6762, 361.1693, 358.4646, 
    358.7562, 359.283, 360.4922, 359.84, 360.6029, 358.9171, 358.0414, 
    357.8154, 357.3928, 357.8251, 357.7899, 358.2036, 358.0707, 359.0634, 
    358.5302, 360.0447, 360.5971, 362.157, 363.1125, 364.0856, 364.5148, 
    364.6454, 364.7 ;

 FSH_R =
  354.1815, 355.0652, 354.8935, 355.6059, 355.2109, 355.6772, 354.3609, 
    355.1, 354.6283, 354.2614, 356.9875, 355.6378, 358.3912, 357.5304, 
    359.6931, 358.257, 359.9827, 359.6522, 360.6481, 360.3628, 361.6351, 
    360.7797, 362.2952, 361.4311, 361.5661, 360.7514, 355.9099, 356.8193, 
    355.8559, 355.9856, 355.9275, 355.2189, 354.8615, 354.1143, 354.25, 
    354.799, 356.044, 355.6217, 356.6868, 356.6628, 357.8479, 357.3136, 
    359.3053, 358.7394, 360.3748, 359.9635, 360.3553, 360.2366, 360.3569, 
    359.7538, 360.0121, 359.4815, 357.4135, 358.0213, 356.2082, 355.1169, 
    354.3932, 353.8792, 353.9519, 354.0903, 354.8022, 355.4719, 355.982, 
    356.3232, 356.6593, 357.6754, 358.2142, 359.4194, 359.2024, 359.5704, 
    359.9226, 360.5132, 360.416, 360.6761, 359.561, 360.302, 359.0787, 
    359.4132, 356.7489, 355.7357, 355.3035, 354.9265, 354.0077, 354.6421, 
    354.392, 354.9874, 355.3654, 355.1785, 356.3325, 355.8838, 358.2461, 
    357.2288, 359.8815, 359.247, 360.0337, 359.6324, 360.3198, 359.7011, 
    360.773, 361.0062, 360.8468, 361.4595, 359.6668, 360.3552, 355.1732, 
    355.2036, 355.3458, 354.7209, 354.6827, 354.1105, 354.6198, 354.8365, 
    355.3874, 355.7129, 356.0224, 356.7029, 357.4625, 358.5248, 359.2881, 
    359.7996, 359.4861, 359.7628, 359.4534, 359.3084, 360.9187, 360.0145, 
    361.3714, 361.2964, 360.6822, 361.3048, 355.2251, 355.0497, 354.4401, 
    354.9171, 354.0482, 354.5344, 354.8138, 355.8928, 356.1302, 356.3499, 
    356.784, 357.3409, 358.3175, 359.1673, 359.9431, 359.8864, 359.9063, 
    360.0794, 359.6504, 360.1499, 360.2336, 360.0146, 361.2863, 360.9231, 
    361.2948, 361.0583, 355.1067, 355.4019, 355.2424, 355.5423, 355.3309, 
    356.2705, 356.5522, 357.8704, 357.3299, 358.1906, 357.4174, 357.5544, 
    358.2179, 357.4594, 359.1201, 357.9936, 360.0862, 358.9608, 360.1566, 
    359.9398, 360.299, 360.6205, 361.0251, 361.7711, 361.5985, 362.2226, 
    355.8422, 356.2249, 356.1915, 356.5922, 356.8884, 357.5309, 358.5606, 
    358.1735, 358.8845, 359.027, 357.9471, 358.6099, 356.4812, 356.8249, 
    356.6205, 355.8722, 358.2622, 357.0356, 359.3007, 358.6365, 360.5746, 
    359.6105, 361.5034, 362.3112, 363.073, 363.961, 356.4341, 356.174, 
    356.64, 357.2839, 357.8822, 358.6769, 358.7584, 358.9072, 359.2929, 
    359.617, 358.9539, 359.6983, 356.9039, 358.3688, 356.0754, 356.7657, 
    357.2461, 357.0357, 358.1293, 358.3869, 359.4334, 358.8927, 362.1116, 
    360.6879, 364.638, 363.5345, 356.0831, 356.4333, 357.6516, 357.0721, 
    358.7302, 359.138, 359.4698, 359.8934, 359.9394, 360.1904, 359.7791, 
    360.1743, 358.6786, 359.3471, 357.5128, 357.9592, 357.7539, 357.5286, 
    358.224, 358.9643, 358.9806, 359.2178, 359.8853, 358.7369, 362.2943, 
    360.0969, 356.8152, 357.489, 357.5859, 357.3248, 359.0971, 358.455, 
    360.1843, 359.7171, 360.4827, 360.1023, 360.0463, 359.5577, 359.2533, 
    358.4843, 357.8586, 357.3627, 357.4781, 358.0228, 359.0097, 359.9433, 
    359.7387, 360.4245, 358.61, 359.3707, 359.0765, 359.8436, 358.1631, 
    359.5926, 357.7974, 357.955, 358.4422, 359.4219, 359.6394, 359.8707, 
    359.7281, 359.0348, 358.9214, 358.4305, 358.2947, 357.9207, 357.6108, 
    357.8938, 358.1909, 359.0353, 359.7958, 360.6249, 360.828, 361.795, 
    361.0071, 362.3064, 361.2007, 363.1151, 359.6762, 361.1693, 358.4646, 
    358.7562, 359.283, 360.4922, 359.84, 360.6029, 358.9171, 358.0414, 
    357.8154, 357.3928, 357.8251, 357.7899, 358.2036, 358.0707, 359.0634, 
    358.5302, 360.0447, 360.5971, 362.157, 363.1125, 364.0856, 364.5148, 
    364.6454, 364.7 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -6.659477, -6.660025, -6.659921, -6.660357, -6.66012, -6.660402, -6.659593, 
    -6.660043, -6.659759, -6.659534, -6.661191, -6.660378, -6.662084, 
    -6.661556, -6.662898, -6.661995, -6.663082, -6.662882, -6.663509, 
    -6.663331, -6.664111, -6.663592, -6.664534, -6.663993, -6.664073, 
    -6.663573, -6.660552, -6.661087, -6.660518, -6.660595, -6.660563, 
    -6.66012, -6.659891, -6.659443, -6.659526, -6.659859, -6.660629, 
    -6.660375, -6.661038, -6.661023, -6.661755, -6.661425, -6.662665, 
    -6.662314, -6.663338, -6.663079, -6.663324, -6.663251, -6.663325, 
    -6.662945, -6.663107, -6.662777, -6.661484, -6.66186, -6.660735, 
    -6.660043, -6.659611, -6.659297, -6.659341, -6.659423, -6.659861, 
    -6.660282, -6.6606, -6.660811, -6.661021, -6.661628, -6.661973, 
    -6.662731, -6.662603, -6.662827, -6.663054, -6.663422, -6.663363, 
    -6.663523, -6.662827, -6.663286, -6.662529, -6.662734, -6.661041, 
    -6.660445, -6.660161, -6.65994, -6.659374, -6.659763, -6.659609, 
    -6.659983, -6.660216, -6.660102, -6.660817, -6.660538, -6.661994, 
    -6.661366, -6.663027, -6.66263, -6.663124, -6.662873, -6.663299, 
    -6.662916, -6.663585, -6.663727, -6.66363, -6.664017, -6.662894, 
    -6.663321, -6.660097, -6.660116, -6.660205, -6.659811, -6.659789, 
    -6.659439, -6.659754, -6.659884, -6.660232, -6.660431, -6.660622, 
    -6.661044, -6.66151, -6.662173, -6.662655, -6.662978, -6.662783, 
    -6.662955, -6.662761, -6.662672, -6.663671, -6.663106, -6.663961, 
    -6.663915, -6.663525, -6.66392, -6.660129, -6.660023, -6.659641, 
    -6.65994, -6.659401, -6.659698, -6.659866, -6.660535, -6.660691, 
    -6.660825, -6.661097, -6.661441, -6.662045, -6.662576, -6.663068, 
    -6.663033, -6.663045, -6.663151, -6.662883, -6.663195, -6.663244, 
    -6.663111, -6.663909, -6.663681, -6.663914, -6.663767, -6.660058, 
    -6.660239, -6.660141, -6.660324, -6.660192, -6.660768, -6.66094, 
    -6.66176, -6.661432, -6.661964, -6.661489, -6.661571, -6.661965, 
    -6.661517, -6.66254, -6.661832, -6.663155, -6.662432, -6.663199, 
    -6.663066, -6.663291, -6.663489, -6.663744, -6.664207, -6.664101, 
    -6.664494, -6.660512, -6.660744, -6.66073, -6.660977, -6.661159, 
    -6.661561, -6.662199, -6.661962, -6.662406, -6.662493, -6.661822, 
    -6.662227, -6.660904, -6.66111, -6.660993, -6.660526, -6.662006, 
    -6.661242, -6.662662, -6.662248, -6.66346, -6.662849, -6.664041, 
    -6.664534, -6.665031, -6.665576, -6.660878, -6.660719, -6.661009, 
    -6.661397, -6.661777, -6.662272, -6.662327, -6.662417, -6.662662, 
    -6.662863, -6.662439, -6.662915, -6.661144, -6.662076, -6.660653, 
    -6.661072, -6.661377, -6.66125, -6.661936, -6.662096, -6.662742, 
    -6.662411, -6.664406, -6.663521, -6.666014, -6.66531, -6.660663, 
    -6.66088, -6.661629, -6.661274, -6.662309, -6.662561, -6.662773, 
    -6.663032, -6.663064, -6.663219, -6.662965, -6.663212, -6.662273, 
    -6.662693, -6.661552, -6.661825, -6.661702, -6.661561, -6.661994, 
    -6.662445, -6.662465, -6.662608, -6.66299, -6.662313, -6.6645, -6.663128, 
    -6.661117, -6.661522, -6.661593, -6.661434, -6.662536, -6.662135, 
    -6.663217, -6.662926, -6.663405, -6.663166, -6.66313, -6.662827, 
    -6.662634, -6.662151, -6.661761, -6.661458, -6.66153, -6.661863, 
    -6.662475, -6.663063, -6.662932, -6.663369, -6.662233, -6.662703, 
    -6.662518, -6.663003, -6.661952, -6.662813, -6.661729, -6.661826, 
    -6.662127, -6.662727, -6.662878, -6.663017, -6.662933, -6.662492, 
    -6.662425, -6.662122, -6.662033, -6.661806, -6.661613, -6.661787, 
    -6.661967, -6.662497, -6.66297, -6.66349, -6.663622, -6.664203, 
    -6.663714, -6.664505, -6.663809, -6.665027, -6.66288, -6.663812, 
    -6.662144, -6.662326, -6.662643, -6.663396, -6.663002, -6.663469, 
    -6.662423, -6.661869, -6.661739, -6.661475, -6.661746, -6.661724, 
    -6.661982, -6.6619, -6.662515, -6.662185, -6.663126, -6.663468, 
    -6.664448, -6.665044, -6.665669, -6.66594, -6.666024, -6.666058 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179 ;

 FSRND =
  0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234 ;

 FSRNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSRNI =
  0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666 ;

 FSRVD =
  0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223 ;

 FSRVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSRVI =
  0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.904545e-44, 0, 3.640714e-41, 
    2.382207e-44, 1.485699e-40, 2.970192e-41, 3.462017e-39, 9.090784e-40, 
    3.043702e-37, 6.372947e-39, 5.297037e-36, 1.228662e-37, 2.240759e-37, 
    5.592868e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 
    5.327737e-42, 3.012792e-43, 9.616453e-40, 1.350768e-40, 8.778827e-40, 
    4.997395e-40, 8.843286e-40, 4.883105e-41, 1.708729e-40, 1.279946e-41, 0, 
    7.006492e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    1.961818e-44, 9.427936e-42, 3.179546e-42, 1.989283e-41, 1.108483e-40, 
    1.845646e-39, 1.168838e-39, 3.948533e-39, 1.895536e-41, 6.828597e-40, 
    1.702578e-42, 9.121052e-42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.242078e-44, 0, 9.087421e-41, 3.976885e-42, 1.893603e-40, 2.691614e-41, 
    7.425691e-40, 3.771455e-41, 6.183549e-39, 1.806158e-38, 8.695494e-39, 
    1.391768e-37, 3.187954e-41, 8.78027e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9.949219e-44, 4.887729e-42, 6.099011e-41, 1.308112e-41, 
    5.099465e-41, 1.112771e-41, 5.404808e-42, 1.210799e-38, 1.728852e-40, 
    9.393621e-38, 6.709526e-38, 4.063952e-39, 6.969254e-38, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3.363116e-44, 2.668072e-42, 1.22367e-40, 9.295093e-41, 
    1.024097e-40, 2.360095e-40, 2.942166e-41, 3.306658e-40, 4.932346e-40, 
    1.727591e-40, 6.41323e-38, 1.233066e-38, 6.661603e-38, 2.286338e-38, 0, 
    0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 1.681558e-44, 0, 0, 1.961818e-44, 0, 
    2.107553e-42, 5.605194e-45, 2.437545e-40, 9.416726e-43, 3.41488e-40, 
    1.20401e-40, 6.718792e-40, 3.047178e-39, 1.966447e-38, 5.518767e-37, 
    2.580681e-37, 3.881303e-36, 0, 0, 0, 0, 0, 0, 1.191104e-43, 1.541428e-44, 
    6.347882e-43, 1.311615e-42, 4.203895e-45, 1.541428e-43, 0, 0, 0, 0, 
    2.522337e-44, 0, 5.205824e-42, 1.765636e-43, 2.460338e-39, 2.425227e-41, 
    1.693173e-37, 5.68547e-36, 1.346246e-34, 4.604947e-33, 0, 0, 0, 0, 
    2.802597e-45, 2.186026e-43, 3.321077e-43, 7.132609e-43, 5.002636e-42, 
    2.496693e-41, 9.066401e-43, 3.719607e-41, 0, 4.344025e-44, 0, 0, 0, 0, 
    1.261169e-44, 4.764415e-44, 1.009916e-41, 6.614129e-43, 2.424143e-36, 
    4.18154e-39, 6.026268e-32, 8.63849e-34, 0, 0, 1.401298e-45, 0, 
    2.872662e-43, 2.299531e-42, 1.206938e-41, 9.634768e-41, 1.20202e-40, 
    4.013333e-40, 5.518173e-41, 3.713385e-40, 2.200039e-43, 6.562281e-42, 0, 
    5.605194e-45, 1.401298e-45, 0, 2.101948e-44, 9.556856e-43, 1.03556e-42, 
    3.440188e-42, 9.359973e-41, 2.970753e-43, 5.321813e-36, 2.591547e-40, 0, 
    0, 0, 0, 1.870733e-42, 6.866362e-44, 3.897558e-40, 4.0789e-41, 
    1.598796e-39, 2.632255e-40, 2.012363e-40, 1.863867e-41, 4.105805e-42, 
    7.987401e-44, 2.802597e-45, 0, 0, 7.006492e-45, 1.203715e-42, 
    1.226613e-40, 4.54329e-41, 1.216202e-39, 1.541428e-43, 7.390448e-42, 
    1.688565e-42, 7.559725e-41, 1.541428e-44, 2.236612e-41, 1.401298e-45, 
    4.203895e-45, 6.445973e-44, 9.556856e-42, 2.787043e-41, 8.629336e-41, 
    4.303107e-41, 1.366266e-42, 7.665103e-43, 6.025583e-44, 2.942727e-44, 
    4.203895e-45, 1.401298e-45, 4.203895e-45, 1.681558e-44, 1.367667e-42, 
    5.998398e-41, 3.113122e-39, 7.966207e-39, 6.155813e-37, 1.82089e-38, 
    5.606511e-36, 4.415561e-38, 1.609795e-34, 3.358352e-41, 3.807932e-38, 
    7.286752e-44, 3.279038e-43, 4.778428e-42, 1.678356e-39, 7.428563e-41, 
    2.815552e-39, 7.496947e-43, 8.407791e-45, 2.802597e-45, 0, 2.802597e-45, 
    1.401298e-45, 1.821688e-44, 8.407791e-45, 1.576461e-42, 1.022948e-43, 
    1.99912e-40, 2.737107e-39, 2.934797e-36, 1.585659e-34, 7.423095e-33, 
    3.795473e-32, 6.187504e-32, 7.582037e-32 ;

 F_DENIT_vr =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.007714e-43, 4.203895e-45, 
    2.945543e-40, 1.975831e-43, 1.20202e-39, 2.403045e-40, 2.800977e-38, 
    7.35498e-39, 2.462535e-36, 5.156091e-38, 4.285616e-35, 9.9406e-37, 
    1.812906e-36, 4.524961e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.242078e-44, 1.401298e-45, 4.310674e-41, 2.438259e-42, 7.78028e-39, 
    1.092854e-39, 7.102588e-39, 4.043189e-39, 7.154737e-39, 3.950737e-40, 
    1.382462e-39, 1.035532e-40, 1.401298e-45, 5.605194e-44, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8.407791e-45, 1.569454e-43, 7.627268e-41, 2.571943e-41, 
    1.609475e-40, 8.96831e-40, 1.493236e-38, 9.456588e-39, 3.194596e-38, 
    1.533637e-40, 5.524734e-39, 1.377056e-41, 7.379798e-41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.863727e-43, 1.401298e-45, 7.352235e-40, 3.218082e-41, 
    1.532035e-39, 2.17766e-40, 6.007822e-39, 3.051285e-40, 5.002857e-38, 
    1.461288e-37, 7.035169e-38, 1.126023e-36, 2.57923e-40, 7.103752e-39, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.802597e-45, 8.043453e-43, 
    3.954464e-41, 4.934504e-40, 1.058289e-40, 4.125801e-40, 9.003203e-41, 
    4.372331e-41, 9.796078e-38, 1.398748e-39, 7.599994e-37, 5.428403e-37, 
    3.287978e-38, 5.638538e-37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.401298e-45, 2.718519e-43, 2.158981e-41, 9.900258e-40, 7.52025e-40, 
    8.285556e-40, 1.90946e-39, 2.380414e-40, 2.675279e-39, 3.990559e-39, 
    1.397721e-39, 5.188682e-37, 9.976233e-38, 5.389631e-37, 1.849783e-37, 0, 
    0, 0, 0, 0, 0, 0, 2.522337e-44, 1.401298e-45, 1.387285e-43, 2.802597e-45, 
    4.203895e-45, 1.611493e-43, 2.802597e-45, 1.70538e-41, 4.904545e-44, 
    1.972117e-39, 7.623064e-42, 2.762845e-39, 9.74114e-40, 5.435895e-39, 
    2.465347e-38, 1.590971e-37, 4.465009e-36, 2.087923e-36, 3.140203e-35, 0, 
    0, 0, 0, 0, 4.203895e-45, 9.668959e-43, 1.261169e-43, 5.130154e-42, 
    1.061203e-41, 3.783506e-44, 1.25136e-42, 0, 0, 0, 0, 2.031883e-43, 0, 
    4.212163e-41, 1.433528e-42, 1.990559e-38, 1.96214e-40, 1.369877e-36, 
    4.599881e-35, 1.089193e-33, 3.725674e-32, 0, 0, 0, 1.401298e-45, 
    2.662467e-44, 1.768439e-42, 2.68769e-42, 5.766343e-42, 4.04695e-41, 
    2.020014e-40, 7.334396e-42, 3.009373e-40, 0, 3.559298e-43, 0, 0, 
    1.401298e-45, 0, 9.949219e-44, 3.89561e-43, 8.170691e-41, 5.350158e-42, 
    1.961275e-35, 3.383113e-38, 4.875606e-31, 6.989049e-33, 0, 0, 
    7.006492e-45, 0, 2.324754e-42, 1.860784e-41, 9.764808e-41, 7.795143e-40, 
    9.724997e-40, 3.247019e-39, 4.464509e-40, 3.004352e-39, 1.783853e-42, 
    5.308959e-41, 4.203895e-45, 4.063766e-44, 1.401298e-44, 4.203895e-45, 
    1.653532e-43, 7.735168e-42, 8.378364e-42, 2.783399e-41, 7.572729e-40, 
    2.406029e-42, 4.305662e-35, 2.09671e-39, 0, 2.802597e-45, 5.605194e-45, 
    1.401298e-45, 1.513683e-41, 5.577168e-43, 3.15336e-39, 3.3001e-40, 
    1.293521e-38, 2.129647e-39, 1.62812e-39, 1.508007e-40, 3.321638e-41, 
    6.502025e-43, 2.382207e-44, 1.401298e-45, 2.802597e-45, 5.745324e-44, 
    9.737623e-42, 9.924024e-40, 3.675802e-40, 9.839797e-39, 1.248557e-42, 
    5.97906e-41, 1.365705e-41, 6.116303e-40, 1.191104e-43, 1.809553e-40, 
    1.681558e-44, 3.923636e-44, 5.21283e-43, 7.732365e-41, 2.254941e-40, 
    6.981605e-40, 3.481456e-40, 1.105624e-41, 6.20495e-42, 4.904545e-43, 
    2.410233e-43, 3.222986e-44, 5.605194e-45, 2.802597e-44, 1.387285e-43, 
    1.107026e-41, 4.853033e-40, 2.5187e-38, 6.445132e-38, 4.980416e-36, 
    1.473207e-37, 4.535999e-35, 3.57245e-37, 1.302419e-33, 2.717132e-40, 
    3.080842e-37, 5.857428e-43, 2.656862e-42, 3.865622e-41, 1.357889e-38, 
    6.010099e-40, 2.277948e-38, 6.06482e-42, 6.305843e-44, 1.821688e-44, 
    1.401298e-45, 1.961818e-44, 1.681558e-44, 1.485376e-43, 7.286752e-44, 
    1.275882e-41, 8.253648e-43, 1.617401e-39, 2.214481e-38, 2.374424e-35, 
    1.282891e-33, 6.005723e-32, 3.070762e-31, 5.006057e-31, 6.134316e-31,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 7.861284e-43, 0, 
    3.210375e-42, 6.417947e-43, 7.479431e-41, 1.96406e-41, 6.575739e-39, 
    1.376832e-40, 1.144394e-37, 2.654452e-39, 4.841027e-39, 1.208312e-40, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.149065e-43, 7.006492e-45, 
    2.077565e-41, 2.918905e-42, 1.896657e-41, 1.0797e-41, 1.91053e-41, 
    1.055178e-42, 3.69102e-42, 2.760558e-43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2.031883e-43, 6.866362e-44, 4.301986e-43, 2.394819e-42, 
    3.987395e-41, 2.52514e-41, 8.530545e-41, 4.091792e-43, 1.475287e-41, 
    3.643376e-44, 1.975831e-43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.963219e-42, 8.547921e-44, 4.09039e-42, 5.815389e-43, 1.604206e-41, 
    8.141544e-43, 1.335914e-40, 3.902098e-40, 1.878609e-40, 3.006833e-39, 
    6.880375e-43, 1.896938e-41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.802597e-45, 1.050974e-43, 1.317221e-42, 2.830623e-43, 1.101421e-42, 
    2.410233e-43, 1.163078e-43, 2.61586e-40, 3.73446e-42, 2.029436e-39, 
    1.449554e-39, 8.779976e-41, 1.505666e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1.401298e-45, 5.745324e-44, 2.64425e-42, 2.008061e-42, 2.21265e-42, 
    5.099325e-42, 6.361895e-43, 7.14382e-42, 1.065547e-41, 3.731658e-42, 
    1.385541e-39, 2.663966e-40, 1.439199e-39, 4.939493e-40, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.484155e-44, 0, 5.26608e-42, 2.101948e-44, 
    7.377836e-42, 2.60081e-42, 1.451605e-41, 6.5833e-41, 4.248387e-40, 
    1.192297e-38, 5.575409e-39, 8.385329e-38, 0, 0, 0, 0, 0, 0, 2.802597e-45, 
    0, 1.401298e-44, 2.802597e-44, 0, 2.802597e-45, 0, 0, 0, 0, 0, 0, 
    1.121039e-43, 4.203895e-45, 5.315405e-41, 5.240856e-43, 3.658001e-39, 
    1.228313e-37, 2.908488e-36, 9.948723e-35, 0, 0, 0, 0, 0, 4.203895e-45, 
    7.006492e-45, 1.541428e-44, 1.079e-43, 5.394999e-43, 1.961818e-44, 
    8.02944e-43, 0, 1.401298e-45, 0, 0, 0, 0, 0, 1.401298e-45, 2.186026e-43, 
    1.401298e-44, 5.237218e-38, 9.034031e-41, 1.30194e-33, 1.866296e-35, 0, 
    0, 0, 0, 5.605194e-45, 4.904545e-44, 2.606415e-43, 2.080928e-42, 
    2.596606e-42, 8.671235e-42, 1.192505e-42, 8.022434e-42, 4.203895e-45, 
    1.415311e-43, 0, 0, 0, 0, 0, 2.101948e-44, 2.242078e-44, 7.426882e-44, 
    2.022074e-42, 7.006492e-45, 1.149747e-37, 5.598187e-42, 0, 0, 0, 0, 
    4.063766e-44, 1.401298e-45, 8.420402e-42, 8.814167e-43, 3.454061e-41, 
    5.686469e-42, 4.348229e-42, 4.021727e-43, 8.82818e-44, 1.401298e-45, 0, 
    0, 0, 0, 2.662467e-44, 2.649855e-42, 9.809089e-43, 2.627575e-41, 
    2.802597e-45, 1.59748e-43, 3.643376e-44, 1.633914e-42, 0, 4.83448e-43, 0, 
    0, 1.401298e-45, 2.059909e-43, 6.025583e-43, 1.863727e-42, 9.290609e-43, 
    2.942727e-44, 1.681558e-44, 1.401298e-45, 0, 0, 0, 0, 0, 2.942727e-44, 
    1.296201e-42, 6.725672e-41, 1.721047e-40, 1.329927e-38, 3.933921e-40, 
    1.211254e-37, 9.539564e-40, 3.477869e-36, 7.258726e-43, 8.226813e-40, 
    1.401298e-45, 7.006492e-45, 1.036961e-43, 3.626e-41, 1.604487e-42, 
    6.082897e-41, 1.681558e-44, 0, 0, 0, 0, 0, 0, 0, 3.363116e-44, 
    2.802597e-45, 4.318802e-42, 5.913339e-41, 6.340457e-38, 3.425724e-36, 
    1.603717e-34, 8.199902e-34, 1.336775e-33, 1.638055e-33 ;

 F_N2O_NIT =
  2.302583e-14, 2.322413e-14, 2.31855e-14, 2.334595e-14, 2.325687e-14, 
    2.336203e-14, 2.306595e-14, 2.323199e-14, 2.312592e-14, 2.304362e-14, 
    2.365893e-14, 2.33531e-14, 2.397887e-14, 2.378218e-14, 2.427788e-14, 
    2.394819e-14, 2.434465e-14, 2.426834e-14, 2.449839e-14, 2.443236e-14, 
    2.472783e-14, 2.452888e-14, 2.488173e-14, 2.468024e-14, 2.471169e-14, 
    2.452232e-14, 2.341451e-14, 2.362076e-14, 2.340231e-14, 2.343166e-14, 
    2.341848e-14, 2.32587e-14, 2.317838e-14, 2.301069e-14, 2.304108e-14, 
    2.316428e-14, 2.344484e-14, 2.33494e-14, 2.359032e-14, 2.358487e-14, 
    2.385456e-14, 2.373276e-14, 2.418848e-14, 2.405849e-14, 2.443511e-14, 
    2.43401e-14, 2.443064e-14, 2.440316e-14, 2.443099e-14, 2.429173e-14, 
    2.435134e-14, 2.422899e-14, 2.375558e-14, 2.389421e-14, 2.348197e-14, 
    2.323588e-14, 2.30732e-14, 2.295812e-14, 2.297437e-14, 2.300536e-14, 
    2.316499e-14, 2.331561e-14, 2.343073e-14, 2.35079e-14, 2.358407e-14, 
    2.38154e-14, 2.393834e-14, 2.421479e-14, 2.416479e-14, 2.424954e-14, 
    2.433066e-14, 2.446716e-14, 2.444467e-14, 2.45049e-14, 2.424729e-14, 
    2.441833e-14, 2.41363e-14, 2.421327e-14, 2.36048e-14, 2.337514e-14, 
    2.327786e-14, 2.31929e-14, 2.298686e-14, 2.312904e-14, 2.307293e-14, 
    2.320652e-14, 2.329162e-14, 2.324951e-14, 2.351001e-14, 2.340855e-14, 
    2.394563e-14, 2.371351e-14, 2.432119e-14, 2.417504e-14, 2.435628e-14, 
    2.426371e-14, 2.442243e-14, 2.427956e-14, 2.452734e-14, 2.458146e-14, 
    2.454446e-14, 2.468675e-14, 2.427163e-14, 2.443061e-14, 2.324834e-14, 
    2.325521e-14, 2.32872e-14, 2.314672e-14, 2.313814e-14, 2.300984e-14, 
    2.312398e-14, 2.317268e-14, 2.329655e-14, 2.336997e-14, 2.343988e-14, 
    2.359399e-14, 2.376672e-14, 2.400936e-14, 2.41845e-14, 2.430226e-14, 
    2.423001e-14, 2.429378e-14, 2.422249e-14, 2.418911e-14, 2.456117e-14, 
    2.435188e-14, 2.466625e-14, 2.46488e-14, 2.450631e-14, 2.465076e-14, 
    2.326002e-14, 2.322053e-14, 2.308368e-14, 2.319074e-14, 2.299588e-14, 
    2.310484e-14, 2.316761e-14, 2.341065e-14, 2.346424e-14, 2.351398e-14, 
    2.361237e-14, 2.373896e-14, 2.39619e-14, 2.415676e-14, 2.433537e-14, 
    2.432226e-14, 2.432687e-14, 2.436685e-14, 2.426786e-14, 2.438312e-14, 
    2.440248e-14, 2.435185e-14, 2.464645e-14, 2.45621e-14, 2.464842e-14, 
    2.459347e-14, 2.323336e-14, 2.329984e-14, 2.32639e-14, 2.33315e-14, 
    2.328386e-14, 2.349608e-14, 2.35599e-14, 2.385977e-14, 2.373647e-14, 
    2.393287e-14, 2.375638e-14, 2.37876e-14, 2.393927e-14, 2.376589e-14, 
    2.414598e-14, 2.388793e-14, 2.43684e-14, 2.410946e-14, 2.438467e-14, 
    2.433458e-14, 2.441754e-14, 2.449197e-14, 2.458578e-14, 2.475937e-14, 
    2.471911e-14, 2.486465e-14, 2.339914e-14, 2.348572e-14, 2.347809e-14, 
    2.356886e-14, 2.36361e-14, 2.378221e-14, 2.401752e-14, 2.392888e-14, 
    2.409173e-14, 2.412449e-14, 2.387713e-14, 2.402884e-14, 2.354373e-14, 
    2.362174e-14, 2.357527e-14, 2.340592e-14, 2.394926e-14, 2.366959e-14, 
    2.418736e-14, 2.403485e-14, 2.448134e-14, 2.425875e-14, 2.469696e-14, 
    2.488553e-14, 2.506373e-14, 2.527277e-14, 2.353304e-14, 2.347413e-14, 
    2.357966e-14, 2.372607e-14, 2.386236e-14, 2.404417e-14, 2.406282e-14, 
    2.409696e-14, 2.418555e-14, 2.426017e-14, 2.410776e-14, 2.427889e-14, 
    2.363984e-14, 2.397362e-14, 2.345184e-14, 2.360831e-14, 2.371739e-14, 
    2.366951e-14, 2.391873e-14, 2.397766e-14, 2.421793e-14, 2.409357e-14, 
    2.483891e-14, 2.450768e-14, 2.543257e-14, 2.517229e-14, 2.345356e-14, 
    2.353283e-14, 2.38098e-14, 2.367781e-14, 2.405633e-14, 2.414999e-14, 
    2.422626e-14, 2.432394e-14, 2.43345e-14, 2.439249e-14, 2.42975e-14, 
    2.438873e-14, 2.404453e-14, 2.419803e-14, 2.377803e-14, 2.387989e-14, 
    2.383301e-14, 2.378162e-14, 2.394038e-14, 2.411012e-14, 2.411376e-14, 
    2.416832e-14, 2.43224e-14, 2.405782e-14, 2.48818e-14, 2.437119e-14, 
    2.361943e-14, 2.377279e-14, 2.379475e-14, 2.373524e-14, 2.414058e-14, 
    2.399329e-14, 2.439107e-14, 2.428323e-14, 2.446006e-14, 2.43721e-14, 
    2.435917e-14, 2.424648e-14, 2.417645e-14, 2.400001e-14, 2.385695e-14, 
    2.374384e-14, 2.377011e-14, 2.389445e-14, 2.412052e-14, 2.433542e-14, 
    2.428825e-14, 2.444656e-14, 2.402872e-14, 2.420346e-14, 2.413584e-14, 
    2.431236e-14, 2.392652e-14, 2.42549e-14, 2.384295e-14, 2.387892e-14, 
    2.399037e-14, 2.421537e-14, 2.426531e-14, 2.431868e-14, 2.428574e-14, 
    2.412629e-14, 2.410022e-14, 2.398764e-14, 2.395659e-14, 2.387106e-14, 
    2.380035e-14, 2.386494e-14, 2.393286e-14, 2.412634e-14, 2.430139e-14, 
    2.4493e-14, 2.454001e-14, 2.476509e-14, 2.458177e-14, 2.488464e-14, 
    2.462699e-14, 2.50739e-14, 2.427401e-14, 2.461951e-14, 2.399545e-14, 
    2.406227e-14, 2.418339e-14, 2.446239e-14, 2.431157e-14, 2.448801e-14, 
    2.40992e-14, 2.389875e-14, 2.384704e-14, 2.37507e-14, 2.384923e-14, 
    2.384121e-14, 2.393568e-14, 2.39053e-14, 2.413277e-14, 2.401044e-14, 
    2.43588e-14, 2.448658e-14, 2.484934e-14, 2.507309e-14, 2.530196e-14, 
    2.540334e-14, 2.543424e-14, 2.544716e-14 ;

 F_NIT =
  3.837638e-11, 3.870687e-11, 3.864251e-11, 3.890991e-11, 3.876146e-11, 
    3.893671e-11, 3.844325e-11, 3.871999e-11, 3.85432e-11, 3.840604e-11, 
    3.943156e-11, 3.892183e-11, 3.996478e-11, 3.963697e-11, 4.046314e-11, 
    3.991366e-11, 4.057441e-11, 4.044724e-11, 4.083065e-11, 4.072061e-11, 
    4.121304e-11, 4.088148e-11, 4.146955e-11, 4.113373e-11, 4.118616e-11, 
    4.087053e-11, 3.902418e-11, 3.936794e-11, 3.900385e-11, 3.905276e-11, 
    3.903081e-11, 3.87645e-11, 3.863064e-11, 3.835115e-11, 3.84018e-11, 
    3.860712e-11, 3.907473e-11, 3.891567e-11, 3.93172e-11, 3.930811e-11, 
    3.97576e-11, 3.95546e-11, 4.031413e-11, 4.009748e-11, 4.072519e-11, 
    4.056684e-11, 4.071773e-11, 4.067194e-11, 4.071832e-11, 4.048622e-11, 
    4.058556e-11, 4.038165e-11, 3.959263e-11, 3.982369e-11, 3.913661e-11, 
    3.872647e-11, 3.845534e-11, 3.826354e-11, 3.829061e-11, 3.834227e-11, 
    3.860832e-11, 3.885935e-11, 3.905122e-11, 3.917984e-11, 3.930679e-11, 
    3.969234e-11, 3.989723e-11, 4.035799e-11, 4.027464e-11, 4.041589e-11, 
    4.05511e-11, 4.077861e-11, 4.074111e-11, 4.08415e-11, 4.041215e-11, 
    4.069722e-11, 4.022717e-11, 4.035544e-11, 3.934133e-11, 3.895857e-11, 
    3.879643e-11, 3.865483e-11, 3.831144e-11, 3.85484e-11, 3.845489e-11, 
    3.867754e-11, 3.881936e-11, 3.874918e-11, 3.918335e-11, 3.901425e-11, 
    3.990938e-11, 3.952251e-11, 4.053532e-11, 4.029174e-11, 4.059381e-11, 
    4.043952e-11, 4.070406e-11, 4.046593e-11, 4.087889e-11, 4.096911e-11, 
    4.090744e-11, 4.114458e-11, 4.045272e-11, 4.071768e-11, 3.874724e-11, 
    3.875868e-11, 3.8812e-11, 3.857787e-11, 3.856357e-11, 3.834973e-11, 
    3.853997e-11, 3.862113e-11, 3.882758e-11, 3.894995e-11, 3.906647e-11, 
    3.932332e-11, 3.96112e-11, 4.001561e-11, 4.030749e-11, 4.050376e-11, 
    4.038335e-11, 4.048964e-11, 4.037082e-11, 4.031519e-11, 4.093528e-11, 
    4.058647e-11, 4.111041e-11, 4.108133e-11, 4.084385e-11, 4.108459e-11, 
    3.87667e-11, 3.870088e-11, 3.847281e-11, 3.865122e-11, 3.832647e-11, 
    3.850806e-11, 3.861268e-11, 3.901776e-11, 3.910706e-11, 3.918996e-11, 
    3.935395e-11, 3.956494e-11, 3.99365e-11, 4.026126e-11, 4.055896e-11, 
    4.053709e-11, 4.054479e-11, 4.061142e-11, 4.044644e-11, 4.063853e-11, 
    4.06708e-11, 4.058642e-11, 4.107742e-11, 4.093683e-11, 4.108069e-11, 
    4.098911e-11, 3.872226e-11, 3.883307e-11, 3.877316e-11, 3.888584e-11, 
    3.880643e-11, 3.916014e-11, 3.926651e-11, 3.976628e-11, 3.956078e-11, 
    3.988811e-11, 3.959396e-11, 3.964599e-11, 3.989878e-11, 3.960982e-11, 
    4.024329e-11, 3.981321e-11, 4.061401e-11, 4.018243e-11, 4.064112e-11, 
    4.055763e-11, 4.06959e-11, 4.081996e-11, 4.09763e-11, 4.126561e-11, 
    4.119851e-11, 4.144108e-11, 3.899858e-11, 3.914286e-11, 3.913015e-11, 
    3.928143e-11, 3.93935e-11, 3.963701e-11, 4.00292e-11, 3.988147e-11, 
    4.015288e-11, 4.020748e-11, 3.979522e-11, 4.004806e-11, 3.923955e-11, 
    3.936957e-11, 3.929213e-11, 3.900987e-11, 3.991543e-11, 3.944932e-11, 
    4.031227e-11, 4.005809e-11, 4.080224e-11, 4.043125e-11, 4.11616e-11, 
    4.147589e-11, 4.177288e-11, 4.212129e-11, 3.922173e-11, 3.912355e-11, 
    3.929944e-11, 3.954346e-11, 3.97706e-11, 4.007362e-11, 4.010469e-11, 
    4.016161e-11, 4.030926e-11, 4.043362e-11, 4.017959e-11, 4.046481e-11, 
    3.939973e-11, 3.995603e-11, 3.908639e-11, 3.934719e-11, 3.952899e-11, 
    3.944919e-11, 3.986455e-11, 3.996277e-11, 4.036321e-11, 4.015595e-11, 
    4.139818e-11, 4.084614e-11, 4.238762e-11, 4.195382e-11, 3.908927e-11, 
    3.922138e-11, 3.968301e-11, 3.946301e-11, 4.009388e-11, 4.024997e-11, 
    4.03771e-11, 4.05399e-11, 4.05575e-11, 4.065415e-11, 4.049583e-11, 
    4.064788e-11, 4.007421e-11, 4.033004e-11, 3.963006e-11, 3.979982e-11, 
    3.972167e-11, 3.963604e-11, 3.990063e-11, 4.018353e-11, 4.018959e-11, 
    4.028053e-11, 4.053733e-11, 4.009636e-11, 4.146967e-11, 4.061865e-11, 
    3.936571e-11, 3.962132e-11, 3.965791e-11, 3.955874e-11, 4.02343e-11, 
    3.998882e-11, 4.065179e-11, 4.047205e-11, 4.076676e-11, 4.062017e-11, 
    4.059861e-11, 4.04108e-11, 4.029408e-11, 4.000002e-11, 3.976158e-11, 
    3.957306e-11, 3.961685e-11, 3.982409e-11, 4.020086e-11, 4.055902e-11, 
    4.048042e-11, 4.074426e-11, 4.004787e-11, 4.03391e-11, 4.02264e-11, 
    4.05206e-11, 3.987753e-11, 4.042483e-11, 3.973825e-11, 3.97982e-11, 
    3.998394e-11, 4.035896e-11, 4.044219e-11, 4.053113e-11, 4.047623e-11, 
    4.021049e-11, 4.016704e-11, 3.997939e-11, 3.992765e-11, 3.97851e-11, 
    3.966726e-11, 3.97749e-11, 3.98881e-11, 4.021057e-11, 4.050232e-11, 
    4.082166e-11, 4.090002e-11, 4.127515e-11, 4.096961e-11, 4.147441e-11, 
    4.104499e-11, 4.178983e-11, 4.045668e-11, 4.103252e-11, 3.999241e-11, 
    4.010379e-11, 4.030565e-11, 4.077065e-11, 4.051928e-11, 4.081335e-11, 
    4.016533e-11, 3.983125e-11, 3.974506e-11, 3.95845e-11, 3.974873e-11, 
    3.973535e-11, 3.989281e-11, 3.984217e-11, 4.022128e-11, 4.00174e-11, 
    4.0598e-11, 4.081097e-11, 4.141557e-11, 4.178849e-11, 4.216993e-11, 
    4.23389e-11, 4.23904e-11, 4.241194e-11 ;

 F_NIT_vr =
  2.454741e-10, 2.465639e-10, 2.463515e-10, 2.47231e-10, 2.467428e-10, 
    2.473182e-10, 2.456938e-10, 2.466052e-10, 2.46023e-10, 2.455701e-10, 
    2.489369e-10, 2.472681e-10, 2.506745e-10, 2.496075e-10, 2.52289e-10, 
    2.505075e-10, 2.526483e-10, 2.522372e-10, 2.534745e-10, 2.531195e-10, 
    2.547023e-10, 2.536375e-10, 2.55524e-10, 2.544477e-10, 2.546155e-10, 
    2.53601e-10, 2.47606e-10, 2.487309e-10, 2.475388e-10, 2.476992e-10, 
    2.47627e-10, 2.467516e-10, 2.463107e-10, 2.453887e-10, 2.455557e-10, 
    2.462327e-10, 2.477693e-10, 2.472472e-10, 2.48563e-10, 2.485333e-10, 
    2.499995e-10, 2.49338e-10, 2.518062e-10, 2.511037e-10, 2.53134e-10, 
    2.526225e-10, 2.531093e-10, 2.529613e-10, 2.531105e-10, 2.523612e-10, 
    2.526816e-10, 2.520227e-10, 2.49465e-10, 2.502172e-10, 2.479736e-10, 
    2.466259e-10, 2.457326e-10, 2.450992e-10, 2.451881e-10, 2.453588e-10, 
    2.462361e-10, 2.47062e-10, 2.476919e-10, 2.48113e-10, 2.485283e-10, 
    2.497862e-10, 2.504531e-10, 2.519475e-10, 2.516778e-10, 2.521343e-10, 
    2.525714e-10, 2.53305e-10, 2.531841e-10, 2.53507e-10, 2.521211e-10, 
    2.530417e-10, 2.515218e-10, 2.519372e-10, 2.486426e-10, 2.473892e-10, 
    2.468558e-10, 2.463899e-10, 2.452567e-10, 2.460389e-10, 2.457301e-10, 
    2.464638e-10, 2.469303e-10, 2.466991e-10, 2.481242e-10, 2.475694e-10, 
    2.504922e-10, 2.492322e-10, 2.525208e-10, 2.517325e-10, 2.52709e-10, 
    2.522106e-10, 2.530641e-10, 2.522954e-10, 2.53627e-10, 2.539171e-10, 
    2.537182e-10, 2.544807e-10, 2.522511e-10, 2.531065e-10, 2.466942e-10, 
    2.467318e-10, 2.469069e-10, 2.461356e-10, 2.460884e-10, 2.453824e-10, 
    2.4601e-10, 2.462774e-10, 2.469567e-10, 2.473582e-10, 2.477402e-10, 
    2.485814e-10, 2.49521e-10, 2.508367e-10, 2.517833e-10, 2.524178e-10, 
    2.520284e-10, 2.523717e-10, 2.519873e-10, 2.518069e-10, 2.538076e-10, 
    2.526835e-10, 2.543702e-10, 2.542769e-10, 2.535125e-10, 2.542866e-10, 
    2.467577e-10, 2.465408e-10, 2.457889e-10, 2.463768e-10, 2.453051e-10, 
    2.459045e-10, 2.462489e-10, 2.475804e-10, 2.478732e-10, 2.481448e-10, 
    2.486811e-10, 2.493698e-10, 2.505794e-10, 2.516329e-10, 2.525958e-10, 
    2.525248e-10, 2.525495e-10, 2.527642e-10, 2.522312e-10, 2.528512e-10, 
    2.529549e-10, 2.526828e-10, 2.542636e-10, 2.538116e-10, 2.542738e-10, 
    2.539791e-10, 2.466109e-10, 2.469749e-10, 2.467776e-10, 2.47148e-10, 
    2.468864e-10, 2.480471e-10, 2.48395e-10, 2.50026e-10, 2.493561e-10, 
    2.504222e-10, 2.494639e-10, 2.496336e-10, 2.504556e-10, 2.49515e-10, 
    2.515736e-10, 2.501765e-10, 2.527723e-10, 2.513752e-10, 2.528593e-10, 
    2.525894e-10, 2.530354e-10, 2.534351e-10, 2.539378e-10, 2.548667e-10, 
    2.54651e-10, 2.554285e-10, 2.475182e-10, 2.479908e-10, 2.479492e-10, 
    2.484442e-10, 2.488103e-10, 2.496053e-10, 2.508808e-10, 2.504005e-10, 
    2.512816e-10, 2.514585e-10, 2.501191e-10, 2.509408e-10, 2.483048e-10, 
    2.487295e-10, 2.484765e-10, 2.475512e-10, 2.505084e-10, 2.489892e-10, 
    2.517956e-10, 2.509712e-10, 2.533773e-10, 2.521797e-10, 2.545324e-10, 
    2.555392e-10, 2.564882e-10, 2.575969e-10, 2.482489e-10, 2.47927e-10, 
    2.485026e-10, 2.492996e-10, 2.500396e-10, 2.510247e-10, 2.511253e-10, 
    2.513094e-10, 2.517876e-10, 2.5219e-10, 2.513669e-10, 2.522902e-10, 
    2.488273e-10, 2.506404e-10, 2.478018e-10, 2.486554e-10, 2.492489e-10, 
    2.489886e-10, 2.503422e-10, 2.506611e-10, 2.51959e-10, 2.512879e-10, 
    2.552896e-10, 2.535172e-10, 2.584422e-10, 2.570637e-10, 2.478144e-10, 
    2.482468e-10, 2.49754e-10, 2.490366e-10, 2.510898e-10, 2.515959e-10, 
    2.52007e-10, 2.525332e-10, 2.525896e-10, 2.529016e-10, 2.523899e-10, 
    2.528809e-10, 2.510238e-10, 2.518532e-10, 2.495789e-10, 2.501314e-10, 
    2.49877e-10, 2.495975e-10, 2.504586e-10, 2.513768e-10, 2.513964e-10, 
    2.516905e-10, 2.525199e-10, 2.510931e-10, 2.555168e-10, 2.527817e-10, 
    2.487187e-10, 2.495524e-10, 2.496717e-10, 2.493485e-10, 2.515443e-10, 
    2.50748e-10, 2.52894e-10, 2.523132e-10, 2.532641e-10, 2.527913e-10, 
    2.527211e-10, 2.521144e-10, 2.51736e-10, 2.507823e-10, 2.500064e-10, 
    2.493922e-10, 2.495344e-10, 2.502093e-10, 2.514322e-10, 2.525913e-10, 
    2.523369e-10, 2.531884e-10, 2.509352e-10, 2.518792e-10, 2.515135e-10, 
    2.524657e-10, 2.503865e-10, 2.521605e-10, 2.499331e-10, 2.501279e-10, 
    2.507314e-10, 2.51947e-10, 2.522161e-10, 2.525035e-10, 2.523257e-10, 
    2.514654e-10, 2.513243e-10, 2.50715e-10, 2.505464e-10, 2.50083e-10, 
    2.496986e-10, 2.500492e-10, 2.504168e-10, 2.514638e-10, 2.524075e-10, 
    2.534374e-10, 2.536897e-10, 2.548935e-10, 2.539125e-10, 2.555306e-10, 
    2.541534e-10, 2.565381e-10, 2.522632e-10, 2.541193e-10, 2.507591e-10, 
    2.511203e-10, 2.51774e-10, 2.532756e-10, 2.524646e-10, 2.53413e-10, 
    2.513187e-10, 2.502329e-10, 2.499523e-10, 2.494291e-10, 2.499638e-10, 
    2.499203e-10, 2.504324e-10, 2.502673e-10, 2.514978e-10, 2.508365e-10, 
    2.527157e-10, 2.534024e-10, 2.553437e-10, 2.565348e-10, 2.577494e-10, 
    2.582854e-10, 2.584487e-10, 2.585166e-10,
  1.247084e-10, 1.256584e-10, 1.254736e-10, 1.262413e-10, 1.258153e-10, 
    1.263183e-10, 1.249009e-10, 1.256961e-10, 1.251883e-10, 1.247939e-10, 
    1.277361e-10, 1.262756e-10, 1.292607e-10, 1.283242e-10, 1.306818e-10, 
    1.291147e-10, 1.309987e-10, 1.306367e-10, 1.317279e-10, 1.31415e-10, 
    1.328139e-10, 1.318724e-10, 1.335415e-10, 1.325889e-10, 1.327377e-10, 
    1.318414e-10, 1.265692e-10, 1.275538e-10, 1.265109e-10, 1.266511e-10, 
    1.265883e-10, 1.25824e-10, 1.254394e-10, 1.24636e-10, 1.247818e-10, 
    1.25372e-10, 1.267142e-10, 1.262581e-10, 1.274092e-10, 1.273832e-10, 
    1.286691e-10, 1.280887e-10, 1.302575e-10, 1.296397e-10, 1.31428e-10, 
    1.309774e-10, 1.314068e-10, 1.312766e-10, 1.314085e-10, 1.307479e-10, 
    1.310308e-10, 1.3045e-10, 1.281973e-10, 1.288577e-10, 1.268916e-10, 
    1.257146e-10, 1.249357e-10, 1.243839e-10, 1.244619e-10, 1.246105e-10, 
    1.253754e-10, 1.260965e-10, 1.26647e-10, 1.270157e-10, 1.273794e-10, 
    1.284823e-10, 1.290679e-10, 1.303824e-10, 1.30145e-10, 1.305475e-10, 
    1.309326e-10, 1.3158e-10, 1.314734e-10, 1.317588e-10, 1.30537e-10, 
    1.313485e-10, 1.300098e-10, 1.303754e-10, 1.274777e-10, 1.263811e-10, 
    1.259155e-10, 1.255091e-10, 1.245218e-10, 1.252032e-10, 1.249344e-10, 
    1.255745e-10, 1.259817e-10, 1.257802e-10, 1.270258e-10, 1.26541e-10, 
    1.291026e-10, 1.279968e-10, 1.308877e-10, 1.301937e-10, 1.310542e-10, 
    1.306149e-10, 1.313679e-10, 1.306902e-10, 1.318652e-10, 1.321215e-10, 
    1.319463e-10, 1.326199e-10, 1.306526e-10, 1.314067e-10, 1.257746e-10, 
    1.258074e-10, 1.259605e-10, 1.252879e-10, 1.252469e-10, 1.24632e-10, 
    1.251791e-10, 1.254123e-10, 1.260054e-10, 1.263565e-10, 1.266907e-10, 
    1.274267e-10, 1.282505e-10, 1.29406e-10, 1.302387e-10, 1.307979e-10, 
    1.304549e-10, 1.307577e-10, 1.304192e-10, 1.302607e-10, 1.320254e-10, 
    1.310334e-10, 1.32523e-10, 1.324404e-10, 1.317656e-10, 1.324497e-10, 
    1.258305e-10, 1.256415e-10, 1.24986e-10, 1.254989e-10, 1.245651e-10, 
    1.250874e-10, 1.25388e-10, 1.265509e-10, 1.268072e-10, 1.270447e-10, 
    1.275145e-10, 1.281184e-10, 1.291802e-10, 1.301069e-10, 1.309551e-10, 
    1.308929e-10, 1.309148e-10, 1.311044e-10, 1.306347e-10, 1.311816e-10, 
    1.312734e-10, 1.310333e-10, 1.324293e-10, 1.320299e-10, 1.324386e-10, 
    1.321786e-10, 1.257029e-10, 1.260211e-10, 1.258491e-10, 1.261725e-10, 
    1.259446e-10, 1.269591e-10, 1.272639e-10, 1.286939e-10, 1.281064e-10, 
    1.29042e-10, 1.282014e-10, 1.283501e-10, 1.290723e-10, 1.282468e-10, 
    1.300556e-10, 1.28828e-10, 1.311118e-10, 1.298819e-10, 1.31189e-10, 
    1.309514e-10, 1.313449e-10, 1.316977e-10, 1.321421e-10, 1.329634e-10, 
    1.327731e-10, 1.334611e-10, 1.26496e-10, 1.269096e-10, 1.268733e-10, 
    1.273068e-10, 1.276277e-10, 1.283245e-10, 1.294449e-10, 1.290232e-10, 
    1.297979e-10, 1.299536e-10, 1.287768e-10, 1.294987e-10, 1.271869e-10, 
    1.275592e-10, 1.273375e-10, 1.265286e-10, 1.291201e-10, 1.277875e-10, 
    1.302524e-10, 1.295275e-10, 1.316474e-10, 1.305914e-10, 1.326683e-10, 
    1.335596e-10, 1.344009e-10, 1.353859e-10, 1.271358e-10, 1.268544e-10, 
    1.273584e-10, 1.280568e-10, 1.287064e-10, 1.295717e-10, 1.296604e-10, 
    1.298228e-10, 1.302438e-10, 1.305982e-10, 1.29874e-10, 1.306871e-10, 
    1.276453e-10, 1.292361e-10, 1.26748e-10, 1.274951e-10, 1.280156e-10, 
    1.277873e-10, 1.28975e-10, 1.292555e-10, 1.303976e-10, 1.298068e-10, 
    1.333393e-10, 1.317721e-10, 1.36138e-10, 1.349127e-10, 1.267562e-10, 
    1.271348e-10, 1.284559e-10, 1.278267e-10, 1.296296e-10, 1.300748e-10, 
    1.304372e-10, 1.309008e-10, 1.30951e-10, 1.31226e-10, 1.307754e-10, 
    1.312083e-10, 1.295735e-10, 1.303031e-10, 1.283048e-10, 1.2879e-10, 
    1.285668e-10, 1.28322e-10, 1.290781e-10, 1.298853e-10, 1.299028e-10, 
    1.30162e-10, 1.308931e-10, 1.296369e-10, 1.335416e-10, 1.311247e-10, 
    1.275482e-10, 1.282795e-10, 1.283843e-10, 1.281007e-10, 1.300301e-10, 
    1.293297e-10, 1.312193e-10, 1.307077e-10, 1.315465e-10, 1.311294e-10, 
    1.310681e-10, 1.305333e-10, 1.302006e-10, 1.293618e-10, 1.286808e-10, 
    1.281419e-10, 1.282671e-10, 1.288594e-10, 1.299348e-10, 1.309554e-10, 
    1.307316e-10, 1.314826e-10, 1.294985e-10, 1.30329e-10, 1.300077e-10, 
    1.308462e-10, 1.290119e-10, 1.305726e-10, 1.28614e-10, 1.287854e-10, 
    1.293158e-10, 1.303853e-10, 1.306227e-10, 1.308759e-10, 1.307197e-10, 
    1.299622e-10, 1.298384e-10, 1.29303e-10, 1.291552e-10, 1.287481e-10, 
    1.284113e-10, 1.287189e-10, 1.290423e-10, 1.299626e-10, 1.30794e-10, 
    1.317027e-10, 1.319255e-10, 1.329903e-10, 1.32123e-10, 1.335551e-10, 
    1.323368e-10, 1.344486e-10, 1.306636e-10, 1.323014e-10, 1.293401e-10, 
    1.29658e-10, 1.302334e-10, 1.315573e-10, 1.308422e-10, 1.316788e-10, 
    1.298335e-10, 1.288797e-10, 1.286337e-10, 1.281746e-10, 1.286442e-10, 
    1.286059e-10, 1.290558e-10, 1.289112e-10, 1.299932e-10, 1.294116e-10, 
    1.310665e-10, 1.316723e-10, 1.333889e-10, 1.344451e-10, 1.355237e-10, 
    1.360008e-10, 1.361461e-10, 1.362069e-10,
  1.174451e-10, 1.184872e-10, 1.182844e-10, 1.191271e-10, 1.186593e-10, 
    1.192116e-10, 1.176561e-10, 1.185286e-10, 1.179714e-10, 1.175389e-10, 
    1.207697e-10, 1.191648e-10, 1.224471e-10, 1.214163e-10, 1.24013e-10, 
    1.222864e-10, 1.243625e-10, 1.239632e-10, 1.251668e-10, 1.248215e-10, 
    1.263661e-10, 1.253263e-10, 1.271701e-10, 1.261175e-10, 1.262819e-10, 
    1.252921e-10, 1.194871e-10, 1.205694e-10, 1.194231e-10, 1.195772e-10, 
    1.195081e-10, 1.186689e-10, 1.18247e-10, 1.173657e-10, 1.175255e-10, 
    1.181729e-10, 1.196465e-10, 1.191455e-10, 1.204101e-10, 1.203815e-10, 
    1.217958e-10, 1.211573e-10, 1.235452e-10, 1.228645e-10, 1.248359e-10, 
    1.243389e-10, 1.248125e-10, 1.246688e-10, 1.248144e-10, 1.240858e-10, 
    1.243977e-10, 1.237574e-10, 1.212767e-10, 1.220035e-10, 1.198413e-10, 
    1.18549e-10, 1.176943e-10, 1.170894e-10, 1.171748e-10, 1.173377e-10, 
    1.181767e-10, 1.18968e-10, 1.195725e-10, 1.199776e-10, 1.203773e-10, 
    1.215904e-10, 1.222349e-10, 1.236829e-10, 1.234212e-10, 1.238648e-10, 
    1.242895e-10, 1.250036e-10, 1.24886e-10, 1.25201e-10, 1.238532e-10, 
    1.247482e-10, 1.232722e-10, 1.236751e-10, 1.204857e-10, 1.192806e-10, 
    1.187695e-10, 1.183233e-10, 1.172405e-10, 1.179878e-10, 1.17693e-10, 
    1.18395e-10, 1.18842e-10, 1.186209e-10, 1.199887e-10, 1.194561e-10, 
    1.222731e-10, 1.210563e-10, 1.242399e-10, 1.234749e-10, 1.244236e-10, 
    1.239391e-10, 1.247697e-10, 1.240221e-10, 1.253184e-10, 1.256013e-10, 
    1.254079e-10, 1.261517e-10, 1.239807e-10, 1.248125e-10, 1.186146e-10, 
    1.186507e-10, 1.188188e-10, 1.180807e-10, 1.180357e-10, 1.173613e-10, 
    1.179613e-10, 1.182172e-10, 1.18868e-10, 1.192536e-10, 1.196206e-10, 
    1.204294e-10, 1.213353e-10, 1.226071e-10, 1.235244e-10, 1.241409e-10, 
    1.237628e-10, 1.240966e-10, 1.237234e-10, 1.235487e-10, 1.254952e-10, 
    1.244006e-10, 1.260446e-10, 1.259534e-10, 1.252085e-10, 1.259637e-10, 
    1.18676e-10, 1.184686e-10, 1.177495e-10, 1.183121e-10, 1.17288e-10, 
    1.178607e-10, 1.181905e-10, 1.194671e-10, 1.197485e-10, 1.200095e-10, 
    1.205259e-10, 1.211899e-10, 1.223585e-10, 1.233792e-10, 1.243142e-10, 
    1.242456e-10, 1.242697e-10, 1.24479e-10, 1.23961e-10, 1.245641e-10, 
    1.246654e-10, 1.244005e-10, 1.259412e-10, 1.255002e-10, 1.259515e-10, 
    1.256643e-10, 1.18536e-10, 1.188852e-10, 1.186965e-10, 1.190515e-10, 
    1.188013e-10, 1.199155e-10, 1.202505e-10, 1.218232e-10, 1.211768e-10, 
    1.222063e-10, 1.212812e-10, 1.214449e-10, 1.222398e-10, 1.213312e-10, 
    1.233227e-10, 1.219709e-10, 1.244871e-10, 1.231315e-10, 1.245722e-10, 
    1.243101e-10, 1.247443e-10, 1.251335e-10, 1.256241e-10, 1.265312e-10, 
    1.263209e-10, 1.270812e-10, 1.194067e-10, 1.198612e-10, 1.198212e-10, 
    1.202975e-10, 1.206504e-10, 1.214166e-10, 1.226499e-10, 1.221855e-10, 
    1.230387e-10, 1.232102e-10, 1.219144e-10, 1.227092e-10, 1.201658e-10, 
    1.205751e-10, 1.203314e-10, 1.194425e-10, 1.222924e-10, 1.208262e-10, 
    1.235396e-10, 1.227409e-10, 1.25078e-10, 1.239133e-10, 1.262052e-10, 
    1.271902e-10, 1.281205e-10, 1.292108e-10, 1.201096e-10, 1.198004e-10, 
    1.203543e-10, 1.211222e-10, 1.218368e-10, 1.227896e-10, 1.228873e-10, 
    1.230661e-10, 1.235301e-10, 1.239207e-10, 1.231226e-10, 1.240187e-10, 
    1.206699e-10, 1.2242e-10, 1.196836e-10, 1.205047e-10, 1.210769e-10, 
    1.208258e-10, 1.221325e-10, 1.224413e-10, 1.236997e-10, 1.230486e-10, 
    1.269467e-10, 1.252157e-10, 1.300439e-10, 1.286869e-10, 1.196925e-10, 
    1.201085e-10, 1.215613e-10, 1.208692e-10, 1.228533e-10, 1.233438e-10, 
    1.237432e-10, 1.242544e-10, 1.243097e-10, 1.246131e-10, 1.241161e-10, 
    1.245935e-10, 1.227916e-10, 1.235954e-10, 1.21395e-10, 1.21929e-10, 
    1.216832e-10, 1.214138e-10, 1.22246e-10, 1.231352e-10, 1.231543e-10, 
    1.2344e-10, 1.242463e-10, 1.228614e-10, 1.271706e-10, 1.245017e-10, 
    1.205629e-10, 1.213672e-10, 1.214825e-10, 1.211705e-10, 1.232946e-10, 
    1.225231e-10, 1.246057e-10, 1.240414e-10, 1.249666e-10, 1.245065e-10, 
    1.244388e-10, 1.238491e-10, 1.234825e-10, 1.225584e-10, 1.218087e-10, 
    1.212157e-10, 1.213535e-10, 1.220053e-10, 1.231897e-10, 1.243147e-10, 
    1.240678e-10, 1.248962e-10, 1.22709e-10, 1.236241e-10, 1.2327e-10, 
    1.241941e-10, 1.221732e-10, 1.238929e-10, 1.217352e-10, 1.219238e-10, 
    1.225078e-10, 1.236861e-10, 1.239477e-10, 1.242269e-10, 1.240546e-10, 
    1.232198e-10, 1.230833e-10, 1.224936e-10, 1.22331e-10, 1.218827e-10, 
    1.215121e-10, 1.218507e-10, 1.222066e-10, 1.232202e-10, 1.241366e-10, 
    1.251391e-10, 1.25385e-10, 1.265612e-10, 1.256032e-10, 1.271855e-10, 
    1.258394e-10, 1.281735e-10, 1.23993e-10, 1.258002e-10, 1.225345e-10, 
    1.228845e-10, 1.235187e-10, 1.249788e-10, 1.241898e-10, 1.251128e-10, 
    1.23078e-10, 1.220277e-10, 1.217568e-10, 1.212517e-10, 1.217684e-10, 
    1.217263e-10, 1.222215e-10, 1.220623e-10, 1.232539e-10, 1.226132e-10, 
    1.244371e-10, 1.251055e-10, 1.270014e-10, 1.281694e-10, 1.293633e-10, 
    1.298917e-10, 1.300528e-10, 1.301201e-10,
  1.205399e-10, 1.216865e-10, 1.214632e-10, 1.22391e-10, 1.218759e-10, 
    1.224841e-10, 1.207719e-10, 1.217321e-10, 1.211187e-10, 1.206429e-10, 
    1.242013e-10, 1.224325e-10, 1.260518e-10, 1.249141e-10, 1.277816e-10, 
    1.258744e-10, 1.281678e-10, 1.277264e-10, 1.290573e-10, 1.286753e-10, 
    1.303848e-10, 1.292338e-10, 1.312752e-10, 1.301095e-10, 1.302915e-10, 
    1.291959e-10, 1.227875e-10, 1.239804e-10, 1.22717e-10, 1.228867e-10, 
    1.228105e-10, 1.218865e-10, 1.214221e-10, 1.204525e-10, 1.206282e-10, 
    1.213406e-10, 1.229631e-10, 1.224112e-10, 1.238045e-10, 1.237729e-10, 
    1.253329e-10, 1.246283e-10, 1.272644e-10, 1.265125e-10, 1.286913e-10, 
    1.281416e-10, 1.286654e-10, 1.285065e-10, 1.286675e-10, 1.278619e-10, 
    1.282067e-10, 1.274989e-10, 1.247601e-10, 1.25562e-10, 1.231777e-10, 
    1.217546e-10, 1.208139e-10, 1.201485e-10, 1.202425e-10, 1.204217e-10, 
    1.213448e-10, 1.222157e-10, 1.228815e-10, 1.233278e-10, 1.237684e-10, 
    1.251064e-10, 1.258175e-10, 1.274167e-10, 1.271274e-10, 1.276177e-10, 
    1.28087e-10, 1.288768e-10, 1.287466e-10, 1.290951e-10, 1.276048e-10, 
    1.285943e-10, 1.269628e-10, 1.27408e-10, 1.238881e-10, 1.225599e-10, 
    1.219974e-10, 1.215061e-10, 1.203148e-10, 1.211369e-10, 1.208125e-10, 
    1.215849e-10, 1.22077e-10, 1.218335e-10, 1.233401e-10, 1.227533e-10, 
    1.258597e-10, 1.245171e-10, 1.280322e-10, 1.271868e-10, 1.282353e-10, 
    1.276998e-10, 1.28618e-10, 1.277914e-10, 1.29225e-10, 1.295381e-10, 
    1.293241e-10, 1.301472e-10, 1.277457e-10, 1.286654e-10, 1.218267e-10, 
    1.218664e-10, 1.220514e-10, 1.212391e-10, 1.211895e-10, 1.204477e-10, 
    1.211077e-10, 1.213893e-10, 1.221056e-10, 1.225302e-10, 1.229345e-10, 
    1.238258e-10, 1.248249e-10, 1.262284e-10, 1.272415e-10, 1.279228e-10, 
    1.275048e-10, 1.278738e-10, 1.274614e-10, 1.272683e-10, 1.294207e-10, 
    1.282099e-10, 1.300287e-10, 1.299277e-10, 1.291034e-10, 1.299391e-10, 
    1.218943e-10, 1.216659e-10, 1.208746e-10, 1.214937e-10, 1.20367e-10, 
    1.20997e-10, 1.2136e-10, 1.227655e-10, 1.230754e-10, 1.233631e-10, 
    1.239322e-10, 1.246644e-10, 1.259539e-10, 1.270811e-10, 1.281144e-10, 
    1.280385e-10, 1.280652e-10, 1.282965e-10, 1.277239e-10, 1.283907e-10, 
    1.285027e-10, 1.282098e-10, 1.299142e-10, 1.294262e-10, 1.299256e-10, 
    1.296077e-10, 1.217401e-10, 1.221246e-10, 1.219168e-10, 1.223077e-10, 
    1.220322e-10, 1.232595e-10, 1.236287e-10, 1.253631e-10, 1.246499e-10, 
    1.257859e-10, 1.247651e-10, 1.249457e-10, 1.25823e-10, 1.248202e-10, 
    1.270188e-10, 1.255261e-10, 1.283055e-10, 1.268076e-10, 1.283997e-10, 
    1.281099e-10, 1.285899e-10, 1.290205e-10, 1.295632e-10, 1.305675e-10, 
    1.303346e-10, 1.311767e-10, 1.226989e-10, 1.231996e-10, 1.231555e-10, 
    1.236805e-10, 1.240694e-10, 1.249145e-10, 1.262756e-10, 1.257629e-10, 
    1.267049e-10, 1.268944e-10, 1.254636e-10, 1.263411e-10, 1.235353e-10, 
    1.239865e-10, 1.237177e-10, 1.227383e-10, 1.258809e-10, 1.242633e-10, 
    1.272583e-10, 1.263761e-10, 1.28959e-10, 1.276713e-10, 1.302065e-10, 
    1.312976e-10, 1.323285e-10, 1.335381e-10, 1.234733e-10, 1.231326e-10, 
    1.23743e-10, 1.245898e-10, 1.253781e-10, 1.264298e-10, 1.265377e-10, 
    1.267352e-10, 1.272477e-10, 1.276794e-10, 1.267977e-10, 1.277877e-10, 
    1.240912e-10, 1.260218e-10, 1.230039e-10, 1.239089e-10, 1.245398e-10, 
    1.242629e-10, 1.257044e-10, 1.260453e-10, 1.274352e-10, 1.267158e-10, 
    1.310278e-10, 1.291115e-10, 1.344628e-10, 1.329568e-10, 1.230137e-10, 
    1.234721e-10, 1.250741e-10, 1.243107e-10, 1.265002e-10, 1.270419e-10, 
    1.274832e-10, 1.280483e-10, 1.281094e-10, 1.284449e-10, 1.278954e-10, 
    1.284231e-10, 1.26432e-10, 1.2732e-10, 1.248906e-10, 1.254798e-10, 
    1.252085e-10, 1.249114e-10, 1.258297e-10, 1.268115e-10, 1.268326e-10, 
    1.271483e-10, 1.280396e-10, 1.265091e-10, 1.312761e-10, 1.28322e-10, 
    1.23973e-10, 1.248601e-10, 1.249871e-10, 1.246429e-10, 1.269876e-10, 
    1.261356e-10, 1.284367e-10, 1.278128e-10, 1.288358e-10, 1.28327e-10, 
    1.282522e-10, 1.276003e-10, 1.271952e-10, 1.261746e-10, 1.253471e-10, 
    1.246928e-10, 1.248448e-10, 1.25564e-10, 1.268717e-10, 1.281149e-10, 
    1.278421e-10, 1.287579e-10, 1.263408e-10, 1.273516e-10, 1.269605e-10, 
    1.279816e-10, 1.257493e-10, 1.276489e-10, 1.252659e-10, 1.25474e-10, 
    1.261187e-10, 1.274203e-10, 1.277092e-10, 1.280179e-10, 1.278274e-10, 
    1.26905e-10, 1.267542e-10, 1.26103e-10, 1.259235e-10, 1.254287e-10, 
    1.250197e-10, 1.253933e-10, 1.257863e-10, 1.269054e-10, 1.279181e-10, 
    1.290266e-10, 1.292986e-10, 1.306008e-10, 1.295402e-10, 1.312926e-10, 
    1.29802e-10, 1.323876e-10, 1.277595e-10, 1.297583e-10, 1.261481e-10, 
    1.265347e-10, 1.272353e-10, 1.288494e-10, 1.279768e-10, 1.289976e-10, 
    1.267483e-10, 1.255888e-10, 1.252897e-10, 1.247325e-10, 1.253025e-10, 
    1.252561e-10, 1.258026e-10, 1.256268e-10, 1.269427e-10, 1.262351e-10, 
    1.282503e-10, 1.289895e-10, 1.310883e-10, 1.323829e-10, 1.337072e-10, 
    1.342938e-10, 1.344726e-10, 1.345473e-10,
  1.315636e-10, 1.327923e-10, 1.325529e-10, 1.335477e-10, 1.329953e-10, 
    1.336475e-10, 1.318122e-10, 1.328412e-10, 1.321838e-10, 1.316739e-10, 
    1.354906e-10, 1.335922e-10, 1.374788e-10, 1.36256e-10, 1.393397e-10, 
    1.372882e-10, 1.397556e-10, 1.392803e-10, 1.407135e-10, 1.403021e-10, 
    1.421447e-10, 1.409037e-10, 1.431054e-10, 1.418478e-10, 1.420441e-10, 
    1.408629e-10, 1.33973e-10, 1.352534e-10, 1.338973e-10, 1.340794e-10, 
    1.339977e-10, 1.330067e-10, 1.32509e-10, 1.314699e-10, 1.316582e-10, 
    1.324215e-10, 1.341614e-10, 1.335693e-10, 1.350643e-10, 1.350304e-10, 
    1.367059e-10, 1.35949e-10, 1.387831e-10, 1.379741e-10, 1.403192e-10, 
    1.397273e-10, 1.402914e-10, 1.401202e-10, 1.402936e-10, 1.394261e-10, 
    1.397974e-10, 1.390354e-10, 1.360906e-10, 1.369523e-10, 1.343916e-10, 
    1.328655e-10, 1.318572e-10, 1.311444e-10, 1.312451e-10, 1.31437e-10, 
    1.32426e-10, 1.333597e-10, 1.340738e-10, 1.345527e-10, 1.350256e-10, 
    1.364627e-10, 1.372269e-10, 1.38947e-10, 1.386356e-10, 1.391633e-10, 
    1.396685e-10, 1.405191e-10, 1.403789e-10, 1.407543e-10, 1.391494e-10, 
    1.402149e-10, 1.384584e-10, 1.389376e-10, 1.351544e-10, 1.337289e-10, 
    1.331257e-10, 1.325989e-10, 1.313225e-10, 1.322032e-10, 1.318556e-10, 
    1.326834e-10, 1.33211e-10, 1.329499e-10, 1.345658e-10, 1.339363e-10, 
    1.372723e-10, 1.358295e-10, 1.396095e-10, 1.386995e-10, 1.398281e-10, 
    1.392515e-10, 1.402404e-10, 1.393503e-10, 1.408942e-10, 1.412318e-10, 
    1.410011e-10, 1.418884e-10, 1.39301e-10, 1.402914e-10, 1.329426e-10, 
    1.329851e-10, 1.331835e-10, 1.323128e-10, 1.322596e-10, 1.314648e-10, 
    1.321719e-10, 1.324737e-10, 1.332416e-10, 1.33697e-10, 1.341307e-10, 
    1.350872e-10, 1.361602e-10, 1.376687e-10, 1.387584e-10, 1.394916e-10, 
    1.390417e-10, 1.394389e-10, 1.38995e-10, 1.387872e-10, 1.411052e-10, 
    1.398009e-10, 1.417606e-10, 1.416517e-10, 1.407633e-10, 1.41664e-10, 
    1.33015e-10, 1.327702e-10, 1.319222e-10, 1.325856e-10, 1.313784e-10, 
    1.320533e-10, 1.324423e-10, 1.339494e-10, 1.342818e-10, 1.345905e-10, 
    1.352014e-10, 1.359877e-10, 1.373734e-10, 1.385858e-10, 1.396979e-10, 
    1.396162e-10, 1.39645e-10, 1.398941e-10, 1.392775e-10, 1.399955e-10, 
    1.401162e-10, 1.398007e-10, 1.416372e-10, 1.411111e-10, 1.416494e-10, 
    1.413067e-10, 1.328497e-10, 1.33262e-10, 1.330391e-10, 1.334584e-10, 
    1.33163e-10, 1.344795e-10, 1.348757e-10, 1.367385e-10, 1.359722e-10, 
    1.371929e-10, 1.360959e-10, 1.362899e-10, 1.372329e-10, 1.36155e-10, 
    1.385188e-10, 1.369137e-10, 1.399038e-10, 1.382917e-10, 1.400052e-10, 
    1.396931e-10, 1.4021e-10, 1.406739e-10, 1.412588e-10, 1.423418e-10, 
    1.420906e-10, 1.42999e-10, 1.338779e-10, 1.344151e-10, 1.343678e-10, 
    1.349312e-10, 1.353488e-10, 1.362563e-10, 1.377193e-10, 1.371681e-10, 
    1.38181e-10, 1.383849e-10, 1.368464e-10, 1.377899e-10, 1.347754e-10, 
    1.352598e-10, 1.349712e-10, 1.339203e-10, 1.372951e-10, 1.355571e-10, 
    1.387764e-10, 1.378274e-10, 1.406077e-10, 1.39221e-10, 1.419524e-10, 
    1.431296e-10, 1.442426e-10, 1.455498e-10, 1.347088e-10, 1.343432e-10, 
    1.349983e-10, 1.359077e-10, 1.367545e-10, 1.378852e-10, 1.380012e-10, 
    1.382137e-10, 1.38765e-10, 1.392296e-10, 1.382809e-10, 1.393462e-10, 
    1.353724e-10, 1.374465e-10, 1.342052e-10, 1.351765e-10, 1.35854e-10, 
    1.355565e-10, 1.371052e-10, 1.374717e-10, 1.389669e-10, 1.381928e-10, 
    1.428385e-10, 1.407721e-10, 1.465497e-10, 1.449214e-10, 1.342156e-10, 
    1.347076e-10, 1.36428e-10, 1.356078e-10, 1.379608e-10, 1.385436e-10, 
    1.390184e-10, 1.396268e-10, 1.396926e-10, 1.400539e-10, 1.394621e-10, 
    1.400304e-10, 1.378876e-10, 1.388428e-10, 1.362306e-10, 1.368638e-10, 
    1.365723e-10, 1.36253e-10, 1.372399e-10, 1.382958e-10, 1.383184e-10, 
    1.386581e-10, 1.396178e-10, 1.379704e-10, 1.431066e-10, 1.399218e-10, 
    1.352452e-10, 1.36198e-10, 1.363344e-10, 1.359646e-10, 1.384851e-10, 
    1.375688e-10, 1.40045e-10, 1.393732e-10, 1.404749e-10, 1.399269e-10, 
    1.398463e-10, 1.391445e-10, 1.387085e-10, 1.376107e-10, 1.367212e-10, 
    1.360182e-10, 1.361815e-10, 1.369544e-10, 1.383606e-10, 1.396985e-10, 
    1.394048e-10, 1.40391e-10, 1.377894e-10, 1.388769e-10, 1.38456e-10, 
    1.39555e-10, 1.371535e-10, 1.391971e-10, 1.36634e-10, 1.368576e-10, 
    1.375506e-10, 1.389509e-10, 1.392617e-10, 1.395941e-10, 1.39389e-10, 
    1.383964e-10, 1.382341e-10, 1.375337e-10, 1.373407e-10, 1.368089e-10, 
    1.363694e-10, 1.367709e-10, 1.371933e-10, 1.383968e-10, 1.394866e-10, 
    1.406805e-10, 1.409736e-10, 1.423779e-10, 1.412342e-10, 1.431245e-10, 
    1.415165e-10, 1.443067e-10, 1.39316e-10, 1.414693e-10, 1.375822e-10, 
    1.379979e-10, 1.387518e-10, 1.404897e-10, 1.395498e-10, 1.406493e-10, 
    1.382278e-10, 1.369811e-10, 1.366596e-10, 1.360609e-10, 1.366733e-10, 
    1.366234e-10, 1.372107e-10, 1.370218e-10, 1.384368e-10, 1.376757e-10, 
    1.398443e-10, 1.406406e-10, 1.429036e-10, 1.443014e-10, 1.457324e-10, 
    1.463669e-10, 1.465603e-10, 1.466412e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24575.68, 24595.97, 24591.99, 24608.59, 24599.35, 24610.27, 24579.76, 
    24596.79, 24585.88, 24577.49, 24641.53, 24609.34, 24676.01, 24654.69, 
    24708.69, 24672.66, 24716.09, 24707.63, 24733.32, 24725.89, 24759.5, 
    24736.77, 24777.39, 24754.02, 24757.63, 24736.03, 24615.75, 24637.48, 
    24614.47, 24617.54, 24616.16, 24599.54, 24591.27, 24574.14, 24577.23, 
    24589.82, 24618.93, 24608.95, 24634.26, 24633.68, 24662.49, 24649.39, 
    24698.84, 24684.68, 24726.2, 24715.59, 24725.7, 24722.62, 24725.74, 
    24710.22, 24716.84, 24703.29, 24651.83, 24666.78, 24622.83, 24597.19, 
    24580.5, 24568.8, 24570.45, 24573.6, 24589.89, 24605.44, 24617.45, 
    24625.56, 24633.6, 24658.27, 24671.59, 24701.73, 24696.25, 24705.56, 
    24714.54, 24729.81, 24727.28, 24734.06, 24705.31, 24724.32, 24693.14, 
    24701.57, 24635.79, 24611.63, 24601.53, 24592.76, 24571.72, 24586.21, 
    24580.48, 24594.16, 24602.95, 24598.59, 24625.79, 24615.13, 24672.38, 
    24647.34, 24713.48, 24697.37, 24717.39, 24707.12, 24724.78, 24708.87, 
    24736.6, 24742.74, 24738.54, 24754.76, 24708, 24725.7, 24598.47, 
    24599.18, 24602.49, 24588.02, 24587.14, 24574.05, 24585.69, 24590.68, 
    24603.46, 24611.1, 24618.41, 24634.65, 24653.04, 24679.35, 24698.41, 
    24711.38, 24703.41, 24710.45, 24702.58, 24698.92, 24740.43, 24716.9, 
    24752.41, 24750.41, 24734.22, 24750.64, 24599.68, 24595.6, 24581.57, 
    24592.54, 24572.64, 24583.73, 24590.16, 24615.35, 24620.97, 24626.21, 
    24636.59, 24650.06, 24674.15, 24695.38, 24715.06, 24713.6, 24714.12, 
    24718.57, 24707.58, 24720.38, 24722.55, 24716.9, 24750.15, 24740.54, 
    24750.37, 24744.1, 24596.93, 24603.8, 24600.08, 24607.09, 24602.15, 
    24624.32, 24631.05, 24663.06, 24649.79, 24670.99, 24651.92, 24655.28, 
    24671.69, 24652.95, 24694.2, 24666.11, 24718.74, 24690.22, 24720.56, 
    24714.97, 24724.23, 24732.61, 24743.23, 24763.14, 24758.49, 24775.4, 
    24614.14, 24623.23, 24622.42, 24631.99, 24639.1, 24654.69, 24680.24, 
    24670.55, 24688.29, 24691.85, 24664.94, 24681.48, 24629.35, 24637.59, 
    24632.67, 24614.86, 24672.78, 24642.67, 24698.73, 24682.13, 24731.41, 
    24706.58, 24755.94, 24777.85, 24798.95, 24824.03, 24628.22, 24622.01, 
    24633.13, 24648.68, 24663.34, 24683.14, 24685.15, 24688.86, 24698.53, 
    24706.73, 24690.04, 24708.8, 24639.51, 24675.44, 24619.67, 24636.17, 
    24647.76, 24642.66, 24669.45, 24675.88, 24702.09, 24688.49, 24772.4, 
    24734.38, 24843.32, 24812, 24619.85, 24628.2, 24657.67, 24643.54, 
    24684.45, 24694.63, 24703, 24713.79, 24714.96, 24721.43, 24710.86, 
    24721.01, 24683.18, 24699.9, 24654.25, 24665.24, 24660.17, 24654.64, 
    24671.81, 24690.3, 24690.69, 24696.65, 24713.64, 24684.62, 24777.42, 
    24719.07, 24637.34, 24653.69, 24656.04, 24649.66, 24693.61, 24677.59, 
    24721.27, 24709.28, 24729.01, 24719.15, 24717.71, 24705.22, 24697.53, 
    24678.33, 24662.76, 24650.58, 24653.4, 24666.82, 24691.43, 24715.07, 
    24709.84, 24727.49, 24681.47, 24700.5, 24693.1, 24712.51, 24670.3, 
    24706.16, 24661.24, 24665.13, 24677.27, 24701.8, 24707.3, 24713.21, 
    24709.56, 24692.05, 24689.22, 24676.97, 24673.58, 24664.28, 24656.65, 
    24663.62, 24670.99, 24692.06, 24711.3, 24732.72, 24738.04, 24763.82, 
    24742.78, 24777.76, 24747.94, 24800.18, 24708.27, 24747.08, 24677.82, 
    24685.1, 24698.29, 24729.28, 24712.42, 24732.16, 24689.11, 24667.29, 
    24661.68, 24651.32, 24661.92, 24661.05, 24671.3, 24668, 24692.76, 
    24679.47, 24717.68, 24732, 24773.61, 24800.08, 24827.53, 24839.77, 
    24843.53, 24845.1 ;

 GC_ICE1 =
  17685.98, 17718.49, 17712.12, 17738.7, 17723.9, 17741.39, 17692.52, 
    17719.79, 17702.33, 17688.88, 17791.44, 17739.9, 17846.59, 17812.49, 
    17898.77, 17841.23, 17910.59, 17897.08, 17938.08, 17926.22, 17979.83, 
    17943.58, 18008.37, 17971.09, 17976.86, 17942.39, 17750.16, 17784.96, 
    17748.12, 17753.04, 17750.83, 17724.21, 17710.95, 17683.51, 17688.47, 
    17708.63, 17755.26, 17739.28, 17779.79, 17778.87, 17824.97, 17804.01, 
    17883.06, 17860.46, 17926.72, 17909.78, 17925.92, 17921, 17925.98, 
    17901.21, 17911.78, 17890.16, 17807.92, 17831.83, 17761.5, 17720.44, 
    17693.71, 17674.96, 17677.6, 17682.65, 17708.75, 17733.66, 17752.89, 
    17765.88, 17778.74, 17818.22, 17839.52, 17887.67, 17878.92, 17893.78, 
    17908.1, 17932.47, 17928.43, 17939.26, 17893.38, 17923.72, 17873.96, 
    17887.41, 17782.26, 17743.57, 17727.39, 17713.34, 17679.63, 17702.84, 
    17693.66, 17715.59, 17729.67, 17722.69, 17766.24, 17749.17, 17840.79, 
    17800.73, 17906.42, 17880.71, 17912.65, 17896.27, 17924.45, 17899.06, 
    17943.3, 17953.1, 17946.4, 17972.28, 17897.67, 17925.92, 17722.49, 
    17723.63, 17728.94, 17705.75, 17704.34, 17683.38, 17702.01, 17710.01, 
    17730.49, 17742.72, 17754.43, 17780.42, 17809.84, 17851.93, 17882.37, 
    17903.07, 17890.34, 17901.58, 17889.02, 17883.17, 17949.42, 17911.88, 
    17968.53, 17965.34, 17939.52, 17965.7, 17724.43, 17717.9, 17695.42, 
    17712.98, 17681.1, 17698.88, 17709.18, 17749.53, 17758.52, 17766.91, 
    17783.53, 17805.08, 17843.62, 17877.52, 17908.94, 17906.62, 17907.43, 
    17914.54, 17897, 17917.43, 17920.89, 17911.87, 17964.92, 17949.59, 
    17965.28, 17955.28, 17720.02, 17731.04, 17725.07, 17736.3, 17728.39, 
    17763.89, 17774.67, 17825.88, 17804.65, 17838.56, 17808.06, 17813.43, 
    17839.69, 17809.7, 17875.65, 17830.76, 17914.81, 17869.3, 17917.71, 
    17908.8, 17923.58, 17936.94, 17953.88, 17985.64, 17978.23, 18005.19, 
    17747.59, 17762.14, 17760.85, 17776.17, 17787.55, 17812.49, 17853.36, 
    17837.87, 17866.21, 17871.9, 17828.88, 17855.35, 17771.95, 17785.12, 
    17777.26, 17748.74, 17841.43, 17793.25, 17882.87, 17856.38, 17935.03, 
    17895.41, 17974.16, 18009.1, 18042.74, 18082.67, 17770.14, 17760.19, 
    17778, 17802.88, 17826.32, 17857.99, 17861.21, 17867.12, 17882.55, 
    17895.65, 17869, 17898.95, 17788.2, 17845.68, 17756.44, 17782.85, 
    17801.4, 17793.23, 17836.11, 17846.38, 17888.23, 17866.54, 18000.4, 
    17939.77, 18113.33, 18063.54, 17756.72, 17770.1, 17817.25, 17794.64, 
    17860.09, 17876.34, 17889.68, 17906.92, 17908.79, 17919.11, 17902.24, 
    17918.43, 17858.05, 17884.74, 17811.78, 17829.36, 17821.25, 17812.4, 
    17839.88, 17869.42, 17870.04, 17879.55, 17906.67, 17860.35, 18008.42, 
    17915.34, 17784.72, 17810.89, 17814.65, 17804.44, 17874.71, 17849.12, 
    17918.85, 17899.71, 17931.2, 17915.47, 17913.17, 17893.24, 17880.96, 
    17850.3, 17825.39, 17805.92, 17810.43, 17831.89, 17871.22, 17908.96, 
    17900.61, 17928.78, 17855.33, 17885.7, 17873.89, 17904.88, 17837.46, 
    17894.74, 17822.96, 17829.19, 17848.61, 17887.78, 17896.56, 17905.99, 
    17900.16, 17872.22, 17867.69, 17848.13, 17842.71, 17827.83, 17815.62, 
    17826.78, 17838.57, 17872.23, 17902.93, 17937.13, 17945.6, 17986.72, 
    17953.17, 18008.95, 17961.4, 18044.71, 17898.1, 17960.02, 17849.49, 
    17861.12, 17882.18, 17931.63, 17904.73, 17936.23, 17867.52, 17832.64, 
    17823.68, 17807.1, 17824.06, 17822.67, 17839.06, 17833.77, 17873.35, 
    17852.13, 17913.12, 17935.98, 18002.34, 18044.54, 18088.24, 18107.7, 
    18113.66, 18116.16 ;

 GC_LIQ1 =
  5232.713, 5234.742, 5234.344, 5236.006, 5235.081, 5236.174, 5233.121, 
    5234.824, 5233.733, 5232.894, 5239.315, 5236.081, 5242.794, 5240.642, 
    5246.144, 5242.456, 5246.906, 5246.036, 5248.679, 5247.914, 5251.38, 
    5249.034, 5253.229, 5250.814, 5251.188, 5248.958, 5236.723, 5238.906, 
    5236.595, 5236.903, 5236.764, 5235.1, 5234.272, 5232.56, 5232.869, 
    5234.127, 5237.042, 5236.042, 5238.581, 5238.522, 5241.43, 5240.108, 
    5245.132, 5243.676, 5247.946, 5246.854, 5247.894, 5247.578, 5247.898, 
    5246.302, 5246.982, 5245.59, 5240.354, 5241.863, 5237.432, 5234.864, 
    5233.195, 5232.028, 5232.192, 5232.506, 5234.134, 5235.69, 5236.893, 
    5237.706, 5238.514, 5241.004, 5242.348, 5245.429, 5244.865, 5245.822, 
    5246.746, 5248.317, 5248.057, 5248.755, 5245.797, 5247.752, 5244.546, 
    5245.412, 5238.736, 5236.311, 5235.298, 5234.421, 5232.319, 5233.766, 
    5233.193, 5234.561, 5235.441, 5235.005, 5237.729, 5236.66, 5242.428, 
    5239.9, 5246.638, 5244.981, 5247.039, 5245.983, 5247.8, 5246.163, 
    5249.017, 5249.65, 5249.217, 5250.892, 5246.073, 5247.895, 5234.993, 
    5235.063, 5235.395, 5233.947, 5233.859, 5232.552, 5233.714, 5234.213, 
    5235.492, 5236.257, 5236.989, 5238.62, 5240.475, 5243.131, 5245.087, 
    5246.421, 5245.601, 5246.325, 5245.516, 5245.139, 5249.412, 5246.989, 
    5250.649, 5250.442, 5248.772, 5250.466, 5235.113, 5234.706, 5233.302, 
    5234.398, 5232.41, 5233.518, 5234.161, 5236.683, 5237.246, 5237.771, 
    5238.816, 5240.175, 5242.607, 5244.775, 5246.8, 5246.65, 5246.703, 
    5247.16, 5246.03, 5247.347, 5247.57, 5246.988, 5250.415, 5249.423, 
    5250.438, 5249.791, 5234.838, 5235.526, 5235.154, 5235.855, 5235.36, 
    5237.582, 5238.258, 5241.487, 5240.148, 5242.288, 5240.363, 5240.701, 
    5242.358, 5240.466, 5244.655, 5241.795, 5247.178, 5244.246, 5247.365, 
    5246.791, 5247.744, 5248.605, 5249.701, 5251.757, 5251.277, 5253.023, 
    5236.562, 5237.472, 5237.392, 5238.353, 5239.07, 5240.643, 5243.222, 
    5242.244, 5244.047, 5244.414, 5241.676, 5243.348, 5238.086, 5238.917, 
    5238.421, 5236.633, 5242.468, 5239.429, 5245.12, 5243.415, 5248.482, 
    5245.928, 5251.014, 5253.277, 5255.458, 5258.077, 5237.973, 5237.35, 
    5238.467, 5240.036, 5241.515, 5243.518, 5243.725, 5244.105, 5245.099, 
    5245.943, 5244.227, 5246.156, 5239.111, 5242.737, 5237.116, 5238.773, 
    5239.943, 5239.428, 5242.132, 5242.781, 5245.465, 5244.068, 5252.713, 
    5248.789, 5260.122, 5256.811, 5237.133, 5237.97, 5240.942, 5239.517, 
    5243.653, 5244.699, 5245.559, 5246.669, 5246.79, 5247.455, 5246.368, 
    5247.412, 5243.522, 5245.24, 5240.598, 5241.707, 5241.195, 5240.637, 
    5242.371, 5244.253, 5244.294, 5244.906, 5246.653, 5243.67, 5253.232, 
    5247.212, 5238.892, 5240.542, 5240.779, 5240.135, 5244.594, 5242.954, 
    5247.438, 5246.205, 5248.235, 5247.221, 5247.072, 5245.788, 5244.997, 
    5243.028, 5241.457, 5240.228, 5240.512, 5241.867, 5244.37, 5246.801, 
    5246.263, 5248.079, 5243.347, 5245.302, 5244.542, 5246.538, 5242.218, 
    5245.884, 5241.303, 5241.696, 5242.921, 5245.437, 5246.001, 5246.609, 
    5246.234, 5244.434, 5244.143, 5242.892, 5242.549, 5241.61, 5240.84, 
    5241.543, 5242.288, 5244.435, 5246.413, 5248.618, 5249.165, 5251.827, 
    5249.655, 5253.268, 5250.188, 5255.586, 5246.101, 5250.098, 5242.978, 
    5243.719, 5245.076, 5248.263, 5246.528, 5248.56, 5244.131, 5241.914, 
    5241.348, 5240.302, 5241.372, 5241.285, 5242.319, 5241.985, 5244.507, 
    5243.144, 5247.069, 5248.543, 5252.839, 5255.575, 5258.447, 5259.745, 
    5260.144, 5260.311 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.728482e-09, 8.766966e-09, 8.759486e-09, 8.790525e-09, 8.773307e-09, 
    8.793632e-09, 8.736285e-09, 8.768493e-09, 8.747932e-09, 8.731948e-09, 
    8.850763e-09, 8.79191e-09, 8.911909e-09, 8.87437e-09, 8.968676e-09, 
    8.906067e-09, 8.981302e-09, 8.966873e-09, 9.010307e-09, 8.997864e-09, 
    9.053418e-09, 9.016051e-09, 9.082221e-09, 9.044496e-09, 9.050396e-09, 
    9.014817e-09, 8.803755e-09, 8.843435e-09, 8.801404e-09, 8.807063e-09, 
    8.804523e-09, 8.773662e-09, 8.758109e-09, 8.725542e-09, 8.731455e-09, 
    8.755375e-09, 8.809606e-09, 8.791198e-09, 8.837596e-09, 8.836548e-09, 
    8.888205e-09, 8.864914e-09, 8.951743e-09, 8.927064e-09, 8.998383e-09, 
    8.980447e-09, 8.99754e-09, 8.992357e-09, 8.997608e-09, 8.971302e-09, 
    8.982572e-09, 8.959426e-09, 8.869276e-09, 8.895769e-09, 8.816755e-09, 
    8.769247e-09, 8.737697e-09, 8.715308e-09, 8.718474e-09, 8.724507e-09, 
    8.755515e-09, 8.784671e-09, 8.80689e-09, 8.821753e-09, 8.836398e-09, 
    8.880725e-09, 8.90419e-09, 8.956733e-09, 8.947252e-09, 8.963315e-09, 
    8.978662e-09, 9.004427e-09, 9.000187e-09, 9.011539e-09, 8.962892e-09, 
    8.995221e-09, 8.941852e-09, 8.956448e-09, 8.840373e-09, 8.796165e-09, 
    8.777369e-09, 8.760923e-09, 8.720908e-09, 8.748541e-09, 8.737647e-09, 
    8.763565e-09, 8.780034e-09, 8.771889e-09, 8.822159e-09, 8.802615e-09, 
    8.905581e-09, 8.861229e-09, 8.976872e-09, 8.949198e-09, 8.983505e-09, 
    8.965999e-09, 8.995995e-09, 8.969e-09, 9.015764e-09, 9.025946e-09, 
    9.018988e-09, 9.045721e-09, 8.967502e-09, 8.99754e-09, 8.77166e-09, 
    8.772989e-09, 8.779177e-09, 8.751972e-09, 8.750308e-09, 8.72538e-09, 
    8.747562e-09, 8.757008e-09, 8.780988e-09, 8.795173e-09, 8.808657e-09, 
    8.838304e-09, 8.871416e-09, 8.917722e-09, 8.950992e-09, 8.973294e-09, 
    8.959619e-09, 8.971692e-09, 8.958196e-09, 8.95187e-09, 9.022131e-09, 
    8.982678e-09, 9.041876e-09, 9.0386e-09, 9.011808e-09, 9.03897e-09, 
    8.773921e-09, 8.766277e-09, 8.739736e-09, 8.760507e-09, 8.722665e-09, 
    8.743846e-09, 8.756025e-09, 8.803021e-09, 8.813349e-09, 8.822924e-09, 
    8.841836e-09, 8.866106e-09, 8.908684e-09, 8.945732e-09, 8.979556e-09, 
    8.977077e-09, 8.97795e-09, 8.985505e-09, 8.966789e-09, 8.988578e-09, 
    8.992234e-09, 8.982673e-09, 9.038161e-09, 9.022309e-09, 9.038531e-09, 
    9.028209e-09, 8.768763e-09, 8.781624e-09, 8.774674e-09, 8.787744e-09, 
    8.778536e-09, 8.819479e-09, 8.831756e-09, 8.889203e-09, 8.865628e-09, 
    8.90315e-09, 8.86944e-09, 8.875412e-09, 8.904371e-09, 8.871262e-09, 
    8.943688e-09, 8.894583e-09, 8.985799e-09, 8.936757e-09, 8.988872e-09, 
    8.979409e-09, 8.995078e-09, 9.009109e-09, 9.026764e-09, 9.059338e-09, 
    9.051796e-09, 9.079039e-09, 8.800801e-09, 8.817485e-09, 8.816016e-09, 
    8.833477e-09, 8.84639e-09, 8.87438e-09, 8.919273e-09, 8.902392e-09, 
    8.933386e-09, 8.939607e-09, 8.892521e-09, 8.92143e-09, 8.828651e-09, 
    8.843639e-09, 8.834716e-09, 8.802116e-09, 8.90628e-09, 8.852821e-09, 
    8.951542e-09, 8.922579e-09, 9.007108e-09, 8.965069e-09, 9.047643e-09, 
    9.082942e-09, 9.116171e-09, 9.154999e-09, 8.826591e-09, 8.815254e-09, 
    8.835554e-09, 8.863637e-09, 8.889699e-09, 8.924346e-09, 8.927891e-09, 
    8.934381e-09, 8.951195e-09, 8.965332e-09, 8.936433e-09, 8.968876e-09, 
    8.847112e-09, 8.910921e-09, 8.810968e-09, 8.841063e-09, 8.861982e-09, 
    8.852806e-09, 8.900463e-09, 8.911694e-09, 8.957338e-09, 8.933744e-09, 
    9.074228e-09, 9.012071e-09, 9.184567e-09, 9.136357e-09, 8.811294e-09, 
    8.826553e-09, 8.879659e-09, 8.854391e-09, 8.926659e-09, 8.944448e-09, 
    8.958911e-09, 8.977397e-09, 8.979393e-09, 8.990346e-09, 8.972398e-09, 
    8.989638e-09, 8.924419e-09, 8.953564e-09, 8.87359e-09, 8.893053e-09, 
    8.8841e-09, 8.874278e-09, 8.904593e-09, 8.936888e-09, 8.93758e-09, 
    8.947935e-09, 8.977112e-09, 8.926953e-09, 9.082248e-09, 8.986334e-09, 
    8.843192e-09, 8.872582e-09, 8.876782e-09, 8.865396e-09, 8.942664e-09, 
    8.914666e-09, 8.99008e-09, 8.969698e-09, 9.003094e-09, 8.986499e-09, 
    8.984057e-09, 8.962743e-09, 8.949474e-09, 8.91595e-09, 8.888675e-09, 
    8.867048e-09, 8.872076e-09, 8.895833e-09, 8.938863e-09, 8.979574e-09, 
    8.970655e-09, 9.000556e-09, 8.921419e-09, 8.954601e-09, 8.941775e-09, 
    8.975218e-09, 8.901943e-09, 8.964334e-09, 8.885995e-09, 8.892864e-09, 
    8.914111e-09, 8.956849e-09, 8.966309e-09, 8.976405e-09, 8.970176e-09, 
    8.939956e-09, 8.935006e-09, 8.913595e-09, 8.907683e-09, 8.891369e-09, 
    8.877862e-09, 8.890201e-09, 8.903161e-09, 8.93997e-09, 8.973141e-09, 
    9.009308e-09, 9.01816e-09, 9.060416e-09, 9.026015e-09, 9.082782e-09, 
    9.034516e-09, 9.118071e-09, 8.967953e-09, 9.0331e-09, 8.915078e-09, 
    8.927793e-09, 8.950789e-09, 9.003536e-09, 8.975061e-09, 9.008363e-09, 
    8.934812e-09, 8.896652e-09, 8.886782e-09, 8.868362e-09, 8.887203e-09, 
    8.885671e-09, 8.903699e-09, 8.897906e-09, 8.941192e-09, 8.91794e-09, 
    8.983995e-09, 9.008101e-09, 9.076182e-09, 9.11792e-09, 9.160412e-09, 
    9.17917e-09, 9.18488e-09, 9.187267e-09 ;

 H2OCAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  6.240021, 6.269336, 6.263629, 6.287323, 6.274172, 6.289697, 6.245955, 
    6.270503, 6.254825, 6.242654, 6.333463, 6.288381, 6.380479, 6.351581, 
    6.424317, 6.375979, 6.434089, 6.422915, 6.456569, 6.446917, 6.490081, 
    6.461026, 6.512516, 6.483133, 6.487726, 6.46007, 6.297435, 6.327841, 
    6.295637, 6.299966, 6.298023, 6.274445, 6.262585, 6.237781, 6.242279, 
    6.260498, 6.301914, 6.287834, 6.323347, 6.322544, 6.36222, 6.344313, 
    6.411217, 6.392159, 6.44732, 6.433422, 6.446667, 6.442649, 6.44672, 
    6.426344, 6.43507, 6.417155, 6.347665, 6.368043, 6.307384, 6.271082, 
    6.247032, 6.230001, 6.232408, 6.236996, 6.260604, 6.282847, 6.299831, 
    6.311207, 6.322428, 6.356475, 6.374532, 6.415077, 6.407745, 6.420166, 
    6.43204, 6.452009, 6.44872, 6.457527, 6.419836, 6.444872, 6.403573, 
    6.414853, 6.325493, 6.29163, 6.27728, 6.264727, 6.234258, 6.25529, 
    6.246994, 6.266739, 6.279306, 6.273088, 6.311519, 6.296562, 6.375603, 
    6.341485, 6.430655, 6.40925, 6.435791, 6.422239, 6.44547, 6.42456, 
    6.460805, 6.468715, 6.463309, 6.484084, 6.423402, 6.446668, 6.272914, 
    6.273929, 6.278652, 6.257905, 6.256636, 6.237659, 6.254542, 6.261741, 
    6.280034, 6.290872, 6.301184, 6.323892, 6.349313, 6.384957, 6.410636, 
    6.427884, 6.417304, 6.426644, 6.416203, 6.411313, 6.465751, 6.435152, 
    6.481093, 6.478546, 6.457736, 6.478833, 6.27464, 6.268807, 6.248583, 
    6.264407, 6.235593, 6.251713, 6.260994, 6.296877, 6.304774, 6.312106, 
    6.326599, 6.345229, 6.37799, 6.406574, 6.432731, 6.430812, 6.431488, 
    6.43734, 6.422851, 6.439721, 6.442555, 6.435146, 6.478204, 6.465886, 
    6.478491, 6.470469, 6.270702, 6.280521, 6.275214, 6.285196, 6.278164, 
    6.309472, 6.318877, 6.362993, 6.344862, 6.373728, 6.34779, 6.352382, 
    6.374676, 6.349189, 6.404998, 6.367135, 6.437568, 6.399649, 6.439949, 
    6.432618, 6.444757, 6.455641, 6.469347, 6.494684, 6.488811, 6.510031, 
    6.295174, 6.307942, 6.306815, 6.32019, 6.330093, 6.351586, 6.386152, 
    6.37314, 6.397037, 6.401841, 6.36554, 6.387816, 6.316494, 6.327987, 
    6.321141, 6.296182, 6.37614, 6.335032, 6.411061, 6.3887, 6.454089, 
    6.421524, 6.48558, 6.513083, 6.539016, 6.56941, 6.314914, 6.306231, 
    6.321781, 6.343337, 6.363369, 6.390063, 6.392797, 6.397807, 6.410792, 
    6.421723, 6.399394, 6.424465, 6.330659, 6.379714, 6.302953, 6.326013, 
    6.342064, 6.335017, 6.371653, 6.380307, 6.415544, 6.397313, 6.50629, 
    6.457944, 6.592597, 6.55481, 6.3032, 6.314883, 6.355649, 6.336233, 
    6.391846, 6.40558, 6.416756, 6.431062, 6.432606, 6.441092, 6.42719, 
    6.440542, 6.39012, 6.412623, 6.350978, 6.365951, 6.35906, 6.351507, 
    6.374834, 6.399745, 6.400274, 6.408276, 6.43086, 6.392072, 6.512553, 
    6.437999, 6.327638, 6.35021, 6.353434, 6.344682, 6.404202, 6.382599, 
    6.440885, 6.425101, 6.450973, 6.438109, 6.436218, 6.419721, 6.409463, 
    6.383589, 6.362582, 6.345951, 6.349815, 6.368092, 6.40127, 6.432747, 
    6.425845, 6.449005, 6.387804, 6.413427, 6.403518, 6.429374, 6.372795, 
    6.420968, 6.360518, 6.365803, 6.38217, 6.41517, 6.422478, 6.430295, 
    6.42547, 6.402113, 6.398289, 6.381772, 6.377217, 6.364652, 6.354262, 
    6.363755, 6.373735, 6.402121, 6.427768, 6.455796, 6.462665, 6.495533, 
    6.468775, 6.51297, 6.475393, 6.540516, 6.42376, 6.474282, 6.382915, 
    6.39272, 6.410483, 6.451323, 6.429252, 6.455067, 6.398139, 6.368725, 
    6.361123, 6.346961, 6.361447, 6.360268, 6.374146, 6.369684, 6.403065, 
    6.385121, 6.436172, 6.454862, 6.507807, 6.540389, 6.573645, 6.588358, 
    6.59284, 6.594715,
  3.950678, 3.97015, 3.966359, 3.981968, 3.973362, 3.983499, 3.954619, 
    3.970926, 3.96051, 3.952426, 4.011738, 3.98265, 4.042078, 4.023426, 
    4.070379, 4.039175, 4.076689, 4.069473, 4.091205, 4.084971, 4.112855, 
    4.094084, 4.127348, 4.108365, 4.111333, 4.093466, 3.988489, 4.008111, 
    3.987329, 3.990123, 3.988868, 3.973544, 3.965667, 3.94919, 3.952177, 
    3.964279, 3.991379, 3.982296, 4.005206, 4.004688, 4.030292, 4.018734, 
    4.06192, 4.049615, 4.085231, 4.076257, 4.08481, 4.082215, 4.084844, 
    4.071686, 4.077321, 4.065753, 4.020898, 4.03405, 3.994908, 3.971312, 
    3.955334, 3.944023, 3.945621, 3.948669, 3.96435, 3.979079, 3.990034, 
    3.997374, 4.004613, 4.026587, 4.038239, 4.064413, 4.059678, 4.067698, 
    4.075365, 4.08826, 4.086135, 4.091824, 4.067484, 4.083652, 4.056983, 
    4.064267, 4.006597, 3.984745, 3.97543, 3.967088, 3.94685, 3.96082, 
    3.95531, 3.968424, 3.976774, 3.972642, 3.997575, 3.987926, 4.03893, 
    4.016911, 4.07447, 4.060649, 4.077786, 4.069035, 4.084038, 4.070534, 
    4.093941, 4.099051, 4.095559, 4.108977, 4.069787, 4.084812, 3.972527, 
    3.973201, 3.976339, 3.962557, 3.961714, 3.949109, 3.960323, 3.965105, 
    3.977257, 3.984256, 3.990908, 4.005558, 4.021962, 4.044968, 4.061544, 
    4.07268, 4.065848, 4.071879, 4.065138, 4.061981, 4.097137, 4.077374, 
    4.107046, 4.1054, 4.09196, 4.105586, 3.973674, 3.969798, 3.956365, 
    3.966875, 3.947737, 3.958444, 3.96461, 3.98813, 3.993223, 3.997954, 
    4.007304, 4.019326, 4.04047, 4.058922, 4.07581, 4.074571, 4.075007, 
    4.078787, 4.06943, 4.080324, 4.082156, 4.07737, 4.10518, 4.097223, 
    4.105365, 4.100183, 3.971057, 3.977579, 3.974055, 3.980595, 3.976015, 
    3.996256, 4.002324, 4.030792, 4.01909, 4.03772, 4.020978, 4.023942, 
    4.038334, 4.021881, 4.057906, 4.033466, 4.078934, 4.054454, 4.080471, 
    4.075737, 4.083576, 4.090606, 4.099458, 4.115827, 4.112032, 4.125742, 
    3.987031, 3.995268, 3.99454, 4.003169, 4.009559, 4.023428, 4.045738, 
    4.037339, 4.052764, 4.055866, 4.032433, 4.046813, 4.000785, 4.008202, 
    4.003783, 3.987682, 4.039277, 4.012747, 4.061819, 4.047383, 4.089603, 
    4.068575, 4.109945, 4.127716, 4.144472, 4.16412, 3.999766, 3.994164, 
    4.004196, 4.018106, 4.031033, 4.048263, 4.050027, 4.053262, 4.061645, 
    4.068702, 4.054287, 4.070472, 4.009929, 4.041584, 3.992049, 4.006928, 
    4.017284, 4.012737, 4.036379, 4.041965, 4.064714, 4.052942, 4.123328, 
    4.092095, 4.179109, 4.154682, 3.992208, 3.999745, 4.026051, 4.013521, 
    4.049413, 4.05828, 4.065495, 4.074733, 4.07573, 4.08121, 4.072232, 
    4.080854, 4.0483, 4.062827, 4.023036, 4.0327, 4.028251, 4.023377, 
    4.038432, 4.054514, 4.054854, 4.060021, 4.074609, 4.049559, 4.127378, 
    4.079218, 4.007975, 4.022542, 4.024621, 4.018972, 4.057391, 4.043445, 
    4.081076, 4.070883, 4.087591, 4.079284, 4.078063, 4.067409, 4.060787, 
    4.044084, 4.030525, 4.019791, 4.022285, 4.034081, 4.055499, 4.075822, 
    4.071365, 4.086319, 4.046804, 4.063347, 4.05695, 4.073643, 4.037117, 
    4.068221, 4.029191, 4.032603, 4.043168, 4.064473, 4.06919, 4.074238, 
    4.071122, 4.056043, 4.053574, 4.04291, 4.039971, 4.03186, 4.025155, 
    4.031282, 4.037724, 4.056047, 4.072607, 4.090707, 4.095142, 4.116378, 
    4.099092, 4.127648, 4.103371, 4.145446, 4.070022, 4.10265, 4.043648, 
    4.049978, 4.061447, 4.08782, 4.073564, 4.090237, 4.053476, 4.034491, 
    4.029583, 4.020443, 4.029792, 4.029031, 4.037988, 4.035108, 4.056656, 
    4.045072, 4.078033, 4.090104, 4.124305, 4.145361, 4.166854, 4.176367, 
    4.179265, 4.180477,
  3.294423, 3.312268, 3.308793, 3.323011, 3.315212, 3.324412, 3.298034, 
    3.312979, 3.303432, 3.296025, 3.350261, 3.323635, 3.378052, 3.360965, 
    3.40399, 3.375391, 3.409775, 3.40316, 3.423088, 3.417371, 3.44295, 
    3.425729, 3.456252, 3.43883, 3.441553, 3.425162, 3.328979, 3.34694, 
    3.327918, 3.330475, 3.329326, 3.315378, 3.308158, 3.293059, 3.295797, 
    3.306887, 3.331625, 3.323312, 3.344282, 3.343807, 3.367254, 3.356669, 
    3.396236, 3.384959, 3.417609, 3.40938, 3.417223, 3.414843, 3.417254, 
    3.405189, 3.410355, 3.39975, 3.358651, 3.370697, 3.334854, 3.313333, 
    3.298689, 3.288326, 3.28979, 3.292582, 3.306952, 3.320368, 3.330394, 
    3.337112, 3.343739, 3.363861, 3.374535, 3.39852, 3.394181, 3.401533, 
    3.408561, 3.420387, 3.418439, 3.423656, 3.401336, 3.416161, 3.391711, 
    3.398387, 3.345554, 3.325552, 3.317084, 3.309461, 3.290916, 3.303716, 
    3.298667, 3.310686, 3.318278, 3.314552, 3.337296, 3.328464, 3.375168, 
    3.354999, 3.407741, 3.395071, 3.410782, 3.402759, 3.416515, 3.404133, 
    3.425598, 3.430285, 3.427082, 3.439393, 3.403447, 3.417224, 3.314446, 
    3.315064, 3.317892, 3.305308, 3.304536, 3.292985, 3.303261, 3.307643, 
    3.318707, 3.325105, 3.331193, 3.344604, 3.359625, 3.3807, 3.395891, 
    3.4061, 3.399837, 3.405366, 3.399186, 3.396292, 3.428529, 3.410404, 
    3.43762, 3.43611, 3.42378, 3.43628, 3.315497, 3.311945, 3.299634, 
    3.309266, 3.291728, 3.301539, 3.307189, 3.328651, 3.333313, 3.337643, 
    3.346203, 3.357211, 3.376579, 3.393488, 3.40897, 3.407834, 3.408234, 
    3.4117, 3.403121, 3.413109, 3.414788, 3.410401, 3.435908, 3.428608, 
    3.436078, 3.431323, 3.313099, 3.318995, 3.315847, 3.321754, 3.317604, 
    3.336088, 3.341643, 3.367712, 3.356994, 3.374059, 3.358724, 3.361439, 
    3.374621, 3.359551, 3.392556, 3.370162, 3.411834, 3.389393, 3.413244, 
    3.408903, 3.416091, 3.422539, 3.430659, 3.445678, 3.442195, 3.454778, 
    3.327645, 3.335184, 3.334518, 3.342417, 3.348268, 3.360968, 3.381406, 
    3.37371, 3.387844, 3.390687, 3.369216, 3.382391, 3.340234, 3.347024, 
    3.342979, 3.32824, 3.375486, 3.351186, 3.396143, 3.382913, 3.421619, 
    3.402336, 3.44028, 3.456589, 3.471973, 3.490019, 3.339301, 3.334173, 
    3.343357, 3.356094, 3.367934, 3.383719, 3.385336, 3.3883, 3.395983, 
    3.402453, 3.38924, 3.404076, 3.348605, 3.377599, 3.332238, 3.345858, 
    3.355341, 3.351177, 3.372831, 3.377949, 3.398797, 3.388008, 3.452561, 
    3.423905, 3.503791, 3.481349, 3.332383, 3.339283, 3.36337, 3.351895, 
    3.384774, 3.3929, 3.399513, 3.407983, 3.408896, 3.413922, 3.40569, 
    3.413595, 3.383753, 3.397068, 3.360608, 3.36946, 3.365385, 3.360921, 
    3.374712, 3.389448, 3.38976, 3.394495, 3.407867, 3.384907, 3.456278, 
    3.412094, 3.346817, 3.360156, 3.36206, 3.356887, 3.392085, 3.379304, 
    3.413799, 3.404453, 3.419773, 3.412155, 3.411035, 3.401268, 3.395197, 
    3.37989, 3.367468, 3.357637, 3.359921, 3.370726, 3.39035, 3.408981, 
    3.404894, 3.418607, 3.382383, 3.397544, 3.39168, 3.406983, 3.373507, 
    3.402011, 3.366247, 3.369372, 3.379051, 3.398576, 3.4029, 3.407528, 
    3.404671, 3.390849, 3.388586, 3.378815, 3.376122, 3.368691, 3.362549, 
    3.368162, 3.374063, 3.390853, 3.406033, 3.422631, 3.4267, 3.446183, 
    3.430322, 3.456526, 3.434247, 3.472867, 3.403662, 3.433586, 3.379491, 
    3.385291, 3.395802, 3.419982, 3.406911, 3.422199, 3.388497, 3.371101, 
    3.366605, 3.358235, 3.366797, 3.3661, 3.374305, 3.371666, 3.391411, 
    3.380796, 3.411008, 3.422078, 3.453459, 3.47279, 3.492532, 3.501272, 
    3.503935, 3.505049,
  3.016801, 3.033729, 3.030432, 3.044127, 3.036524, 3.0455, 3.020226, 
    3.034404, 3.025347, 3.01832, 3.070836, 3.044739, 3.098105, 3.081336, 
    3.123583, 3.095493, 3.129268, 3.122767, 3.142358, 3.136736, 3.161451, 
    3.144955, 3.174125, 3.157528, 3.160121, 3.144397, 3.049975, 3.067579, 
    3.048935, 3.05144, 3.050315, 3.036681, 3.02983, 3.015508, 3.018104, 
    3.028623, 3.052567, 3.044422, 3.064974, 3.064509, 3.087507, 3.077122, 
    3.115964, 3.104887, 3.13697, 3.12888, 3.13659, 3.134251, 3.136621, 
    3.124761, 3.129839, 3.119416, 3.079066, 3.090886, 3.055732, 3.034739, 
    3.020847, 3.01102, 3.012408, 3.015055, 3.028685, 3.041538, 3.051361, 
    3.057945, 3.064442, 3.084176, 3.094652, 3.118208, 3.113945, 3.121168, 
    3.128076, 3.139702, 3.137785, 3.142916, 3.120975, 3.135545, 3.111519, 
    3.118078, 3.066219, 3.046617, 3.038321, 3.031066, 3.013475, 3.025616, 
    3.020826, 3.032228, 3.039491, 3.035897, 3.058125, 3.04947, 3.095274, 
    3.075483, 3.127269, 3.11482, 3.130258, 3.122373, 3.135894, 3.123723, 
    3.144826, 3.149391, 3.146285, 3.158064, 3.12305, 3.136591, 3.035797, 
    3.036383, 3.039113, 3.027126, 3.026393, 3.015437, 3.025183, 3.029341, 
    3.039912, 3.046179, 3.052144, 3.06529, 3.080021, 3.100705, 3.115626, 
    3.125657, 3.119503, 3.124936, 3.118863, 3.116019, 3.147709, 3.129887, 
    3.156376, 3.154938, 3.143038, 3.1551, 3.036794, 3.033423, 3.021743, 
    3.030881, 3.014246, 3.02355, 3.02891, 3.049653, 3.054221, 3.058465, 
    3.066857, 3.077653, 3.096659, 3.113264, 3.128478, 3.127361, 3.127754, 
    3.13116, 3.122729, 3.132546, 3.134197, 3.129883, 3.154745, 3.147787, 
    3.154907, 3.15038, 3.034518, 3.040194, 3.037126, 3.042897, 3.038831, 
    3.056941, 3.062386, 3.087956, 3.077441, 3.094186, 3.079138, 3.081801, 
    3.094737, 3.079949, 3.112349, 3.090359, 3.131293, 3.109241, 3.132679, 
    3.128412, 3.135478, 3.141817, 3.149747, 3.16405, 3.160733, 3.172721, 
    3.048667, 3.056055, 3.055403, 3.063146, 3.068882, 3.081339, 3.101398, 
    3.093844, 3.107721, 3.110513, 3.089433, 3.102365, 3.061006, 3.067662, 
    3.063696, 3.049251, 3.095586, 3.071744, 3.115873, 3.102878, 3.140913, 
    3.121958, 3.158909, 3.174446, 3.189113, 3.206328, 3.060091, 3.055065, 
    3.064067, 3.076557, 3.088174, 3.10367, 3.105258, 3.108169, 3.115716, 
    3.122073, 3.109092, 3.123668, 3.069211, 3.097661, 3.053168, 3.066519, 
    3.075819, 3.071735, 3.092981, 3.098004, 3.11848, 3.107882, 3.170608, 
    3.14316, 3.219476, 3.198056, 3.053311, 3.060073, 3.083695, 3.072439, 
    3.104706, 3.112687, 3.119184, 3.127507, 3.128405, 3.133344, 3.125253, 
    3.133024, 3.103703, 3.116781, 3.080986, 3.089672, 3.085674, 3.081293, 
    3.094827, 3.109296, 3.109603, 3.114254, 3.127391, 3.104837, 3.174149, 
    3.131546, 3.067459, 3.080542, 3.082411, 3.077336, 3.111886, 3.099335, 
    3.133224, 3.124038, 3.139098, 3.131608, 3.130507, 3.120908, 3.114944, 
    3.09991, 3.087717, 3.078071, 3.080312, 3.090914, 3.110182, 3.128488, 
    3.124471, 3.137952, 3.102358, 3.117249, 3.111488, 3.126524, 3.093644, 
    3.121636, 3.086519, 3.089586, 3.099087, 3.118263, 3.122512, 3.12706, 
    3.124253, 3.110672, 3.108449, 3.098855, 3.096211, 3.088918, 3.082891, 
    3.088398, 3.094189, 3.110676, 3.12559, 3.141908, 3.14591, 3.164531, 
    3.149426, 3.174385, 3.153162, 3.189964, 3.123259, 3.152534, 3.099518, 
    3.105214, 3.115537, 3.139303, 3.126453, 3.141483, 3.108362, 3.091282, 
    3.08687, 3.078658, 3.087058, 3.086374, 3.094427, 3.091838, 3.111225, 
    3.1008, 3.13048, 3.141364, 3.171464, 3.189891, 3.208727, 3.21707, 
    3.219613, 3.220676,
  2.987448, 3.004083, 3.000842, 3.014311, 3.006831, 3.015661, 2.990813, 
    3.004746, 2.995844, 2.988941, 3.040615, 3.014912, 3.067525, 3.050972, 
    3.092714, 3.064945, 3.098342, 3.091908, 3.111254, 3.105738, 3.130008, 
    3.113745, 3.142593, 3.126115, 3.128688, 3.11321, 3.020066, 3.037404, 
    3.019042, 3.021508, 3.020401, 3.006986, 3.000249, 2.986179, 2.988728, 
    2.999064, 3.022617, 3.014601, 3.034839, 3.03438, 3.057061, 3.046815, 
    3.085177, 3.074227, 3.10597, 3.097958, 3.105594, 3.103276, 3.105624, 
    3.093881, 3.098907, 3.088593, 3.048732, 3.060396, 3.025734, 3.005076, 
    2.991423, 2.981772, 2.983135, 2.985734, 2.999125, 3.011764, 3.021431, 
    3.027914, 3.034315, 3.053773, 3.064115, 3.087397, 3.083181, 3.090325, 
    3.097162, 3.108676, 3.106778, 3.111789, 3.090135, 3.104558, 3.080782, 
    3.087268, 3.036064, 3.016761, 3.008598, 3.001465, 2.984183, 2.996108, 
    2.991402, 3.002608, 3.00975, 3.006216, 3.028091, 3.019569, 3.064729, 
    3.045198, 3.096364, 3.084046, 3.099323, 3.091518, 3.104903, 3.092854, 
    3.113621, 3.118044, 3.115021, 3.126647, 3.092188, 3.105594, 3.006117, 
    3.006693, 3.009378, 2.997592, 2.996872, 2.986109, 2.995683, 2.99977, 
    3.010164, 3.01633, 3.022202, 3.03515, 3.049674, 3.070094, 3.084843, 
    3.094768, 3.088678, 3.094054, 3.088045, 3.085232, 3.116387, 3.098955, 
    3.124972, 3.123546, 3.111907, 3.123706, 3.007098, 3.003783, 2.992303, 
    3.001283, 2.98494, 2.994079, 2.999346, 3.019748, 3.024247, 3.028426, 
    3.036695, 3.047339, 3.066097, 3.082507, 3.09756, 3.096454, 3.096843, 
    3.100216, 3.09187, 3.101588, 3.103223, 3.098952, 3.123355, 3.116462, 
    3.123515, 3.119025, 3.00486, 3.010441, 3.007424, 3.0131, 3.009101, 
    3.026925, 3.032288, 3.057504, 3.047129, 3.063654, 3.048804, 3.05143, 
    3.064198, 3.049604, 3.081602, 3.059876, 3.100347, 3.078528, 3.101719, 
    3.097495, 3.104492, 3.110735, 3.118398, 3.132587, 3.129296, 3.141198, 
    3.018779, 3.026053, 3.02541, 3.033037, 3.03869, 3.050975, 3.070779, 
    3.063317, 3.077028, 3.079788, 3.058962, 3.071734, 3.030929, 3.037488, 
    3.03358, 3.019353, 3.065037, 3.041511, 3.085088, 3.072241, 3.109868, 
    3.091106, 3.127485, 3.142911, 3.157492, 3.174625, 3.030028, 3.025078, 
    3.033945, 3.046257, 3.057719, 3.073024, 3.074593, 3.07747, 3.084932, 
    3.091221, 3.078381, 3.092799, 3.039013, 3.067086, 3.02321, 3.03636, 
    3.045529, 3.041502, 3.062465, 3.067426, 3.087666, 3.077186, 3.139098, 
    3.112023, 3.187728, 3.166389, 3.02335, 3.03001, 3.053299, 3.042197, 
    3.074047, 3.081936, 3.088363, 3.096599, 3.097488, 3.102379, 3.094368, 
    3.102061, 3.073056, 3.085986, 3.050627, 3.059198, 3.055252, 3.05093, 
    3.064288, 3.078583, 3.078887, 3.083486, 3.096482, 3.074177, 3.142614, 
    3.100596, 3.037288, 3.050188, 3.052032, 3.047026, 3.081145, 3.068741, 
    3.102259, 3.093165, 3.108078, 3.100659, 3.099569, 3.090069, 3.084168, 
    3.069309, 3.057268, 3.047751, 3.049962, 3.060424, 3.079459, 3.097569, 
    3.093594, 3.106942, 3.071727, 3.086448, 3.080751, 3.095626, 3.063119, 
    3.090787, 3.056086, 3.059113, 3.068495, 3.087451, 3.091656, 3.096156, 
    3.093378, 3.079944, 3.077747, 3.068266, 3.065654, 3.058454, 3.052506, 
    3.05794, 3.063658, 3.079948, 3.094701, 3.110822, 3.114661, 3.133064, 
    3.118078, 3.142849, 3.121781, 3.158337, 3.092394, 3.121159, 3.068922, 
    3.074549, 3.084755, 3.10828, 3.095556, 3.110415, 3.077661, 3.060787, 
    3.056433, 3.04833, 3.056618, 3.055943, 3.063894, 3.061337, 3.080491, 
    3.070188, 3.099543, 3.1103, 3.139949, 3.158266, 3.177016, 3.185331, 
    3.187865, 3.188926,
  2.97751, 2.995923, 2.992336, 3.007253, 2.998966, 3.00875, 2.981246, 
    2.996657, 2.986807, 2.979177, 3.036467, 3.00792, 3.066467, 3.048, 
    3.094654, 3.063586, 3.100966, 3.09375, 3.115527, 3.109269, 3.137339, 
    3.118421, 3.152014, 3.132807, 3.135803, 3.1178, 3.013636, 3.032895, 
    3.012501, 3.015236, 3.014008, 2.999138, 2.991679, 2.976062, 2.978943, 
    2.990368, 3.016467, 3.007575, 3.030044, 3.029534, 3.054789, 3.04337, 
    3.08621, 3.073957, 3.109529, 3.100535, 3.109107, 3.106504, 3.109141, 
    3.095963, 3.1016, 3.090035, 3.045505, 3.058509, 3.019928, 2.997021, 
    2.98192, 2.971034, 2.972588, 2.975554, 2.990435, 3.004431, 3.015151, 
    3.022348, 3.029461, 3.051121, 3.062659, 3.088696, 3.083975, 3.091976, 
    3.099642, 3.112569, 3.110436, 3.116149, 3.091763, 3.107944, 3.08129, 
    3.088552, 3.031405, 3.009971, 3.000922, 2.993025, 2.973784, 2.987099, 
    2.981896, 2.99429, 3.002199, 2.998284, 3.022546, 3.013085, 3.063345, 
    3.041569, 3.098747, 3.084943, 3.102067, 3.093314, 3.108331, 3.094811, 
    3.118278, 3.123418, 3.119904, 3.133427, 3.094064, 3.109107, 2.998175, 
    2.998813, 3.001787, 2.98874, 2.987944, 2.975982, 2.986629, 2.991149, 
    3.002658, 3.009492, 3.016006, 3.030389, 3.046555, 3.069337, 3.085835, 
    3.096957, 3.090131, 3.096156, 3.089422, 3.086271, 3.121491, 3.101653, 
    3.131477, 3.129817, 3.116285, 3.130004, 2.999261, 2.99559, 2.982892, 
    2.992824, 2.974647, 2.984855, 2.99068, 3.013284, 3.018276, 3.022917, 
    3.032107, 3.043953, 3.064873, 3.08322, 3.100089, 3.098849, 3.099285, 
    3.103069, 3.093708, 3.104609, 3.106444, 3.10165, 3.129595, 3.121579, 
    3.129782, 3.124559, 2.996783, 3.002964, 2.999622, 3.005911, 3.00148, 
    3.021249, 3.027208, 3.055282, 3.04372, 3.062145, 3.045585, 3.048511, 
    3.062752, 3.046476, 3.082207, 3.057929, 3.103216, 3.078767, 3.104756, 
    3.100015, 3.107869, 3.114925, 3.123829, 3.140346, 3.136511, 3.150386, 
    3.012208, 3.020281, 3.019568, 3.028041, 3.034327, 3.048004, 3.070103, 
    3.061769, 3.077089, 3.080177, 3.056909, 3.07117, 3.025697, 3.032989, 
    3.028644, 3.012845, 3.063689, 3.037465, 3.086109, 3.071738, 3.113918, 
    3.092852, 3.134403, 3.152385, 3.169423, 3.188978, 3.024696, 3.019199, 
    3.02905, 3.042748, 3.055523, 3.072612, 3.074366, 3.077584, 3.085936, 
    3.092981, 3.078603, 3.09475, 3.034685, 3.065978, 3.017125, 3.031735, 
    3.041938, 3.037456, 3.060818, 3.066357, 3.088997, 3.077267, 3.147936, 
    3.11642, 3.203873, 3.179632, 3.017281, 3.024677, 3.050594, 3.038228, 
    3.073756, 3.082582, 3.089778, 3.09901, 3.100008, 3.105496, 3.096509, 
    3.10514, 3.072649, 3.087115, 3.047616, 3.057173, 3.052771, 3.047953, 
    3.062853, 3.078829, 3.07917, 3.084316, 3.098879, 3.073901, 3.152037, 
    3.103494, 3.032767, 3.047126, 3.049182, 3.043605, 3.081695, 3.067826, 
    3.105362, 3.09516, 3.111897, 3.103566, 3.102343, 3.091689, 3.08508, 
    3.06846, 3.05502, 3.044413, 3.046875, 3.058541, 3.079809, 3.100099, 
    3.095641, 3.110621, 3.071163, 3.087633, 3.081255, 3.097919, 3.061548, 
    3.092493, 3.053702, 3.057078, 3.067551, 3.088755, 3.093468, 3.098514, 
    3.095399, 3.080351, 3.077894, 3.067296, 3.064378, 3.056342, 3.04971, 
    3.05577, 3.06215, 3.080357, 3.096882, 3.115026, 3.119486, 3.1409, 
    3.123457, 3.152311, 3.127763, 3.17041, 3.094295, 3.12704, 3.068028, 
    3.074317, 3.085737, 3.112124, 3.097841, 3.114552, 3.077798, 3.058945, 
    3.054088, 3.045057, 3.054295, 3.053542, 3.062413, 3.059559, 3.080964, 
    3.069443, 3.102313, 3.114419, 3.148929, 3.170327, 3.191694, 3.201145, 
    3.204029, 3.205236,
  3.255258, 3.278734, 3.274146, 3.293253, 3.282629, 3.295176, 3.259992, 
    3.279673, 3.267085, 3.257358, 3.330445, 3.29411, 3.368219, 3.344929, 
    3.404013, 3.364576, 3.41207, 3.402861, 3.430716, 3.422692, 3.458801, 
    3.434431, 3.477803, 3.45295, 3.456816, 3.433633, 3.301454, 3.32597, 
    3.299994, 3.303512, 3.301932, 3.282849, 3.273307, 3.253474, 3.257059, 
    3.271632, 3.305096, 3.293667, 3.322401, 3.321763, 3.353476, 3.339108, 
    3.393258, 3.377701, 3.423026, 3.41152, 3.422484, 3.419152, 3.422528, 
    3.405683, 3.412881, 3.398128, 3.341791, 3.358167, 3.309551, 3.280139, 
    3.260852, 3.247287, 3.249199, 3.252849, 3.271718, 3.289632, 3.303402, 
    3.312671, 3.321671, 3.348856, 3.363406, 3.396422, 3.390417, 3.4006, 
    3.410379, 3.426921, 3.424188, 3.431513, 3.400329, 3.420995, 3.387005, 
    3.396239, 3.324104, 3.296743, 3.285135, 3.275027, 3.25067, 3.267457, 
    3.260822, 3.276645, 3.286771, 3.281756, 3.312925, 3.300745, 3.364272, 
    3.336847, 3.409236, 3.391647, 3.413477, 3.402304, 3.421491, 3.404214, 
    3.434247, 3.440854, 3.436336, 3.453749, 3.403261, 3.422485, 3.281616, 
    3.282433, 3.286243, 3.269552, 3.268536, 3.253376, 3.266858, 3.27263, 
    3.287359, 3.296128, 3.304502, 3.322834, 3.34311, 3.37185, 3.392782, 
    3.406951, 3.398249, 3.40593, 3.397346, 3.393337, 3.438376, 3.412949, 
    3.451234, 3.449094, 3.431688, 3.449335, 3.283007, 3.278308, 3.262091, 
    3.27477, 3.251733, 3.264594, 3.27203, 3.301001, 3.307425, 3.313404, 
    3.324984, 3.339841, 3.366204, 3.389458, 3.410949, 3.409366, 3.409923, 
    3.414758, 3.402807, 3.416727, 3.419075, 3.412945, 3.448808, 3.438489, 
    3.449049, 3.442322, 3.279834, 3.287752, 3.283469, 3.291532, 3.285849, 
    3.311254, 3.318854, 3.354097, 3.339548, 3.362757, 3.341891, 3.345571, 
    3.363523, 3.343012, 3.38817, 3.357434, 3.414946, 3.383802, 3.416916, 
    3.410856, 3.420899, 3.429943, 3.441383, 3.462687, 3.457731, 3.475691, 
    3.299619, 3.310007, 3.309088, 3.319896, 3.327763, 3.344933, 3.372819, 
    3.362282, 3.381673, 3.385592, 3.356149, 3.374171, 3.316966, 3.326087, 
    3.32065, 3.300437, 3.364707, 3.331697, 3.393131, 3.374889, 3.428651, 
    3.401716, 3.455009, 3.478284, 3.500459, 3.526731, 3.315699, 3.308613, 
    3.321158, 3.338327, 3.354401, 3.375997, 3.37822, 3.3823, 3.39291, 
    3.40188, 3.383594, 3.404136, 3.328213, 3.3676, 3.305942, 3.324518, 
    3.33731, 3.331686, 3.361081, 3.36808, 3.396805, 3.381898, 3.472513, 
    3.431861, 3.546629, 3.514072, 3.306144, 3.315673, 3.348192, 3.332655, 
    3.377447, 3.388646, 3.3978, 3.409572, 3.410846, 3.417863, 3.40638, 
    3.417407, 3.376043, 3.39441, 3.344445, 3.356481, 3.350934, 3.34487, 
    3.363651, 3.383881, 3.384313, 3.39085, 3.409404, 3.37763, 3.477833, 
    3.415302, 3.32581, 3.343829, 3.346415, 3.339404, 3.38752, 3.369937, 
    3.417691, 3.404659, 3.42606, 3.415394, 3.41383, 3.400234, 3.391822, 
    3.37074, 3.353767, 3.340419, 3.343513, 3.358207, 3.385125, 3.410963, 
    3.405272, 3.424425, 3.374161, 3.395069, 3.38696, 3.40818, 3.362003, 
    3.401258, 3.352106, 3.356362, 3.36959, 3.396498, 3.402501, 3.408939, 
    3.404963, 3.385813, 3.382694, 3.369267, 3.365578, 3.355434, 3.34708, 
    3.354712, 3.362762, 3.38582, 3.406856, 3.430072, 3.435799, 3.463403, 
    3.440904, 3.478188, 3.446447, 3.501747, 3.403555, 3.445516, 3.370193, 
    3.378158, 3.392657, 3.426351, 3.408079, 3.429465, 3.382571, 3.358717, 
    3.352593, 3.341228, 3.352854, 3.351905, 3.363095, 3.359491, 3.38659, 
    3.371983, 3.413792, 3.429294, 3.473801, 3.501639, 3.530418, 3.543027, 
    3.546836, 3.548431,
  3.812406, 3.852937, 3.844965, 3.878337, 3.859726, 3.88172, 3.820528, 
    3.854572, 3.832743, 3.816005, 3.945441, 3.879844, 4.01692, 3.972602, 
    4.084903, 4.009935, 4.100404, 4.082694, 4.136674, 4.120997, 4.192388, 
    4.14397, 4.230848, 4.18067, 4.188406, 4.142401, 3.892799, 3.937109, 
    3.890218, 3.896441, 3.893644, 3.860109, 3.843509, 3.809353, 3.815492, 
    3.840606, 3.899248, 3.879065, 3.930483, 3.929301, 3.988774, 3.961651, 
    4.064368, 4.034976, 4.121648, 4.099343, 4.120593, 4.114115, 4.120677, 
    4.088106, 4.101969, 4.073643, 3.966693, 3.997694, 3.90716, 3.855384, 
    3.822005, 3.798792, 3.802051, 3.808284, 3.840755, 3.871978, 3.896246, 
    3.912715, 3.929131, 3.980019, 4.007696, 4.07039, 4.058971, 4.078366, 
    4.097143, 4.129248, 4.123912, 4.138238, 4.077848, 4.117695, 4.05251, 
    4.070041, 3.933642, 3.884481, 3.864103, 3.846494, 3.804561, 3.833386, 
    3.821953, 3.849304, 3.866965, 3.858202, 3.913168, 3.891545, 4.009353, 
    3.95741, 4.09494, 4.061307, 4.103121, 4.081628, 4.11866, 4.085288, 
    4.143606, 4.156633, 4.147718, 4.182268, 4.083461, 4.120595, 3.857958, 
    3.859383, 3.866041, 3.837007, 3.835249, 3.809186, 3.832352, 3.842335, 
    3.867995, 3.883397, 3.898195, 3.931285, 3.969176, 4.023901, 4.063463, 
    4.090544, 4.073875, 4.088581, 4.072153, 4.064517, 4.151739, 4.1021, 
    4.177247, 4.172982, 4.138582, 4.173461, 3.860385, 3.852197, 3.824137, 
    3.846049, 3.806376, 3.828447, 3.841297, 3.891997, 3.90338, 3.914023, 
    3.935276, 3.963027, 4.013053, 4.057154, 4.098242, 4.09519, 4.096264, 
    4.105598, 4.082592, 4.109411, 4.113965, 4.102093, 4.172411, 4.151962, 
    4.172891, 4.159538, 3.854853, 3.868683, 3.861193, 3.875312, 3.865352, 
    3.910191, 3.923916, 3.989954, 3.962476, 4.006454, 3.966881, 3.973815, 
    4.007919, 3.968991, 4.054713, 3.996299, 4.105962, 4.046459, 4.109776, 
    4.098062, 4.117509, 4.135159, 4.15768, 4.200201, 4.19024, 4.226542, 
    3.889555, 3.90797, 3.906336, 3.925843, 3.940444, 3.972611, 4.025769, 
    4.005546, 4.042445, 4.049838, 3.993853, 4.028357, 3.920427, 3.937326, 
    3.927238, 3.891, 4.010185, 3.947776, 4.064125, 4.029702, 4.13263, 
    4.080501, 4.184787, 4.231832, 4.277551, 4.33226, 3.918119, 3.905491, 
    3.92818, 3.960185, 3.99053, 4.031778, 4.03595, 4.043627, 4.063706, 
    4.080816, 4.046066, 4.085137, 3.941281, 4.015732, 3.900748, 3.93441, 
    3.958277, 3.947755, 4.003252, 4.016653, 4.07112, 4.042869, 4.220078, 
    4.138921, 4.374619, 4.306071, 3.901106, 3.918074, 3.978765, 3.949565, 
    4.034498, 4.055615, 4.073017, 4.095587, 4.098043, 4.111612, 4.089446, 
    4.110729, 4.031865, 4.066559, 3.971692, 3.994484, 3.983953, 3.972491, 
    4.008164, 4.046607, 4.047422, 4.059793, 4.095263, 4.034843, 4.23091, 
    4.10665, 3.936811, 3.97053, 3.975406, 3.962206, 4.053484, 4.020221, 
    4.111279, 4.086142, 4.127565, 4.106829, 4.103805, 4.077667, 4.061638, 
    4.021766, 3.989326, 3.964112, 3.969935, 3.99777, 4.048956, 4.098268, 
    4.087317, 4.124374, 4.028339, 4.067813, 4.052425, 4.092906, 4.005013, 
    4.079626, 3.986174, 3.994257, 4.019554, 4.070534, 4.082006, 4.094367, 
    4.086725, 4.050256, 4.044369, 4.018932, 4.011855, 3.992493, 3.976662, 
    3.991121, 4.006465, 4.050269, 4.09036, 4.135413, 4.146659, 4.201644, 
    4.156732, 4.231634, 4.167717, 4.280235, 4.084025, 4.165868, 4.020714, 
    4.035834, 4.063224, 4.128133, 4.092713, 4.134223, 4.044138, 3.998743, 
    3.987098, 3.965633, 3.987593, 3.985794, 4.007101, 4.000218, 4.051726, 
    4.024158, 4.10373, 4.133889, 4.222696, 4.280009, 4.33991, 4.366787, 
    4.37507, 4.378548,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24858.28, 24879.12, 24875.04, 24892.09, 24882.59, 24893.81, 24862.47, 
    24879.96, 24868.76, 24860.13, 24925.93, 24892.85, 24961.35, 24939.45, 
    24994.93, 24957.91, 25002.54, 24993.84, 25020.24, 25012.61, 25047.14, 
    25023.78, 25065.53, 25041.51, 25045.23, 25023.02, 24899.44, 24921.77, 
    24898.13, 24901.28, 24899.87, 24882.79, 24874.29, 24856.69, 24859.87, 
    24872.8, 24902.71, 24892.46, 24918.45, 24917.86, 24947.46, 24934, 
    24984.81, 24970.26, 25012.92, 25002.02, 25012.41, 25009.24, 25012.45, 
    24996.5, 25003.3, 24989.39, 24936.51, 24951.87, 24906.71, 24880.37, 
    24863.23, 24851.21, 24852.9, 24856.14, 24872.88, 24888.85, 24901.19, 
    24909.52, 24917.77, 24943.12, 24956.8, 24987.78, 24982.15, 24991.71, 
    25000.94, 25016.63, 25014.03, 25021, 24991.46, 25010.99, 24978.95, 
    24987.61, 24920.03, 24895.21, 24884.83, 24875.82, 24854.21, 24869.09, 
    24863.2, 24877.26, 24886.29, 24881.81, 24909.75, 24898.8, 24957.62, 
    24931.89, 24999.86, 24983.3, 25003.87, 24993.32, 25011.46, 24995.12, 
    25023.61, 25029.91, 25025.6, 25042.28, 24994.22, 25012.41, 24881.69, 
    24882.42, 24885.82, 24870.95, 24870.05, 24856.61, 24868.56, 24873.69, 
    24886.82, 24894.66, 24902.17, 24918.85, 24937.74, 24964.78, 24984.37, 
    24997.7, 24989.5, 24996.73, 24988.65, 24984.89, 25027.55, 25003.37, 
    25039.86, 25037.8, 25021.17, 25038.04, 24882.93, 24878.74, 24864.33, 
    24875.59, 24855.15, 24866.55, 24873.15, 24899.03, 24904.8, 24910.18, 
    24920.85, 24934.69, 24959.44, 24981.25, 25001.47, 24999.98, 25000.51, 
    25005.08, 24993.79, 25006.95, 25009.17, 25003.36, 25037.53, 25027.65, 
    25037.76, 25031.32, 24880.1, 24887.17, 24883.35, 24890.55, 24885.47, 
    24908.25, 24915.16, 24948.04, 24934.41, 24956.19, 24936.6, 24940.05, 
    24956.91, 24937.65, 24980.04, 24951.18, 25005.26, 24975.96, 25007.12, 
    25001.39, 25010.9, 25019.5, 25030.42, 25050.88, 25046.11, 25063.48, 
    24897.79, 24907.12, 24906.3, 24916.13, 24923.43, 24939.45, 24965.7, 
    24955.74, 24973.97, 24977.63, 24949.97, 24966.97, 24913.41, 24921.88, 
    24916.83, 24898.52, 24958.03, 24927.09, 24984.69, 24967.64, 25018.28, 
    24992.76, 25043.49, 25066, 25087.68, 25113.45, 24912.25, 24905.87, 
    24917.3, 24933.28, 24948.33, 24968.67, 24970.74, 24974.55, 24984.48, 
    24992.92, 24975.76, 24995.04, 24923.85, 24960.76, 24903.47, 24920.42, 
    24932.32, 24927.08, 24954.61, 24961.21, 24988.14, 24974.18, 25060.39, 
    25021.33, 25133.29, 25101.09, 24903.65, 24912.23, 24942.5, 24927.98, 
    24970.02, 24980.49, 24989.08, 25000.17, 25001.38, 25008.02, 24997.16, 
    25007.59, 24968.71, 24985.89, 24938.99, 24950.28, 24945.07, 24939.39, 
    24957.04, 24976.03, 24976.43, 24982.55, 25000.02, 24970.19, 25065.56, 
    25005.59, 24921.62, 24938.42, 24940.84, 24934.28, 24979.43, 24962.97, 
    25007.86, 24995.54, 25015.81, 25005.68, 25004.2, 24991.37, 24983.46, 
    24963.73, 24947.73, 24935.23, 24938.12, 24951.91, 24977.19, 25001.49, 
    24996.11, 25014.25, 24966.96, 24986.51, 24978.91, 24998.86, 24955.48, 
    24992.33, 24946.17, 24950.17, 24962.64, 24987.85, 24993.5, 24999.58, 
    24995.82, 24977.84, 24974.92, 24962.34, 24958.85, 24949.3, 24941.46, 
    24948.62, 24956.2, 24977.84, 24997.61, 25019.63, 25025.09, 25051.58, 
    25029.96, 25065.9, 25035.27, 25088.95, 24994.5, 25034.38, 24963.21, 
    24970.69, 24984.25, 25016.09, 24998.76, 25019.05, 24974.8, 24952.39, 
    24946.63, 24935.98, 24946.88, 24945.98, 24956.51, 24953.12, 24978.56, 
    24964.9, 25004.16, 25018.89, 25061.64, 25088.84, 25117.06, 25129.64, 
    25133.49, 25135.11 ;

 HCSOI =
  24858.28, 24879.12, 24875.04, 24892.09, 24882.59, 24893.81, 24862.47, 
    24879.96, 24868.76, 24860.13, 24925.93, 24892.85, 24961.35, 24939.45, 
    24994.93, 24957.91, 25002.54, 24993.84, 25020.24, 25012.61, 25047.14, 
    25023.78, 25065.53, 25041.51, 25045.23, 25023.02, 24899.44, 24921.77, 
    24898.13, 24901.28, 24899.87, 24882.79, 24874.29, 24856.69, 24859.87, 
    24872.8, 24902.71, 24892.46, 24918.45, 24917.86, 24947.46, 24934, 
    24984.81, 24970.26, 25012.92, 25002.02, 25012.41, 25009.24, 25012.45, 
    24996.5, 25003.3, 24989.39, 24936.51, 24951.87, 24906.71, 24880.37, 
    24863.23, 24851.21, 24852.9, 24856.14, 24872.88, 24888.85, 24901.19, 
    24909.52, 24917.77, 24943.12, 24956.8, 24987.78, 24982.15, 24991.71, 
    25000.94, 25016.63, 25014.03, 25021, 24991.46, 25010.99, 24978.95, 
    24987.61, 24920.03, 24895.21, 24884.83, 24875.82, 24854.21, 24869.09, 
    24863.2, 24877.26, 24886.29, 24881.81, 24909.75, 24898.8, 24957.62, 
    24931.89, 24999.86, 24983.3, 25003.87, 24993.32, 25011.46, 24995.12, 
    25023.61, 25029.91, 25025.6, 25042.28, 24994.22, 25012.41, 24881.69, 
    24882.42, 24885.82, 24870.95, 24870.05, 24856.61, 24868.56, 24873.69, 
    24886.82, 24894.66, 24902.17, 24918.85, 24937.74, 24964.78, 24984.37, 
    24997.7, 24989.5, 24996.73, 24988.65, 24984.89, 25027.55, 25003.37, 
    25039.86, 25037.8, 25021.17, 25038.04, 24882.93, 24878.74, 24864.33, 
    24875.59, 24855.15, 24866.55, 24873.15, 24899.03, 24904.8, 24910.18, 
    24920.85, 24934.69, 24959.44, 24981.25, 25001.47, 24999.98, 25000.51, 
    25005.08, 24993.79, 25006.95, 25009.17, 25003.36, 25037.53, 25027.65, 
    25037.76, 25031.32, 24880.1, 24887.17, 24883.35, 24890.55, 24885.47, 
    24908.25, 24915.16, 24948.04, 24934.41, 24956.19, 24936.6, 24940.05, 
    24956.91, 24937.65, 24980.04, 24951.18, 25005.26, 24975.96, 25007.12, 
    25001.39, 25010.9, 25019.5, 25030.42, 25050.88, 25046.11, 25063.48, 
    24897.79, 24907.12, 24906.3, 24916.13, 24923.43, 24939.45, 24965.7, 
    24955.74, 24973.97, 24977.63, 24949.97, 24966.97, 24913.41, 24921.88, 
    24916.83, 24898.52, 24958.03, 24927.09, 24984.69, 24967.64, 25018.28, 
    24992.76, 25043.49, 25066, 25087.68, 25113.45, 24912.25, 24905.87, 
    24917.3, 24933.28, 24948.33, 24968.67, 24970.74, 24974.55, 24984.48, 
    24992.92, 24975.76, 24995.04, 24923.85, 24960.76, 24903.47, 24920.42, 
    24932.32, 24927.08, 24954.61, 24961.21, 24988.14, 24974.18, 25060.39, 
    25021.33, 25133.29, 25101.09, 24903.65, 24912.23, 24942.5, 24927.98, 
    24970.02, 24980.49, 24989.08, 25000.17, 25001.38, 25008.02, 24997.16, 
    25007.59, 24968.71, 24985.89, 24938.99, 24950.28, 24945.07, 24939.39, 
    24957.04, 24976.03, 24976.43, 24982.55, 25000.02, 24970.19, 25065.56, 
    25005.59, 24921.62, 24938.42, 24940.84, 24934.28, 24979.43, 24962.97, 
    25007.86, 24995.54, 25015.81, 25005.68, 25004.2, 24991.37, 24983.46, 
    24963.73, 24947.73, 24935.23, 24938.12, 24951.91, 24977.19, 25001.49, 
    24996.11, 25014.25, 24966.96, 24986.51, 24978.91, 24998.86, 24955.48, 
    24992.33, 24946.17, 24950.17, 24962.64, 24987.85, 24993.5, 24999.58, 
    24995.82, 24977.84, 24974.92, 24962.34, 24958.85, 24949.3, 24941.46, 
    24948.62, 24956.2, 24977.84, 24997.61, 25019.63, 25025.09, 25051.58, 
    25029.96, 25065.9, 25035.27, 25088.95, 24994.5, 25034.38, 24963.21, 
    24970.69, 24984.25, 25016.09, 24998.76, 25019.05, 24974.8, 24952.39, 
    24946.63, 24935.98, 24946.88, 24945.98, 24956.51, 24953.12, 24978.56, 
    24964.9, 25004.16, 25018.89, 25061.64, 25088.84, 25117.06, 25129.64, 
    25133.49, 25135.11 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 HR_vr =
  2.694543e-07, 2.70184e-07, 2.700423e-07, 2.706303e-07, 2.703043e-07, 
    2.706891e-07, 2.696024e-07, 2.702129e-07, 2.698233e-07, 2.695202e-07, 
    2.717696e-07, 2.706565e-07, 2.729249e-07, 2.722163e-07, 2.739952e-07, 
    2.728145e-07, 2.74233e-07, 2.739614e-07, 2.747792e-07, 2.74545e-07, 
    2.755894e-07, 2.748872e-07, 2.761305e-07, 2.754219e-07, 2.755327e-07, 
    2.74864e-07, 2.708809e-07, 2.716311e-07, 2.708364e-07, 2.709434e-07, 
    2.708954e-07, 2.703109e-07, 2.70016e-07, 2.693987e-07, 2.695108e-07, 
    2.699643e-07, 2.709916e-07, 2.706432e-07, 2.715213e-07, 2.715015e-07, 
    2.724776e-07, 2.720377e-07, 2.736763e-07, 2.73211e-07, 2.745548e-07, 
    2.742171e-07, 2.745389e-07, 2.744414e-07, 2.745402e-07, 2.740448e-07, 
    2.742571e-07, 2.738211e-07, 2.7212e-07, 2.726204e-07, 2.711269e-07, 
    2.70227e-07, 2.696292e-07, 2.692045e-07, 2.692645e-07, 2.693789e-07, 
    2.69967e-07, 2.705196e-07, 2.709403e-07, 2.712216e-07, 2.714986e-07, 
    2.723359e-07, 2.727792e-07, 2.737702e-07, 2.735917e-07, 2.738943e-07, 
    2.741835e-07, 2.746685e-07, 2.745887e-07, 2.748023e-07, 2.738865e-07, 
    2.744952e-07, 2.734899e-07, 2.73765e-07, 2.715731e-07, 2.707372e-07, 
    2.703809e-07, 2.700695e-07, 2.693107e-07, 2.698348e-07, 2.696282e-07, 
    2.701197e-07, 2.704317e-07, 2.702774e-07, 2.712293e-07, 2.708593e-07, 
    2.728055e-07, 2.719679e-07, 2.741498e-07, 2.736284e-07, 2.742747e-07, 
    2.73945e-07, 2.745098e-07, 2.740015e-07, 2.748818e-07, 2.750732e-07, 
    2.749424e-07, 2.754451e-07, 2.739733e-07, 2.745388e-07, 2.702731e-07, 
    2.702982e-07, 2.704155e-07, 2.698998e-07, 2.698683e-07, 2.693956e-07, 
    2.698163e-07, 2.699953e-07, 2.704498e-07, 2.707184e-07, 2.709737e-07, 
    2.715346e-07, 2.721604e-07, 2.730347e-07, 2.736622e-07, 2.740824e-07, 
    2.738248e-07, 2.740522e-07, 2.73798e-07, 2.736788e-07, 2.750014e-07, 
    2.74259e-07, 2.753728e-07, 2.753112e-07, 2.748073e-07, 2.753182e-07, 
    2.703159e-07, 2.701711e-07, 2.696679e-07, 2.700617e-07, 2.693441e-07, 
    2.697458e-07, 2.699766e-07, 2.708669e-07, 2.710626e-07, 2.712437e-07, 
    2.716014e-07, 2.720602e-07, 2.728641e-07, 2.73563e-07, 2.742004e-07, 
    2.741537e-07, 2.741701e-07, 2.743124e-07, 2.739599e-07, 2.743702e-07, 
    2.74439e-07, 2.74259e-07, 2.75303e-07, 2.750049e-07, 2.753099e-07, 
    2.751159e-07, 2.702182e-07, 2.704619e-07, 2.703302e-07, 2.705777e-07, 
    2.704033e-07, 2.711784e-07, 2.714106e-07, 2.724963e-07, 2.720511e-07, 
    2.727597e-07, 2.721232e-07, 2.72236e-07, 2.727824e-07, 2.721576e-07, 
    2.735243e-07, 2.725978e-07, 2.743179e-07, 2.733935e-07, 2.743757e-07, 
    2.741976e-07, 2.744926e-07, 2.747566e-07, 2.750887e-07, 2.757008e-07, 
    2.755591e-07, 2.760708e-07, 2.70825e-07, 2.711407e-07, 2.71113e-07, 
    2.714434e-07, 2.716875e-07, 2.722165e-07, 2.73064e-07, 2.727455e-07, 
    2.733303e-07, 2.734476e-07, 2.725592e-07, 2.731046e-07, 2.71352e-07, 
    2.716353e-07, 2.714667e-07, 2.708498e-07, 2.728187e-07, 2.718089e-07, 
    2.736725e-07, 2.731264e-07, 2.747189e-07, 2.739273e-07, 2.754811e-07, 
    2.761438e-07, 2.767675e-07, 2.774948e-07, 2.713131e-07, 2.710986e-07, 
    2.714827e-07, 2.720134e-07, 2.725058e-07, 2.731597e-07, 2.732266e-07, 
    2.73349e-07, 2.736661e-07, 2.739324e-07, 2.733876e-07, 2.739992e-07, 
    2.717007e-07, 2.729064e-07, 2.710174e-07, 2.715866e-07, 2.719821e-07, 
    2.718088e-07, 2.727091e-07, 2.729211e-07, 2.737817e-07, 2.73337e-07, 
    2.759802e-07, 2.748121e-07, 2.780485e-07, 2.771457e-07, 2.710237e-07, 
    2.713124e-07, 2.723161e-07, 2.718388e-07, 2.732034e-07, 2.735388e-07, 
    2.738115e-07, 2.741596e-07, 2.741973e-07, 2.744035e-07, 2.740655e-07, 
    2.743902e-07, 2.731611e-07, 2.737107e-07, 2.722016e-07, 2.725692e-07, 
    2.724002e-07, 2.722146e-07, 2.72787e-07, 2.733961e-07, 2.734093e-07, 
    2.736045e-07, 2.741536e-07, 2.732089e-07, 2.761303e-07, 2.743273e-07, 
    2.716271e-07, 2.721823e-07, 2.722619e-07, 2.720468e-07, 2.735052e-07, 
    2.729771e-07, 2.743985e-07, 2.740147e-07, 2.746435e-07, 2.743311e-07, 
    2.742851e-07, 2.738837e-07, 2.736336e-07, 2.730013e-07, 2.724865e-07, 
    2.72078e-07, 2.721731e-07, 2.726216e-07, 2.734334e-07, 2.742006e-07, 
    2.740326e-07, 2.745957e-07, 2.731045e-07, 2.737301e-07, 2.734883e-07, 
    2.741186e-07, 2.72737e-07, 2.73913e-07, 2.72436e-07, 2.725656e-07, 
    2.729666e-07, 2.737723e-07, 2.739508e-07, 2.741409e-07, 2.740237e-07, 
    2.73454e-07, 2.733608e-07, 2.72957e-07, 2.728453e-07, 2.725374e-07, 
    2.722823e-07, 2.725154e-07, 2.727599e-07, 2.734544e-07, 2.740794e-07, 
    2.747603e-07, 2.749269e-07, 2.757207e-07, 2.750743e-07, 2.761403e-07, 
    2.752336e-07, 2.768026e-07, 2.739814e-07, 2.752074e-07, 2.729849e-07, 
    2.732248e-07, 2.736581e-07, 2.746515e-07, 2.741157e-07, 2.747424e-07, 
    2.733571e-07, 2.72637e-07, 2.724508e-07, 2.721029e-07, 2.724587e-07, 
    2.724298e-07, 2.727702e-07, 2.726609e-07, 2.734774e-07, 2.730389e-07, 
    2.742839e-07, 2.747375e-07, 2.760171e-07, 2.768001e-07, 2.775965e-07, 
    2.779476e-07, 2.780545e-07, 2.780991e-07,
  2.336853e-07, 2.345734e-07, 2.344009e-07, 2.351167e-07, 2.347197e-07, 
    2.351883e-07, 2.338655e-07, 2.346086e-07, 2.341343e-07, 2.337654e-07, 
    2.365042e-07, 2.351486e-07, 2.37911e-07, 2.370478e-07, 2.392149e-07, 
    2.377766e-07, 2.395046e-07, 2.391736e-07, 2.401701e-07, 2.398847e-07, 
    2.411577e-07, 2.403017e-07, 2.418172e-07, 2.409535e-07, 2.410886e-07, 
    2.402735e-07, 2.354218e-07, 2.363355e-07, 2.353676e-07, 2.354979e-07, 
    2.354395e-07, 2.347279e-07, 2.34369e-07, 2.336175e-07, 2.33754e-07, 
    2.34306e-07, 2.355565e-07, 2.351323e-07, 2.362014e-07, 2.361773e-07, 
    2.373661e-07, 2.368302e-07, 2.388263e-07, 2.382594e-07, 2.398966e-07, 
    2.394851e-07, 2.398773e-07, 2.397584e-07, 2.398788e-07, 2.392753e-07, 
    2.395339e-07, 2.390027e-07, 2.369306e-07, 2.3754e-07, 2.357213e-07, 
    2.346259e-07, 2.338981e-07, 2.333811e-07, 2.334542e-07, 2.335935e-07, 
    2.343092e-07, 2.349818e-07, 2.35494e-07, 2.358365e-07, 2.361738e-07, 
    2.371937e-07, 2.377335e-07, 2.389407e-07, 2.387231e-07, 2.390919e-07, 
    2.394442e-07, 2.400352e-07, 2.39938e-07, 2.401983e-07, 2.390823e-07, 
    2.39824e-07, 2.385991e-07, 2.389343e-07, 2.362649e-07, 2.352468e-07, 
    2.348132e-07, 2.34434e-07, 2.335104e-07, 2.341483e-07, 2.338969e-07, 
    2.344951e-07, 2.348749e-07, 2.346871e-07, 2.358458e-07, 2.353955e-07, 
    2.377655e-07, 2.367454e-07, 2.394031e-07, 2.387678e-07, 2.395553e-07, 
    2.391536e-07, 2.398418e-07, 2.392225e-07, 2.402952e-07, 2.405285e-07, 
    2.40369e-07, 2.409816e-07, 2.391881e-07, 2.398772e-07, 2.346818e-07, 
    2.347124e-07, 2.348552e-07, 2.342275e-07, 2.341891e-07, 2.336137e-07, 
    2.341258e-07, 2.343437e-07, 2.348969e-07, 2.352239e-07, 2.355347e-07, 
    2.362177e-07, 2.369798e-07, 2.380446e-07, 2.38809e-07, 2.39321e-07, 
    2.390071e-07, 2.392842e-07, 2.389745e-07, 2.388292e-07, 2.40441e-07, 
    2.395363e-07, 2.408935e-07, 2.408185e-07, 2.402044e-07, 2.40827e-07, 
    2.347339e-07, 2.345576e-07, 2.339451e-07, 2.344245e-07, 2.33551e-07, 
    2.3404e-07, 2.34321e-07, 2.354048e-07, 2.356429e-07, 2.358634e-07, 
    2.36299e-07, 2.368577e-07, 2.378369e-07, 2.386882e-07, 2.394647e-07, 
    2.394079e-07, 2.394279e-07, 2.396012e-07, 2.391717e-07, 2.396717e-07, 
    2.397555e-07, 2.395362e-07, 2.408085e-07, 2.404452e-07, 2.408169e-07, 
    2.405804e-07, 2.34615e-07, 2.349116e-07, 2.347513e-07, 2.350527e-07, 
    2.348403e-07, 2.35784e-07, 2.360667e-07, 2.373889e-07, 2.368466e-07, 
    2.377097e-07, 2.369344e-07, 2.370718e-07, 2.377376e-07, 2.369763e-07, 
    2.386411e-07, 2.375126e-07, 2.396079e-07, 2.384818e-07, 2.396784e-07, 
    2.394613e-07, 2.398208e-07, 2.401426e-07, 2.405473e-07, 2.412934e-07, 
    2.411207e-07, 2.417445e-07, 2.353537e-07, 2.357381e-07, 2.357043e-07, 
    2.361065e-07, 2.364038e-07, 2.370481e-07, 2.380803e-07, 2.376923e-07, 
    2.384047e-07, 2.385476e-07, 2.374654e-07, 2.381299e-07, 2.359953e-07, 
    2.363404e-07, 2.36135e-07, 2.353839e-07, 2.377816e-07, 2.365518e-07, 
    2.388216e-07, 2.381563e-07, 2.400967e-07, 2.391321e-07, 2.410256e-07, 
    2.418336e-07, 2.425939e-07, 2.43481e-07, 2.359479e-07, 2.356868e-07, 
    2.361544e-07, 2.368007e-07, 2.374004e-07, 2.381969e-07, 2.382784e-07, 
    2.384275e-07, 2.388137e-07, 2.391383e-07, 2.384745e-07, 2.392196e-07, 
    2.364202e-07, 2.378883e-07, 2.355879e-07, 2.362811e-07, 2.367627e-07, 
    2.365516e-07, 2.37648e-07, 2.379062e-07, 2.389547e-07, 2.384129e-07, 
    2.416342e-07, 2.402103e-07, 2.441562e-07, 2.430552e-07, 2.355955e-07, 
    2.359471e-07, 2.371694e-07, 2.36588e-07, 2.382501e-07, 2.386587e-07, 
    2.389909e-07, 2.394151e-07, 2.39461e-07, 2.397123e-07, 2.393004e-07, 
    2.39696e-07, 2.381986e-07, 2.388681e-07, 2.370299e-07, 2.374776e-07, 
    2.372717e-07, 2.370458e-07, 2.377429e-07, 2.384849e-07, 2.38501e-07, 
    2.387387e-07, 2.394081e-07, 2.382568e-07, 2.418174e-07, 2.396198e-07, 
    2.363303e-07, 2.370065e-07, 2.371033e-07, 2.368414e-07, 2.386178e-07, 
    2.379745e-07, 2.397061e-07, 2.392385e-07, 2.400047e-07, 2.39624e-07, 
    2.39568e-07, 2.390788e-07, 2.387742e-07, 2.380039e-07, 2.373769e-07, 
    2.368794e-07, 2.369951e-07, 2.375415e-07, 2.385304e-07, 2.39465e-07, 
    2.392604e-07, 2.399465e-07, 2.381297e-07, 2.388918e-07, 2.385973e-07, 
    2.393652e-07, 2.37682e-07, 2.391149e-07, 2.373153e-07, 2.374733e-07, 
    2.379617e-07, 2.389434e-07, 2.391607e-07, 2.393923e-07, 2.392494e-07, 
    2.385555e-07, 2.384418e-07, 2.379499e-07, 2.378139e-07, 2.374389e-07, 
    2.371282e-07, 2.37412e-07, 2.3771e-07, 2.385559e-07, 2.393174e-07, 
    2.401471e-07, 2.403501e-07, 2.413179e-07, 2.405299e-07, 2.418296e-07, 
    2.407244e-07, 2.426369e-07, 2.391982e-07, 2.406922e-07, 2.37984e-07, 
    2.382762e-07, 2.388042e-07, 2.400146e-07, 2.393616e-07, 2.401254e-07, 
    2.384374e-07, 2.375602e-07, 2.373334e-07, 2.369096e-07, 2.373431e-07, 
    2.373078e-07, 2.377224e-07, 2.375892e-07, 2.385839e-07, 2.380498e-07, 
    2.395665e-07, 2.401194e-07, 2.416791e-07, 2.426337e-07, 2.436048e-07, 
    2.440331e-07, 2.441634e-07, 2.442178e-07,
  2.190408e-07, 2.200111e-07, 2.198226e-07, 2.206048e-07, 2.20171e-07, 
    2.206831e-07, 2.192376e-07, 2.200496e-07, 2.195313e-07, 2.191283e-07, 
    2.221216e-07, 2.206397e-07, 2.236599e-07, 2.227158e-07, 2.250865e-07, 
    2.23513e-07, 2.254036e-07, 2.250412e-07, 2.261318e-07, 2.258195e-07, 
    2.272133e-07, 2.26276e-07, 2.279356e-07, 2.269896e-07, 2.271376e-07, 
    2.26245e-07, 2.209381e-07, 2.219371e-07, 2.208789e-07, 2.210214e-07, 
    2.209575e-07, 2.201799e-07, 2.197878e-07, 2.189667e-07, 2.191158e-07, 
    2.197189e-07, 2.210855e-07, 2.206218e-07, 2.217903e-07, 2.21764e-07, 
    2.230639e-07, 2.224779e-07, 2.246612e-07, 2.24041e-07, 2.258325e-07, 
    2.253822e-07, 2.258114e-07, 2.256812e-07, 2.258131e-07, 2.251525e-07, 
    2.254355e-07, 2.248542e-07, 2.225876e-07, 2.23254e-07, 2.212656e-07, 
    2.200685e-07, 2.192732e-07, 2.187086e-07, 2.187884e-07, 2.189406e-07, 
    2.197225e-07, 2.204573e-07, 2.210171e-07, 2.213914e-07, 2.217602e-07, 
    2.228755e-07, 2.234658e-07, 2.247865e-07, 2.245483e-07, 2.249518e-07, 
    2.253373e-07, 2.259843e-07, 2.258778e-07, 2.261627e-07, 2.249413e-07, 
    2.257531e-07, 2.244126e-07, 2.247794e-07, 2.2186e-07, 2.207469e-07, 
    2.202733e-07, 2.198588e-07, 2.188498e-07, 2.195466e-07, 2.19272e-07, 
    2.199254e-07, 2.203405e-07, 2.201352e-07, 2.214017e-07, 2.209094e-07, 
    2.235008e-07, 2.223851e-07, 2.252924e-07, 2.245972e-07, 2.25459e-07, 
    2.250193e-07, 2.257725e-07, 2.250947e-07, 2.262688e-07, 2.265243e-07, 
    2.263497e-07, 2.270204e-07, 2.250571e-07, 2.258113e-07, 2.201295e-07, 
    2.201629e-07, 2.203189e-07, 2.196332e-07, 2.195912e-07, 2.189626e-07, 
    2.19522e-07, 2.197601e-07, 2.203646e-07, 2.207219e-07, 2.210616e-07, 
    2.218082e-07, 2.226415e-07, 2.238061e-07, 2.246423e-07, 2.252025e-07, 
    2.248591e-07, 2.251623e-07, 2.248233e-07, 2.246644e-07, 2.264285e-07, 
    2.254382e-07, 2.269239e-07, 2.268418e-07, 2.261695e-07, 2.26851e-07, 
    2.201865e-07, 2.199938e-07, 2.193247e-07, 2.198484e-07, 2.188942e-07, 
    2.194283e-07, 2.197353e-07, 2.209196e-07, 2.211798e-07, 2.214209e-07, 
    2.218971e-07, 2.225079e-07, 2.235788e-07, 2.245101e-07, 2.253598e-07, 
    2.252976e-07, 2.253195e-07, 2.255092e-07, 2.250391e-07, 2.255863e-07, 
    2.256781e-07, 2.254381e-07, 2.268308e-07, 2.26433e-07, 2.2684e-07, 
    2.265811e-07, 2.200564e-07, 2.203806e-07, 2.202054e-07, 2.205348e-07, 
    2.203027e-07, 2.213341e-07, 2.216432e-07, 2.230889e-07, 2.224958e-07, 
    2.234397e-07, 2.225918e-07, 2.22742e-07, 2.234703e-07, 2.226376e-07, 
    2.244587e-07, 2.232242e-07, 2.255165e-07, 2.242844e-07, 2.255937e-07, 
    2.253561e-07, 2.257495e-07, 2.261017e-07, 2.265448e-07, 2.273619e-07, 
    2.271727e-07, 2.278558e-07, 2.208637e-07, 2.212839e-07, 2.21247e-07, 
    2.216866e-07, 2.220117e-07, 2.227161e-07, 2.238451e-07, 2.234207e-07, 
    2.241999e-07, 2.243562e-07, 2.231724e-07, 2.238993e-07, 2.215651e-07, 
    2.219424e-07, 2.217178e-07, 2.208968e-07, 2.235184e-07, 2.221735e-07, 
    2.246561e-07, 2.239282e-07, 2.260515e-07, 2.249959e-07, 2.270686e-07, 
    2.279536e-07, 2.287863e-07, 2.297585e-07, 2.215132e-07, 2.212278e-07, 
    2.217389e-07, 2.224457e-07, 2.231014e-07, 2.239726e-07, 2.240618e-07, 
    2.242249e-07, 2.246474e-07, 2.250026e-07, 2.242764e-07, 2.250916e-07, 
    2.220297e-07, 2.236351e-07, 2.211198e-07, 2.218775e-07, 2.224041e-07, 
    2.221732e-07, 2.233722e-07, 2.236546e-07, 2.248017e-07, 2.242089e-07, 
    2.277351e-07, 2.26176e-07, 2.304985e-07, 2.292918e-07, 2.21128e-07, 
    2.215123e-07, 2.228488e-07, 2.222131e-07, 2.240308e-07, 2.244778e-07, 
    2.248413e-07, 2.253055e-07, 2.253557e-07, 2.256307e-07, 2.2518e-07, 
    2.25613e-07, 2.239745e-07, 2.247069e-07, 2.226962e-07, 2.231858e-07, 
    2.229606e-07, 2.227135e-07, 2.23476e-07, 2.242878e-07, 2.243053e-07, 
    2.245654e-07, 2.252982e-07, 2.240381e-07, 2.27936e-07, 2.255298e-07, 
    2.219312e-07, 2.226707e-07, 2.227765e-07, 2.2249e-07, 2.24433e-07, 
    2.237293e-07, 2.25624e-07, 2.251122e-07, 2.259508e-07, 2.255341e-07, 
    2.254728e-07, 2.249375e-07, 2.246041e-07, 2.237615e-07, 2.230756e-07, 
    2.225316e-07, 2.226581e-07, 2.232557e-07, 2.243375e-07, 2.253602e-07, 
    2.251362e-07, 2.258871e-07, 2.238991e-07, 2.247329e-07, 2.244107e-07, 
    2.252508e-07, 2.234094e-07, 2.249773e-07, 2.230083e-07, 2.23181e-07, 
    2.237153e-07, 2.247894e-07, 2.250271e-07, 2.252806e-07, 2.251242e-07, 
    2.243649e-07, 2.242406e-07, 2.237024e-07, 2.235537e-07, 2.231434e-07, 
    2.228037e-07, 2.231141e-07, 2.2344e-07, 2.243653e-07, 2.251987e-07, 
    2.261067e-07, 2.263289e-07, 2.273888e-07, 2.265259e-07, 2.279494e-07, 
    2.26739e-07, 2.288337e-07, 2.250683e-07, 2.267036e-07, 2.237397e-07, 
    2.240593e-07, 2.246371e-07, 2.259618e-07, 2.252469e-07, 2.26083e-07, 
    2.242357e-07, 2.232763e-07, 2.230281e-07, 2.225647e-07, 2.230387e-07, 
    2.230001e-07, 2.234536e-07, 2.233079e-07, 2.24396e-07, 2.238116e-07, 
    2.254713e-07, 2.260764e-07, 2.277842e-07, 2.2883e-07, 2.298941e-07, 
    2.303635e-07, 2.305064e-07, 2.305661e-07,
  2.100066e-07, 2.11004e-07, 2.108101e-07, 2.116145e-07, 2.111684e-07, 
    2.11695e-07, 2.102088e-07, 2.110436e-07, 2.105107e-07, 2.100964e-07, 
    2.131753e-07, 2.116504e-07, 2.147591e-07, 2.137868e-07, 2.162291e-07, 
    2.146078e-07, 2.16556e-07, 2.161824e-07, 2.173068e-07, 2.169847e-07, 
    2.184227e-07, 2.174555e-07, 2.191681e-07, 2.181918e-07, 2.183445e-07, 
    2.174236e-07, 2.119574e-07, 2.129855e-07, 2.118964e-07, 2.120431e-07, 
    2.119773e-07, 2.111776e-07, 2.107745e-07, 2.099304e-07, 2.100836e-07, 
    2.107036e-07, 2.12109e-07, 2.11632e-07, 2.128342e-07, 2.12807e-07, 
    2.141452e-07, 2.135419e-07, 2.157906e-07, 2.151516e-07, 2.169982e-07, 
    2.165338e-07, 2.169764e-07, 2.168422e-07, 2.169781e-07, 2.162971e-07, 
    2.165889e-07, 2.159896e-07, 2.136548e-07, 2.143411e-07, 2.122942e-07, 
    2.110632e-07, 2.102454e-07, 2.096651e-07, 2.097472e-07, 2.099036e-07, 
    2.107072e-07, 2.114628e-07, 2.120386e-07, 2.124237e-07, 2.128031e-07, 
    2.139514e-07, 2.145592e-07, 2.159198e-07, 2.156744e-07, 2.160903e-07, 
    2.164876e-07, 2.171546e-07, 2.170449e-07, 2.173387e-07, 2.160793e-07, 
    2.169163e-07, 2.155345e-07, 2.159125e-07, 2.129061e-07, 2.117607e-07, 
    2.112736e-07, 2.108474e-07, 2.098102e-07, 2.105265e-07, 2.102441e-07, 
    2.109159e-07, 2.113427e-07, 2.111316e-07, 2.124342e-07, 2.119278e-07, 
    2.145952e-07, 2.134464e-07, 2.164413e-07, 2.157248e-07, 2.16613e-07, 
    2.161598e-07, 2.169363e-07, 2.162375e-07, 2.174481e-07, 2.177117e-07, 
    2.175316e-07, 2.182235e-07, 2.161987e-07, 2.169763e-07, 2.111257e-07, 
    2.111601e-07, 2.113205e-07, 2.106154e-07, 2.105723e-07, 2.099262e-07, 
    2.105011e-07, 2.107459e-07, 2.113674e-07, 2.11735e-07, 2.120844e-07, 
    2.128525e-07, 2.137103e-07, 2.149096e-07, 2.157712e-07, 2.163486e-07, 
    2.159946e-07, 2.163072e-07, 2.159577e-07, 2.157939e-07, 2.176129e-07, 
    2.165916e-07, 2.18124e-07, 2.180392e-07, 2.173457e-07, 2.180487e-07, 
    2.111843e-07, 2.109862e-07, 2.102983e-07, 2.108366e-07, 2.098558e-07, 
    2.104048e-07, 2.107205e-07, 2.119384e-07, 2.12206e-07, 2.12454e-07, 
    2.12944e-07, 2.135727e-07, 2.146756e-07, 2.15635e-07, 2.165107e-07, 
    2.164466e-07, 2.164692e-07, 2.166648e-07, 2.161802e-07, 2.167443e-07, 
    2.16839e-07, 2.165915e-07, 2.180278e-07, 2.176175e-07, 2.180374e-07, 
    2.177702e-07, 2.110506e-07, 2.113839e-07, 2.112038e-07, 2.115425e-07, 
    2.113039e-07, 2.123648e-07, 2.126829e-07, 2.14171e-07, 2.135604e-07, 
    2.145323e-07, 2.136591e-07, 2.138138e-07, 2.145639e-07, 2.137063e-07, 
    2.155821e-07, 2.143104e-07, 2.166724e-07, 2.154026e-07, 2.167519e-07, 
    2.16507e-07, 2.169126e-07, 2.172758e-07, 2.177328e-07, 2.185759e-07, 
    2.183807e-07, 2.190857e-07, 2.118808e-07, 2.123131e-07, 2.122751e-07, 
    2.127274e-07, 2.13062e-07, 2.137871e-07, 2.149498e-07, 2.145126e-07, 
    2.153153e-07, 2.154764e-07, 2.14257e-07, 2.150057e-07, 2.126024e-07, 
    2.129907e-07, 2.127595e-07, 2.119149e-07, 2.146133e-07, 2.132286e-07, 
    2.157854e-07, 2.150354e-07, 2.17224e-07, 2.161357e-07, 2.182732e-07, 
    2.191867e-07, 2.200465e-07, 2.210509e-07, 2.12549e-07, 2.122553e-07, 
    2.127813e-07, 2.135088e-07, 2.141839e-07, 2.150812e-07, 2.15173e-07, 
    2.153411e-07, 2.157765e-07, 2.161425e-07, 2.153942e-07, 2.162343e-07, 
    2.130807e-07, 2.147335e-07, 2.121443e-07, 2.12924e-07, 2.134659e-07, 
    2.132282e-07, 2.144626e-07, 2.147536e-07, 2.159355e-07, 2.153246e-07, 
    2.189613e-07, 2.173525e-07, 2.218157e-07, 2.205688e-07, 2.121527e-07, 
    2.12548e-07, 2.139238e-07, 2.132693e-07, 2.151411e-07, 2.156017e-07, 
    2.159762e-07, 2.164549e-07, 2.165065e-07, 2.167901e-07, 2.163254e-07, 
    2.167718e-07, 2.150831e-07, 2.158378e-07, 2.137666e-07, 2.142708e-07, 
    2.140388e-07, 2.137844e-07, 2.145696e-07, 2.15406e-07, 2.154239e-07, 
    2.15692e-07, 2.164475e-07, 2.151487e-07, 2.191688e-07, 2.166863e-07, 
    2.129791e-07, 2.137405e-07, 2.138493e-07, 2.135544e-07, 2.155556e-07, 
    2.148305e-07, 2.167832e-07, 2.162555e-07, 2.171201e-07, 2.166905e-07, 
    2.166273e-07, 2.160755e-07, 2.157319e-07, 2.148638e-07, 2.141573e-07, 
    2.135971e-07, 2.137274e-07, 2.143428e-07, 2.154571e-07, 2.165112e-07, 
    2.162803e-07, 2.170544e-07, 2.150054e-07, 2.158646e-07, 2.155325e-07, 
    2.163985e-07, 2.14501e-07, 2.161167e-07, 2.140879e-07, 2.142658e-07, 
    2.148161e-07, 2.159229e-07, 2.161678e-07, 2.164292e-07, 2.162679e-07, 
    2.154854e-07, 2.153572e-07, 2.148028e-07, 2.146496e-07, 2.142271e-07, 
    2.138773e-07, 2.141969e-07, 2.145325e-07, 2.154858e-07, 2.163447e-07, 
    2.17281e-07, 2.175101e-07, 2.186038e-07, 2.177135e-07, 2.191826e-07, 
    2.179335e-07, 2.200957e-07, 2.162104e-07, 2.178968e-07, 2.148412e-07, 
    2.151704e-07, 2.157659e-07, 2.171316e-07, 2.163944e-07, 2.172565e-07, 
    2.153522e-07, 2.14364e-07, 2.141083e-07, 2.136312e-07, 2.141192e-07, 
    2.140795e-07, 2.145465e-07, 2.143964e-07, 2.155174e-07, 2.149153e-07, 
    2.166257e-07, 2.172497e-07, 2.190118e-07, 2.200918e-07, 2.211909e-07, 
    2.216761e-07, 2.218238e-07, 2.218855e-07,
  2.030027e-07, 2.039495e-07, 2.037654e-07, 2.045295e-07, 2.041056e-07, 
    2.04606e-07, 2.031946e-07, 2.039871e-07, 2.034812e-07, 2.030879e-07, 
    2.060135e-07, 2.045636e-07, 2.075213e-07, 2.065953e-07, 2.089227e-07, 
    2.073772e-07, 2.092346e-07, 2.088781e-07, 2.099513e-07, 2.096438e-07, 
    2.110176e-07, 2.100933e-07, 2.117303e-07, 2.107968e-07, 2.109428e-07, 
    2.100628e-07, 2.048552e-07, 2.058329e-07, 2.047973e-07, 2.049367e-07, 
    2.048741e-07, 2.041143e-07, 2.037316e-07, 2.029304e-07, 2.030758e-07, 
    2.036643e-07, 2.049994e-07, 2.04546e-07, 2.056888e-07, 2.05663e-07, 
    2.069365e-07, 2.063622e-07, 2.085045e-07, 2.078952e-07, 2.096566e-07, 
    2.092134e-07, 2.096358e-07, 2.095077e-07, 2.096375e-07, 2.089875e-07, 
    2.092659e-07, 2.086942e-07, 2.064697e-07, 2.071231e-07, 2.051754e-07, 
    2.040058e-07, 2.032294e-07, 2.026787e-07, 2.027566e-07, 2.02905e-07, 
    2.036677e-07, 2.043853e-07, 2.049324e-07, 2.052985e-07, 2.056593e-07, 
    2.067521e-07, 2.073309e-07, 2.086277e-07, 2.083936e-07, 2.087903e-07, 
    2.091693e-07, 2.09806e-07, 2.097012e-07, 2.099818e-07, 2.087798e-07, 
    2.095785e-07, 2.082602e-07, 2.086206e-07, 2.057575e-07, 2.046683e-07, 
    2.042057e-07, 2.038008e-07, 2.028164e-07, 2.034961e-07, 2.032281e-07, 
    2.038658e-07, 2.042711e-07, 2.040706e-07, 2.053085e-07, 2.048271e-07, 
    2.073652e-07, 2.062714e-07, 2.091251e-07, 2.084416e-07, 2.09289e-07, 
    2.088565e-07, 2.095976e-07, 2.089306e-07, 2.100862e-07, 2.10338e-07, 
    2.10166e-07, 2.10827e-07, 2.088937e-07, 2.096358e-07, 2.04065e-07, 
    2.040977e-07, 2.042501e-07, 2.035806e-07, 2.035396e-07, 2.029264e-07, 
    2.03472e-07, 2.037044e-07, 2.042946e-07, 2.046439e-07, 2.049759e-07, 
    2.057063e-07, 2.065225e-07, 2.076647e-07, 2.084859e-07, 2.090367e-07, 
    2.086989e-07, 2.089971e-07, 2.086638e-07, 2.085076e-07, 2.102437e-07, 
    2.092685e-07, 2.107319e-07, 2.106509e-07, 2.099885e-07, 2.1066e-07, 
    2.041207e-07, 2.039325e-07, 2.032795e-07, 2.037905e-07, 2.028596e-07, 
    2.033806e-07, 2.036803e-07, 2.048372e-07, 2.050915e-07, 2.053274e-07, 
    2.057933e-07, 2.063915e-07, 2.074417e-07, 2.083561e-07, 2.091914e-07, 
    2.091301e-07, 2.091517e-07, 2.093384e-07, 2.08876e-07, 2.094143e-07, 
    2.095047e-07, 2.092684e-07, 2.106401e-07, 2.10248e-07, 2.106492e-07, 
    2.103939e-07, 2.039937e-07, 2.043103e-07, 2.041392e-07, 2.04461e-07, 
    2.042343e-07, 2.052426e-07, 2.05545e-07, 2.069612e-07, 2.063798e-07, 
    2.073052e-07, 2.064737e-07, 2.06621e-07, 2.073354e-07, 2.065186e-07, 
    2.083057e-07, 2.070939e-07, 2.093456e-07, 2.081346e-07, 2.094216e-07, 
    2.091878e-07, 2.095749e-07, 2.099217e-07, 2.103582e-07, 2.11164e-07, 
    2.109773e-07, 2.116515e-07, 2.047824e-07, 2.051934e-07, 2.051572e-07, 
    2.055873e-07, 2.059056e-07, 2.065955e-07, 2.07703e-07, 2.072864e-07, 
    2.080512e-07, 2.082049e-07, 2.070429e-07, 2.077562e-07, 2.054685e-07, 
    2.058378e-07, 2.056179e-07, 2.048149e-07, 2.073824e-07, 2.060641e-07, 
    2.084995e-07, 2.077845e-07, 2.098723e-07, 2.088336e-07, 2.108746e-07, 
    2.117482e-07, 2.125709e-07, 2.135331e-07, 2.054177e-07, 2.051384e-07, 
    2.056385e-07, 2.063308e-07, 2.069733e-07, 2.078281e-07, 2.079156e-07, 
    2.080758e-07, 2.084909e-07, 2.0884e-07, 2.081265e-07, 2.089276e-07, 
    2.059235e-07, 2.074969e-07, 2.050328e-07, 2.057744e-07, 2.062899e-07, 
    2.060637e-07, 2.072388e-07, 2.075159e-07, 2.086427e-07, 2.080601e-07, 
    2.115325e-07, 2.09995e-07, 2.142662e-07, 2.130711e-07, 2.050408e-07, 
    2.054167e-07, 2.067258e-07, 2.061028e-07, 2.078852e-07, 2.083244e-07, 
    2.086814e-07, 2.091381e-07, 2.091874e-07, 2.09458e-07, 2.090146e-07, 
    2.094405e-07, 2.0783e-07, 2.085494e-07, 2.06576e-07, 2.070561e-07, 
    2.068352e-07, 2.06593e-07, 2.073407e-07, 2.081378e-07, 2.081548e-07, 
    2.084105e-07, 2.091313e-07, 2.078925e-07, 2.117312e-07, 2.093591e-07, 
    2.058267e-07, 2.065513e-07, 2.066548e-07, 2.06374e-07, 2.082803e-07, 
    2.075893e-07, 2.094514e-07, 2.089479e-07, 2.09773e-07, 2.093629e-07, 
    2.093026e-07, 2.087761e-07, 2.084484e-07, 2.07621e-07, 2.069481e-07, 
    2.064147e-07, 2.065387e-07, 2.071247e-07, 2.081865e-07, 2.091919e-07, 
    2.089716e-07, 2.097103e-07, 2.077559e-07, 2.085751e-07, 2.082584e-07, 
    2.090842e-07, 2.072754e-07, 2.088156e-07, 2.068819e-07, 2.070514e-07, 
    2.075756e-07, 2.086307e-07, 2.088642e-07, 2.091136e-07, 2.089597e-07, 
    2.082135e-07, 2.080913e-07, 2.075628e-07, 2.07417e-07, 2.070145e-07, 
    2.066814e-07, 2.069857e-07, 2.073054e-07, 2.082138e-07, 2.09033e-07, 
    2.099267e-07, 2.101455e-07, 2.111908e-07, 2.103398e-07, 2.117444e-07, 
    2.105502e-07, 2.126181e-07, 2.089049e-07, 2.10515e-07, 2.075994e-07, 
    2.079132e-07, 2.08481e-07, 2.097841e-07, 2.090804e-07, 2.099034e-07, 
    2.080865e-07, 2.071449e-07, 2.069014e-07, 2.064472e-07, 2.069117e-07, 
    2.068739e-07, 2.073186e-07, 2.071757e-07, 2.08244e-07, 2.0767e-07, 
    2.093011e-07, 2.098969e-07, 2.115808e-07, 2.126143e-07, 2.136671e-07, 
    2.141323e-07, 2.142739e-07, 2.143331e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  9.652399e-13, 9.678468e-13, 9.673404e-13, 9.69441e-13, 9.682762e-13, 
    9.696512e-13, 9.65769e-13, 9.679499e-13, 9.665581e-13, 9.654752e-13, 
    9.735113e-13, 9.695348e-13, 9.776379e-13, 9.751066e-13, 9.814612e-13, 
    9.772438e-13, 9.823108e-13, 9.813404e-13, 9.842616e-13, 9.834251e-13, 
    9.871558e-13, 9.846476e-13, 9.890884e-13, 9.865574e-13, 9.869532e-13, 
    9.845646e-13, 9.703362e-13, 9.730164e-13, 9.701772e-13, 9.705597e-13, 
    9.703883e-13, 9.683001e-13, 9.672466e-13, 9.650411e-13, 9.654418e-13, 
    9.670618e-13, 9.707316e-13, 9.69487e-13, 9.726239e-13, 9.725531e-13, 
    9.760401e-13, 9.744686e-13, 9.803222e-13, 9.786601e-13, 9.834602e-13, 
    9.822538e-13, 9.834034e-13, 9.830549e-13, 9.834079e-13, 9.816385e-13, 
    9.823967e-13, 9.808393e-13, 9.747628e-13, 9.765501e-13, 9.712151e-13, 
    9.680003e-13, 9.658645e-13, 9.643473e-13, 9.645619e-13, 9.649706e-13, 
    9.670714e-13, 9.690454e-13, 9.705484e-13, 9.715532e-13, 9.725429e-13, 
    9.755342e-13, 9.771176e-13, 9.806576e-13, 9.800199e-13, 9.811007e-13, 
    9.821338e-13, 9.838663e-13, 9.835813e-13, 9.843441e-13, 9.810728e-13, 
    9.832472e-13, 9.796564e-13, 9.80639e-13, 9.728094e-13, 9.69823e-13, 
    9.685502e-13, 9.674376e-13, 9.647268e-13, 9.66599e-13, 9.658611e-13, 
    9.676169e-13, 9.687315e-13, 9.681804e-13, 9.715807e-13, 9.702592e-13, 
    9.772114e-13, 9.742194e-13, 9.820133e-13, 9.801509e-13, 9.824597e-13, 
    9.812819e-13, 9.832993e-13, 9.814838e-13, 9.846282e-13, 9.85312e-13, 
    9.848446e-13, 9.866401e-13, 9.813831e-13, 9.83403e-13, 9.681649e-13, 
    9.682548e-13, 9.686737e-13, 9.668314e-13, 9.667188e-13, 9.650299e-13, 
    9.66533e-13, 9.671725e-13, 9.687963e-13, 9.697559e-13, 9.706678e-13, 
    9.726715e-13, 9.74907e-13, 9.7803e-13, 9.802715e-13, 9.817727e-13, 
    9.808526e-13, 9.816649e-13, 9.807566e-13, 9.803309e-13, 9.850556e-13, 
    9.824036e-13, 9.86382e-13, 9.861621e-13, 9.843621e-13, 9.861868e-13, 
    9.683179e-13, 9.678006e-13, 9.660028e-13, 9.674099e-13, 9.64846e-13, 
    9.662811e-13, 9.671057e-13, 9.702864e-13, 9.709851e-13, 9.716322e-13, 
    9.729102e-13, 9.74549e-13, 9.774209e-13, 9.799172e-13, 9.82194e-13, 
    9.820273e-13, 9.820859e-13, 9.82594e-13, 9.813349e-13, 9.828006e-13, 
    9.830463e-13, 9.824036e-13, 9.861326e-13, 9.850679e-13, 9.861574e-13, 
    9.854643e-13, 9.679688e-13, 9.688393e-13, 9.683689e-13, 9.692532e-13, 
    9.6863e-13, 9.71399e-13, 9.722285e-13, 9.761069e-13, 9.745166e-13, 
    9.770478e-13, 9.747741e-13, 9.75177e-13, 9.771292e-13, 9.748971e-13, 
    9.797791e-13, 9.764694e-13, 9.826137e-13, 9.793118e-13, 9.828205e-13, 
    9.821842e-13, 9.832379e-13, 9.841808e-13, 9.853672e-13, 9.875536e-13, 
    9.870476e-13, 9.888752e-13, 9.701366e-13, 9.712643e-13, 9.711655e-13, 
    9.723455e-13, 9.732176e-13, 9.751076e-13, 9.781349e-13, 9.769971e-13, 
    9.790861e-13, 9.79505e-13, 9.763315e-13, 9.782801e-13, 9.720191e-13, 
    9.730312e-13, 9.724291e-13, 9.702253e-13, 9.772586e-13, 9.736515e-13, 
    9.803085e-13, 9.783578e-13, 9.840464e-13, 9.812186e-13, 9.867688e-13, 
    9.891361e-13, 9.913638e-13, 9.939616e-13, 9.7188e-13, 9.71114e-13, 
    9.724859e-13, 9.743818e-13, 9.761409e-13, 9.784767e-13, 9.787158e-13, 
    9.79153e-13, 9.802855e-13, 9.81237e-13, 9.792907e-13, 9.814755e-13, 
    9.73265e-13, 9.775718e-13, 9.708239e-13, 9.728572e-13, 9.742703e-13, 
    9.73651e-13, 9.768671e-13, 9.776243e-13, 9.806985e-13, 9.791101e-13, 
    9.885516e-13, 9.843794e-13, 9.959391e-13, 9.927146e-13, 9.708461e-13, 
    9.718776e-13, 9.754633e-13, 9.73758e-13, 9.786328e-13, 9.798309e-13, 
    9.808048e-13, 9.820484e-13, 9.821831e-13, 9.829196e-13, 9.817124e-13, 
    9.828721e-13, 9.784816e-13, 9.804448e-13, 9.750543e-13, 9.763672e-13, 
    9.757635e-13, 9.751008e-13, 9.771456e-13, 9.793212e-13, 9.793685e-13, 
    9.800655e-13, 9.820272e-13, 9.786526e-13, 9.89088e-13, 9.826478e-13, 
    9.730018e-13, 9.749854e-13, 9.752695e-13, 9.745013e-13, 9.797108e-13, 
    9.778245e-13, 9.829017e-13, 9.815308e-13, 9.837768e-13, 9.826609e-13, 
    9.824966e-13, 9.810628e-13, 9.801694e-13, 9.779108e-13, 9.760718e-13, 
    9.746128e-13, 9.749522e-13, 9.765546e-13, 9.794544e-13, 9.821949e-13, 
    9.815947e-13, 9.836062e-13, 9.782796e-13, 9.805143e-13, 9.796506e-13, 
    9.819021e-13, 9.769667e-13, 9.811677e-13, 9.758914e-13, 9.763546e-13, 
    9.77787e-13, 9.806652e-13, 9.813027e-13, 9.819817e-13, 9.815629e-13, 
    9.795281e-13, 9.791949e-13, 9.777524e-13, 9.773535e-13, 9.762538e-13, 
    9.753425e-13, 9.76175e-13, 9.770486e-13, 9.795293e-13, 9.817621e-13, 
    9.841942e-13, 9.847893e-13, 9.876248e-13, 9.853158e-13, 9.891237e-13, 
    9.85885e-13, 9.914891e-13, 9.814121e-13, 9.857913e-13, 9.778525e-13, 
    9.787092e-13, 9.802573e-13, 9.838056e-13, 9.818915e-13, 9.841302e-13, 
    9.791819e-13, 9.766094e-13, 9.759444e-13, 9.747013e-13, 9.759728e-13, 
    9.758695e-13, 9.770854e-13, 9.766947e-13, 9.796117e-13, 9.780453e-13, 
    9.824923e-13, 9.841127e-13, 9.886835e-13, 9.914802e-13, 9.943246e-13, 
    9.955787e-13, 9.959604e-13, 9.961199e-13 ;

 LITR1C =
  3.066846e-05, 3.066834e-05, 3.066836e-05, 3.066827e-05, 3.066832e-05, 
    3.066826e-05, 3.066843e-05, 3.066833e-05, 3.06684e-05, 3.066845e-05, 
    3.066808e-05, 3.066826e-05, 3.06679e-05, 3.066801e-05, 3.066772e-05, 
    3.066791e-05, 3.066768e-05, 3.066773e-05, 3.066759e-05, 3.066763e-05, 
    3.066746e-05, 3.066758e-05, 3.066738e-05, 3.066749e-05, 3.066747e-05, 
    3.066758e-05, 3.066823e-05, 3.06681e-05, 3.066823e-05, 3.066822e-05, 
    3.066822e-05, 3.066832e-05, 3.066837e-05, 3.066846e-05, 3.066845e-05, 
    3.066837e-05, 3.066821e-05, 3.066826e-05, 3.066812e-05, 3.066812e-05, 
    3.066797e-05, 3.066804e-05, 3.066777e-05, 3.066785e-05, 3.066763e-05, 
    3.066768e-05, 3.066763e-05, 3.066765e-05, 3.066763e-05, 3.066771e-05, 
    3.066768e-05, 3.066775e-05, 3.066802e-05, 3.066794e-05, 3.066819e-05, 
    3.066833e-05, 3.066843e-05, 3.06685e-05, 3.066849e-05, 3.066847e-05, 
    3.066837e-05, 3.066829e-05, 3.066822e-05, 3.066817e-05, 3.066812e-05, 
    3.066799e-05, 3.066792e-05, 3.066776e-05, 3.066779e-05, 3.066774e-05, 
    3.066769e-05, 3.066761e-05, 3.066763e-05, 3.066759e-05, 3.066774e-05, 
    3.066764e-05, 3.06678e-05, 3.066776e-05, 3.066811e-05, 3.066825e-05, 
    3.066831e-05, 3.066836e-05, 3.066848e-05, 3.066839e-05, 3.066843e-05, 
    3.066835e-05, 3.06683e-05, 3.066832e-05, 3.066817e-05, 3.066823e-05, 
    3.066791e-05, 3.066805e-05, 3.06677e-05, 3.066778e-05, 3.066768e-05, 
    3.066773e-05, 3.066764e-05, 3.066772e-05, 3.066758e-05, 3.066755e-05, 
    3.066757e-05, 3.066749e-05, 3.066772e-05, 3.066763e-05, 3.066833e-05, 
    3.066832e-05, 3.06683e-05, 3.066838e-05, 3.066839e-05, 3.066847e-05, 
    3.06684e-05, 3.066837e-05, 3.06683e-05, 3.066825e-05, 3.066821e-05, 
    3.066812e-05, 3.066802e-05, 3.066788e-05, 3.066778e-05, 3.066771e-05, 
    3.066775e-05, 3.066771e-05, 3.066775e-05, 3.066777e-05, 3.066756e-05, 
    3.066768e-05, 3.06675e-05, 3.066751e-05, 3.066759e-05, 3.066751e-05, 
    3.066832e-05, 3.066834e-05, 3.066842e-05, 3.066836e-05, 3.066847e-05, 
    3.066841e-05, 3.066837e-05, 3.066823e-05, 3.066819e-05, 3.066816e-05, 
    3.066811e-05, 3.066803e-05, 3.06679e-05, 3.066779e-05, 3.066769e-05, 
    3.06677e-05, 3.066769e-05, 3.066767e-05, 3.066773e-05, 3.066766e-05, 
    3.066765e-05, 3.066768e-05, 3.066751e-05, 3.066756e-05, 3.066751e-05, 
    3.066754e-05, 3.066833e-05, 3.066829e-05, 3.066831e-05, 3.066827e-05, 
    3.06683e-05, 3.066818e-05, 3.066814e-05, 3.066796e-05, 3.066804e-05, 
    3.066792e-05, 3.066802e-05, 3.0668e-05, 3.066792e-05, 3.066802e-05, 
    3.06678e-05, 3.066795e-05, 3.066767e-05, 3.066782e-05, 3.066766e-05, 
    3.066769e-05, 3.066764e-05, 3.06676e-05, 3.066755e-05, 3.066744e-05, 
    3.066747e-05, 3.066739e-05, 3.066823e-05, 3.066818e-05, 3.066819e-05, 
    3.066814e-05, 3.06681e-05, 3.066801e-05, 3.066787e-05, 3.066792e-05, 
    3.066783e-05, 3.066781e-05, 3.066795e-05, 3.066787e-05, 3.066815e-05, 
    3.06681e-05, 3.066813e-05, 3.066823e-05, 3.066791e-05, 3.066807e-05, 
    3.066777e-05, 3.066786e-05, 3.06676e-05, 3.066773e-05, 3.066748e-05, 
    3.066738e-05, 3.066727e-05, 3.066716e-05, 3.066815e-05, 3.066819e-05, 
    3.066813e-05, 3.066804e-05, 3.066796e-05, 3.066786e-05, 3.066784e-05, 
    3.066783e-05, 3.066778e-05, 3.066773e-05, 3.066782e-05, 3.066772e-05, 
    3.066809e-05, 3.06679e-05, 3.06682e-05, 3.066811e-05, 3.066805e-05, 
    3.066807e-05, 3.066793e-05, 3.06679e-05, 3.066776e-05, 3.066783e-05, 
    3.06674e-05, 3.066759e-05, 3.066707e-05, 3.066721e-05, 3.06682e-05, 
    3.066815e-05, 3.066799e-05, 3.066807e-05, 3.066785e-05, 3.066779e-05, 
    3.066775e-05, 3.06677e-05, 3.066769e-05, 3.066766e-05, 3.066771e-05, 
    3.066766e-05, 3.066786e-05, 3.066777e-05, 3.066801e-05, 3.066795e-05, 
    3.066798e-05, 3.066801e-05, 3.066792e-05, 3.066782e-05, 3.066782e-05, 
    3.066779e-05, 3.06677e-05, 3.066785e-05, 3.066738e-05, 3.066767e-05, 
    3.06681e-05, 3.066802e-05, 3.0668e-05, 3.066804e-05, 3.06678e-05, 
    3.066788e-05, 3.066766e-05, 3.066772e-05, 3.066762e-05, 3.066767e-05, 
    3.066767e-05, 3.066774e-05, 3.066778e-05, 3.066788e-05, 3.066796e-05, 
    3.066803e-05, 3.066802e-05, 3.066794e-05, 3.066781e-05, 3.066769e-05, 
    3.066771e-05, 3.066762e-05, 3.066787e-05, 3.066776e-05, 3.06678e-05, 
    3.06677e-05, 3.066792e-05, 3.066774e-05, 3.066797e-05, 3.066795e-05, 
    3.066789e-05, 3.066776e-05, 3.066773e-05, 3.06677e-05, 3.066772e-05, 
    3.066781e-05, 3.066782e-05, 3.066789e-05, 3.066791e-05, 3.066796e-05, 
    3.0668e-05, 3.066796e-05, 3.066792e-05, 3.066781e-05, 3.066771e-05, 
    3.06676e-05, 3.066757e-05, 3.066744e-05, 3.066755e-05, 3.066738e-05, 
    3.066752e-05, 3.066727e-05, 3.066772e-05, 3.066752e-05, 3.066788e-05, 
    3.066784e-05, 3.066778e-05, 3.066762e-05, 3.06677e-05, 3.06676e-05, 
    3.066783e-05, 3.066794e-05, 3.066797e-05, 3.066803e-05, 3.066797e-05, 
    3.066798e-05, 3.066792e-05, 3.066794e-05, 3.06678e-05, 3.066788e-05, 
    3.066767e-05, 3.06676e-05, 3.066739e-05, 3.066727e-05, 3.066714e-05, 
    3.066708e-05, 3.066707e-05, 3.066706e-05 ;

 LITR1C_TO_SOIL1C =
  6.428924e-13, 6.446283e-13, 6.442911e-13, 6.456899e-13, 6.449143e-13, 
    6.458299e-13, 6.432447e-13, 6.44697e-13, 6.437701e-13, 6.43049e-13, 
    6.484004e-13, 6.457524e-13, 6.511484e-13, 6.494627e-13, 6.536944e-13, 
    6.508859e-13, 6.542601e-13, 6.536139e-13, 6.555592e-13, 6.550022e-13, 
    6.574864e-13, 6.558162e-13, 6.587734e-13, 6.57088e-13, 6.573516e-13, 
    6.55761e-13, 6.462861e-13, 6.480708e-13, 6.461802e-13, 6.464348e-13, 
    6.463207e-13, 6.449302e-13, 6.442286e-13, 6.427599e-13, 6.430268e-13, 
    6.441056e-13, 6.465494e-13, 6.457206e-13, 6.478095e-13, 6.477623e-13, 
    6.500844e-13, 6.490378e-13, 6.529358e-13, 6.518291e-13, 6.550255e-13, 
    6.542222e-13, 6.549877e-13, 6.547557e-13, 6.549907e-13, 6.538124e-13, 
    6.543173e-13, 6.532803e-13, 6.492338e-13, 6.50424e-13, 6.468713e-13, 
    6.447306e-13, 6.433083e-13, 6.422979e-13, 6.424408e-13, 6.42713e-13, 
    6.441119e-13, 6.454265e-13, 6.464274e-13, 6.470965e-13, 6.477556e-13, 
    6.497475e-13, 6.508019e-13, 6.531593e-13, 6.527345e-13, 6.534543e-13, 
    6.541423e-13, 6.552959e-13, 6.551062e-13, 6.556141e-13, 6.534356e-13, 
    6.548837e-13, 6.524924e-13, 6.531468e-13, 6.47933e-13, 6.459443e-13, 
    6.450968e-13, 6.443559e-13, 6.425506e-13, 6.437974e-13, 6.43306e-13, 
    6.444752e-13, 6.452175e-13, 6.448505e-13, 6.471148e-13, 6.462348e-13, 
    6.508643e-13, 6.48872e-13, 6.54062e-13, 6.528218e-13, 6.543592e-13, 
    6.53575e-13, 6.549183e-13, 6.537094e-13, 6.558033e-13, 6.562586e-13, 
    6.559474e-13, 6.571431e-13, 6.536423e-13, 6.549875e-13, 6.448401e-13, 
    6.449e-13, 6.45179e-13, 6.439522e-13, 6.438771e-13, 6.427526e-13, 
    6.437534e-13, 6.441793e-13, 6.452606e-13, 6.458996e-13, 6.465068e-13, 
    6.478412e-13, 6.493298e-13, 6.514095e-13, 6.529022e-13, 6.539018e-13, 
    6.532891e-13, 6.538301e-13, 6.532252e-13, 6.529417e-13, 6.560879e-13, 
    6.543219e-13, 6.569712e-13, 6.568247e-13, 6.556262e-13, 6.568412e-13, 
    6.44942e-13, 6.445975e-13, 6.434004e-13, 6.443373e-13, 6.4263e-13, 
    6.435857e-13, 6.441348e-13, 6.462529e-13, 6.467182e-13, 6.471491e-13, 
    6.480001e-13, 6.490914e-13, 6.510039e-13, 6.526662e-13, 6.541823e-13, 
    6.540714e-13, 6.541104e-13, 6.544487e-13, 6.536103e-13, 6.545864e-13, 
    6.5475e-13, 6.543219e-13, 6.568051e-13, 6.560962e-13, 6.568216e-13, 
    6.563601e-13, 6.447095e-13, 6.452892e-13, 6.44976e-13, 6.455649e-13, 
    6.451499e-13, 6.469937e-13, 6.475461e-13, 6.501289e-13, 6.490698e-13, 
    6.507554e-13, 6.492413e-13, 6.495096e-13, 6.508096e-13, 6.493233e-13, 
    6.525742e-13, 6.503703e-13, 6.544619e-13, 6.52263e-13, 6.545995e-13, 
    6.541758e-13, 6.548775e-13, 6.555054e-13, 6.562954e-13, 6.577514e-13, 
    6.574144e-13, 6.586315e-13, 6.461531e-13, 6.469041e-13, 6.468383e-13, 
    6.47624e-13, 6.482049e-13, 6.494634e-13, 6.514794e-13, 6.507217e-13, 
    6.521127e-13, 6.523917e-13, 6.502784e-13, 6.51576e-13, 6.474067e-13, 
    6.480808e-13, 6.476797e-13, 6.462122e-13, 6.508958e-13, 6.484937e-13, 
    6.529268e-13, 6.516277e-13, 6.554159e-13, 6.535328e-13, 6.572288e-13, 
    6.588052e-13, 6.602886e-13, 6.620186e-13, 6.473141e-13, 6.46804e-13, 
    6.477176e-13, 6.489801e-13, 6.501515e-13, 6.517069e-13, 6.518662e-13, 
    6.521573e-13, 6.529114e-13, 6.53545e-13, 6.52249e-13, 6.537039e-13, 
    6.482364e-13, 6.511043e-13, 6.466108e-13, 6.479648e-13, 6.489058e-13, 
    6.484934e-13, 6.506351e-13, 6.511394e-13, 6.531865e-13, 6.521287e-13, 
    6.584159e-13, 6.556376e-13, 6.633354e-13, 6.611882e-13, 6.466257e-13, 
    6.473126e-13, 6.497003e-13, 6.485647e-13, 6.518109e-13, 6.526087e-13, 
    6.532573e-13, 6.540854e-13, 6.541751e-13, 6.546655e-13, 6.538617e-13, 
    6.546339e-13, 6.517102e-13, 6.530175e-13, 6.494279e-13, 6.503022e-13, 
    6.499002e-13, 6.494588e-13, 6.508205e-13, 6.522693e-13, 6.523008e-13, 
    6.52765e-13, 6.540713e-13, 6.51824e-13, 6.587732e-13, 6.544845e-13, 
    6.480611e-13, 6.49382e-13, 6.495712e-13, 6.490596e-13, 6.525288e-13, 
    6.512726e-13, 6.546536e-13, 6.537407e-13, 6.552363e-13, 6.544933e-13, 
    6.543839e-13, 6.53429e-13, 6.528341e-13, 6.513301e-13, 6.501055e-13, 
    6.491339e-13, 6.493599e-13, 6.50427e-13, 6.52358e-13, 6.541829e-13, 
    6.537833e-13, 6.551227e-13, 6.515757e-13, 6.530638e-13, 6.524886e-13, 
    6.539879e-13, 6.507014e-13, 6.53499e-13, 6.499853e-13, 6.502938e-13, 
    6.512477e-13, 6.531643e-13, 6.535888e-13, 6.54041e-13, 6.537621e-13, 
    6.524071e-13, 6.521852e-13, 6.512246e-13, 6.50959e-13, 6.502267e-13, 
    6.496199e-13, 6.501742e-13, 6.50756e-13, 6.524079e-13, 6.538947e-13, 
    6.555143e-13, 6.559105e-13, 6.577988e-13, 6.562612e-13, 6.587969e-13, 
    6.566403e-13, 6.603721e-13, 6.536617e-13, 6.565778e-13, 6.512912e-13, 
    6.518618e-13, 6.528927e-13, 6.552555e-13, 6.539809e-13, 6.554717e-13, 
    6.521766e-13, 6.504635e-13, 6.500206e-13, 6.491929e-13, 6.500395e-13, 
    6.499707e-13, 6.507804e-13, 6.505203e-13, 6.524627e-13, 6.514197e-13, 
    6.54381e-13, 6.554601e-13, 6.585038e-13, 6.603661e-13, 6.622603e-13, 
    6.630954e-13, 6.633495e-13, 6.634557e-13 ;

 LITR1C_vr =
  0.001751201, 0.001751194, 0.001751195, 0.00175119, 0.001751193, 
    0.001751189, 0.001751199, 0.001751194, 0.001751197, 0.0017512, 
    0.001751179, 0.001751189, 0.001751169, 0.001751175, 0.001751159, 
    0.001751169, 0.001751156, 0.001751159, 0.001751151, 0.001751153, 
    0.001751144, 0.00175115, 0.001751139, 0.001751145, 0.001751144, 
    0.001751151, 0.001751187, 0.00175118, 0.001751188, 0.001751187, 
    0.001751187, 0.001751193, 0.001751195, 0.001751201, 0.0017512, 
    0.001751196, 0.001751186, 0.00175119, 0.001751181, 0.001751182, 
    0.001751173, 0.001751177, 0.001751162, 0.001751166, 0.001751153, 
    0.001751157, 0.001751154, 0.001751154, 0.001751154, 0.001751158, 
    0.001751156, 0.00175116, 0.001751176, 0.001751171, 0.001751185, 
    0.001751193, 0.001751199, 0.001751203, 0.001751202, 0.001751201, 
    0.001751196, 0.001751191, 0.001751187, 0.001751184, 0.001751182, 
    0.001751174, 0.00175117, 0.001751161, 0.001751162, 0.00175116, 
    0.001751157, 0.001751152, 0.001751153, 0.001751151, 0.00175116, 
    0.001751154, 0.001751163, 0.001751161, 0.001751181, 0.001751189, 
    0.001751192, 0.001751195, 0.001751202, 0.001751197, 0.001751199, 
    0.001751194, 0.001751191, 0.001751193, 0.001751184, 0.001751188, 
    0.00175117, 0.001751177, 0.001751157, 0.001751162, 0.001751156, 
    0.001751159, 0.001751154, 0.001751159, 0.00175115, 0.001751149, 
    0.00175115, 0.001751145, 0.001751159, 0.001751154, 0.001751193, 
    0.001751193, 0.001751192, 0.001751196, 0.001751197, 0.001751201, 
    0.001751197, 0.001751196, 0.001751191, 0.001751189, 0.001751186, 
    0.001751181, 0.001751175, 0.001751167, 0.001751162, 0.001751158, 
    0.00175116, 0.001751158, 0.00175116, 0.001751162, 0.001751149, 
    0.001751156, 0.001751146, 0.001751146, 0.001751151, 0.001751146, 
    0.001751193, 0.001751194, 0.001751199, 0.001751195, 0.001751202, 
    0.001751198, 0.001751196, 0.001751187, 0.001751186, 0.001751184, 
    0.001751181, 0.001751176, 0.001751169, 0.001751163, 0.001751157, 
    0.001751157, 0.001751157, 0.001751156, 0.001751159, 0.001751155, 
    0.001751155, 0.001751156, 0.001751147, 0.001751149, 0.001751147, 
    0.001751148, 0.001751193, 0.001751191, 0.001751192, 0.00175119, 
    0.001751192, 0.001751185, 0.001751182, 0.001751172, 0.001751177, 
    0.00175117, 0.001751176, 0.001751175, 0.00175117, 0.001751176, 
    0.001751163, 0.001751172, 0.001751156, 0.001751164, 0.001751155, 
    0.001751157, 0.001751154, 0.001751152, 0.001751148, 0.001751143, 
    0.001751144, 0.001751139, 0.001751188, 0.001751185, 0.001751185, 
    0.001751182, 0.00175118, 0.001751175, 0.001751167, 0.00175117, 
    0.001751165, 0.001751164, 0.001751172, 0.001751167, 0.001751183, 
    0.00175118, 0.001751182, 0.001751188, 0.001751169, 0.001751179, 
    0.001751162, 0.001751167, 0.001751152, 0.001751159, 0.001751145, 
    0.001751139, 0.001751133, 0.001751126, 0.001751183, 0.001751185, 
    0.001751182, 0.001751177, 0.001751172, 0.001751166, 0.001751166, 
    0.001751165, 0.001751162, 0.001751159, 0.001751164, 0.001751159, 
    0.00175118, 0.001751169, 0.001751186, 0.001751181, 0.001751177, 
    0.001751179, 0.00175117, 0.001751169, 0.001751161, 0.001751165, 
    0.00175114, 0.001751151, 0.001751121, 0.00175113, 0.001751186, 
    0.001751183, 0.001751174, 0.001751179, 0.001751166, 0.001751163, 
    0.00175116, 0.001751157, 0.001751157, 0.001751155, 0.001751158, 
    0.001751155, 0.001751166, 0.001751161, 0.001751175, 0.001751172, 
    0.001751173, 0.001751175, 0.00175117, 0.001751164, 0.001751164, 
    0.001751162, 0.001751157, 0.001751166, 0.001751139, 0.001751155, 
    0.001751181, 0.001751175, 0.001751175, 0.001751177, 0.001751163, 
    0.001751168, 0.001751155, 0.001751158, 0.001751153, 0.001751155, 
    0.001751156, 0.00175116, 0.001751162, 0.001751168, 0.001751172, 
    0.001751176, 0.001751175, 0.001751171, 0.001751164, 0.001751157, 
    0.001751158, 0.001751153, 0.001751167, 0.001751161, 0.001751163, 
    0.001751157, 0.00175117, 0.001751159, 0.001751173, 0.001751172, 
    0.001751168, 0.001751161, 0.001751159, 0.001751157, 0.001751158, 
    0.001751164, 0.001751164, 0.001751168, 0.001751169, 0.001751172, 
    0.001751174, 0.001751172, 0.00175117, 0.001751164, 0.001751158, 
    0.001751152, 0.00175115, 0.001751143, 0.001751149, 0.001751139, 
    0.001751147, 0.001751133, 0.001751159, 0.001751147, 0.001751168, 
    0.001751166, 0.001751162, 0.001751153, 0.001751157, 0.001751152, 
    0.001751164, 0.001751171, 0.001751173, 0.001751176, 0.001751173, 
    0.001751173, 0.00175117, 0.001751171, 0.001751163, 0.001751167, 
    0.001751156, 0.001751152, 0.00175114, 0.001751133, 0.001751125, 
    0.001751122, 0.001751121, 0.001751121,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.733029e-07, 9.732992e-07, 9.732998e-07, 9.732968e-07, 9.732985e-07, 
    9.732966e-07, 9.733021e-07, 9.732989e-07, 9.73301e-07, 9.733026e-07, 
    9.73291e-07, 9.732967e-07, 9.732851e-07, 9.732887e-07, 9.732796e-07, 
    9.732856e-07, 9.732784e-07, 9.732797e-07, 9.732755e-07, 9.732768e-07, 
    9.732714e-07, 9.73275e-07, 9.732686e-07, 9.732722e-07, 9.732717e-07, 
    9.732751e-07, 9.732955e-07, 9.732917e-07, 9.732958e-07, 9.732952e-07, 
    9.732955e-07, 9.732985e-07, 9.733e-07, 9.733031e-07, 9.733026e-07, 
    9.733003e-07, 9.73295e-07, 9.732968e-07, 9.732922e-07, 9.732923e-07, 
    9.732873e-07, 9.732896e-07, 9.732812e-07, 9.732836e-07, 9.732767e-07, 
    9.732785e-07, 9.732768e-07, 9.732772e-07, 9.732768e-07, 9.732793e-07, 
    9.732782e-07, 9.732804e-07, 9.732892e-07, 9.732867e-07, 9.732943e-07, 
    9.732989e-07, 9.73302e-07, 9.733042e-07, 9.733038e-07, 9.733033e-07, 
    9.733002e-07, 9.732973e-07, 9.732952e-07, 9.732938e-07, 9.732923e-07, 
    9.732881e-07, 9.732858e-07, 9.732807e-07, 9.732817e-07, 9.732801e-07, 
    9.732786e-07, 9.732761e-07, 9.732765e-07, 9.732754e-07, 9.732802e-07, 
    9.73277e-07, 9.732821e-07, 9.732807e-07, 9.73292e-07, 9.732963e-07, 
    9.732981e-07, 9.732997e-07, 9.733036e-07, 9.733009e-07, 9.73302e-07, 
    9.732995e-07, 9.732978e-07, 9.732986e-07, 9.732937e-07, 9.732956e-07, 
    9.732856e-07, 9.7329e-07, 9.732788e-07, 9.732814e-07, 9.732781e-07, 
    9.732798e-07, 9.732769e-07, 9.732795e-07, 9.732751e-07, 9.73274e-07, 
    9.732747e-07, 9.732721e-07, 9.732797e-07, 9.732768e-07, 9.732987e-07, 
    9.732985e-07, 9.732979e-07, 9.733005e-07, 9.733008e-07, 9.733031e-07, 
    9.73301e-07, 9.733001e-07, 9.732978e-07, 9.732964e-07, 9.732951e-07, 
    9.732922e-07, 9.732889e-07, 9.732845e-07, 9.732813e-07, 9.732792e-07, 
    9.732804e-07, 9.732793e-07, 9.732806e-07, 9.732812e-07, 9.732744e-07, 
    9.732782e-07, 9.732724e-07, 9.732728e-07, 9.732754e-07, 9.732728e-07, 
    9.732985e-07, 9.732992e-07, 9.733018e-07, 9.732997e-07, 9.733035e-07, 
    9.733013e-07, 9.733002e-07, 9.732956e-07, 9.732946e-07, 9.732937e-07, 
    9.732919e-07, 9.732895e-07, 9.732854e-07, 9.732818e-07, 9.732785e-07, 
    9.732787e-07, 9.732787e-07, 9.732779e-07, 9.732797e-07, 9.732777e-07, 
    9.732773e-07, 9.732782e-07, 9.732729e-07, 9.732744e-07, 9.732728e-07, 
    9.732738e-07, 9.732989e-07, 9.732977e-07, 9.732984e-07, 9.732971e-07, 
    9.73298e-07, 9.73294e-07, 9.732928e-07, 9.732872e-07, 9.732895e-07, 
    9.732859e-07, 9.732892e-07, 9.732886e-07, 9.732858e-07, 9.73289e-07, 
    9.73282e-07, 9.732868e-07, 9.732779e-07, 9.732827e-07, 9.732776e-07, 
    9.732785e-07, 9.73277e-07, 9.732756e-07, 9.732739e-07, 9.732709e-07, 
    9.732715e-07, 9.732689e-07, 9.732959e-07, 9.732942e-07, 9.732944e-07, 
    9.732927e-07, 9.732914e-07, 9.732887e-07, 9.732844e-07, 9.73286e-07, 
    9.73283e-07, 9.732823e-07, 9.732869e-07, 9.732842e-07, 9.732931e-07, 
    9.732917e-07, 9.732926e-07, 9.732958e-07, 9.732856e-07, 9.732908e-07, 
    9.732812e-07, 9.73284e-07, 9.732759e-07, 9.7328e-07, 9.73272e-07, 
    9.732686e-07, 9.732653e-07, 9.732616e-07, 9.732934e-07, 9.732944e-07, 
    9.732925e-07, 9.732897e-07, 9.732872e-07, 9.732838e-07, 9.732835e-07, 
    9.732829e-07, 9.732812e-07, 9.732798e-07, 9.732827e-07, 9.732795e-07, 
    9.732913e-07, 9.732852e-07, 9.732948e-07, 9.732919e-07, 9.732898e-07, 
    9.732908e-07, 9.732862e-07, 9.732851e-07, 9.732806e-07, 9.732829e-07, 
    9.732694e-07, 9.732754e-07, 9.732588e-07, 9.732634e-07, 9.732948e-07, 
    9.732934e-07, 9.732881e-07, 9.732906e-07, 9.732836e-07, 9.732819e-07, 
    9.732805e-07, 9.732787e-07, 9.732785e-07, 9.732775e-07, 9.732792e-07, 
    9.732776e-07, 9.732838e-07, 9.73281e-07, 9.732888e-07, 9.732869e-07, 
    9.732878e-07, 9.732887e-07, 9.732858e-07, 9.732827e-07, 9.732826e-07, 
    9.732815e-07, 9.732787e-07, 9.732836e-07, 9.732686e-07, 9.732779e-07, 
    9.732917e-07, 9.732888e-07, 9.732885e-07, 9.732896e-07, 9.732821e-07, 
    9.732848e-07, 9.732775e-07, 9.732795e-07, 9.732762e-07, 9.732778e-07, 
    9.732781e-07, 9.732802e-07, 9.732814e-07, 9.732846e-07, 9.732873e-07, 
    9.732894e-07, 9.732889e-07, 9.732867e-07, 9.732825e-07, 9.732785e-07, 
    9.732794e-07, 9.732764e-07, 9.732842e-07, 9.73281e-07, 9.732821e-07, 
    9.732789e-07, 9.73286e-07, 9.7328e-07, 9.732876e-07, 9.732869e-07, 
    9.732848e-07, 9.732807e-07, 9.732798e-07, 9.732788e-07, 9.732794e-07, 
    9.732823e-07, 9.732828e-07, 9.732848e-07, 9.732855e-07, 9.73287e-07, 
    9.732884e-07, 9.732871e-07, 9.732859e-07, 9.732823e-07, 9.732792e-07, 
    9.732756e-07, 9.732748e-07, 9.732707e-07, 9.73274e-07, 9.732686e-07, 
    9.732732e-07, 9.732652e-07, 9.732796e-07, 9.732734e-07, 9.732847e-07, 
    9.732835e-07, 9.732813e-07, 9.732762e-07, 9.732789e-07, 9.732757e-07, 
    9.732828e-07, 9.732865e-07, 9.732875e-07, 9.732893e-07, 9.732875e-07, 
    9.732876e-07, 9.732859e-07, 9.732864e-07, 9.732822e-07, 9.732845e-07, 
    9.732781e-07, 9.732757e-07, 9.732692e-07, 9.732652e-07, 9.732611e-07, 
    9.732593e-07, 9.732587e-07, 9.732585e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  6.715481e-25, 2.156797e-25, -5.490028e-25, 6.764499e-25, -7.401734e-25, 
    6.862535e-26, 2.254833e-25, 1.862688e-25, -1.372507e-25, -5.588064e-25, 
    1.764652e-25, -1.960724e-25, 3.823413e-25, 3.529304e-25, 3.061136e-41, 
    3.061136e-41, -5.19592e-25, 2.745014e-25, -2.156797e-25, -2.843051e-25, 
    -1.176435e-25, 1.176435e-24, -1.024478e-24, 2.058761e-25, -1.960724e-26, 
    4.901811e-26, -1.156827e-24, -3.061136e-41, 8.431115e-25, -2.941087e-25, 
    -5.19592e-25, 8.82326e-25, -6.372354e-26, 1.470543e-26, -1.862688e-25, 
    9.117368e-25, 3.088141e-25, 3.823413e-25, 3.137159e-25, 6.078246e-25, 
    6.323336e-25, 2.646978e-25, 7.842898e-26, 1.470543e-25, 9.313441e-25, 
    6.568427e-25, -1.666616e-25, 1.122515e-24, 4.264576e-25, 7.156644e-25, 
    5.146902e-25, -3.872431e-25, 6.715481e-25, -6.862535e-25, 1.372507e-25, 
    3.088141e-25, 5.19592e-25, 7.842898e-26, 6.862535e-26, 6.47039e-25, 
    -1.960724e-25, -7.058608e-25, 3.529304e-25, 3.137159e-25, -5.882173e-25, 
    -2.058761e-25, 3.872431e-25, 6.421373e-25, 5.244938e-25, 1.764652e-25, 
    5.490028e-25, -1.078398e-25, 4.019485e-25, -4.901811e-25, 5.882173e-26, 
    5.391992e-25, -1.862688e-25, -1.911706e-25, 6.764499e-25, 4.901811e-26, 
    -1.764652e-25, -7.352717e-25, 3.431268e-25, 2.450905e-26, 6.715481e-25, 
    -6.862535e-26, 6.078246e-25, 1.960724e-25, 6.813517e-25, -2.058761e-25, 
    -1.81367e-25, -1.960724e-26, 2.254833e-25, 5.735119e-25, 4.901811e-26, 
    -3.333231e-25, 5.882173e-26, 5.784137e-25, 6.862535e-26, 3.921449e-26, 
    3.480286e-25, -9.803622e-27, -2.352869e-25, 1.333293e-24, 2.646978e-25, 
    -1.56858e-25, 6.372354e-25, -4.901811e-26, 4.607703e-25, 7.548789e-25, 
    -9.803622e-26, -3.431268e-26, -2.352869e-25, 5.882173e-26, 1.098006e-24, 
    1.960724e-26, 1.56858e-25, -1.715634e-25, 5.097883e-25, -3.480286e-25, 
    7.25468e-25, -1.470543e-25, 1.078398e-25, 1.666616e-25, 3.725376e-25, 
    2.548942e-25, 2.058761e-25, 4.607703e-25, 3.431268e-26, 2.646978e-25, 
    -9.313441e-26, 3.529304e-25, 5.735119e-25, -8.186024e-25, -5.490028e-25, 
    1.470543e-25, -6.078246e-25, -2.745014e-25, -3.676358e-25, 4.509666e-25, 
    4.117521e-25, 2.941087e-26, 7.842898e-25, -1.421525e-25, 2.156797e-25, 
    -9.803622e-26, 2.401887e-25, 6.47039e-25, -6.862535e-26, -1.617598e-25, 
    -9.068351e-25, 8.235043e-25, 7.450753e-25, -7.352717e-25, 5.293956e-25, 
    2.941087e-25, 3.725376e-25, 6.274318e-25, 1.274471e-25, 6.323336e-25, 
    2.009742e-25, -5.784137e-25, 5.490028e-25, 5.391992e-25, -2.646978e-25, 
    -2.352869e-25, 1.960724e-26, 7.842898e-26, 2.745014e-25, 1.56858e-25, 
    8.725224e-25, -7.842898e-25, 2.352869e-25, 1.470543e-25, -5.882173e-26, 
    -2.205815e-25, -3.872431e-25, 2.843051e-25, -3.529304e-25, -4.019485e-25, 
    -3.333231e-25, 7.989952e-25, 3.529304e-25, -1.02938e-24, 4.117521e-25, 
    6.372354e-26, 4.901811e-26, -1.117613e-24, 6.666463e-25, 1.666616e-25, 
    9.60755e-25, 3.725376e-25, 3.235195e-25, 7.00959e-25, -3.284213e-25, 
    -8.725224e-25, -5.293956e-25, 8.82326e-25, 5.19592e-25, 1.24506e-24, 
    4.509666e-25, 5.293956e-25, -6.176282e-25, 2.941087e-26, 2.156797e-25, 
    -3.921449e-26, 9.803622e-26, 3.039123e-25, -6.862535e-26, -3.62734e-25, 
    -1.088202e-24, 4.313593e-25, 2.745014e-25, 2.695996e-25, 1.862688e-25, 
    2.59796e-25, -1.911706e-25, 1.176435e-24, 3.431268e-25, -6.274318e-25, 
    1.960724e-25, -4.705739e-25, -2.107779e-25, 1.960724e-25, 1.764652e-25, 
    6.666463e-25, 3.137159e-25, -2.941087e-25, 8.431115e-25, 4.362612e-25, 
    -4.313593e-25, 4.41163e-25, 7.352717e-25, 3.186177e-25, 4.901811e-26, 
    1.666616e-25, 7.058608e-25, -1.960724e-25, 9.460495e-25, -2.107779e-25, 
    -1.56858e-25, 7.744861e-25, -1.470543e-25, -6.568427e-25, 1.372507e-25, 
    5.686101e-25, 1.470543e-25, -2.205815e-25, 3.823413e-25, -9.313441e-25, 
    -1.176435e-25, 3.921449e-26, 4.901811e-26, -8.82326e-26, 1.666616e-25, 
    -3.921449e-26, -2.548942e-25, -2.107779e-25, 6.862535e-26, 1.176435e-25, 
    4.901811e-25, -1.960724e-25, -4.803775e-25, 3.62734e-25, 6.078246e-25, 
    -2.843051e-25, -1.421525e-25, -6.078246e-25, -2.303851e-25, 6.862535e-26, 
    1.078398e-25, 3.921449e-26, -1.666616e-25, -9.803622e-26, -6.862535e-26, 
    2.646978e-25, 2.107779e-25, -2.254833e-25, 2.745014e-25, 2.450905e-26, 
    1.862688e-25, 5.98021e-25, 2.695996e-25, 5.882173e-25, -2.941087e-26, 
    7.450753e-25, 7.842898e-26, -4.901811e-26, -1.078398e-24, 1.470543e-26, 
    3.137159e-25, -1.215649e-24, 8.137007e-25, -1.078398e-25, 1.372507e-25, 
    -3.333231e-25, -4.313593e-25, 7.352717e-26, -1.960724e-25, -3.431268e-25, 
    -5.391992e-25, -2.156797e-25, 1.666616e-25, -4.509666e-25, 4.313593e-25, 
    -4.901811e-25, -2.646978e-25, 1.343096e-24, 5.293956e-25, -4.950829e-25, 
    9.362459e-25, 6.960572e-25, 3.235195e-25, -1.715634e-25, -8.82326e-26, 
    -7.842898e-26, 3.62734e-25, 5.735119e-25, -3.137159e-25, 4.803775e-25, 
    -6.862535e-26, -9.411477e-25, 2.548942e-25, 5.833155e-25, -8.82326e-26, 
    -2.058761e-25, 4.362612e-25, -9.803622e-27, -5.391992e-26, -1.862688e-25, 
    4.803775e-25, 6.372354e-25, 4.803775e-25, 2.843051e-25, 2.401887e-25, 
    -4.117521e-25, 6.274318e-25, -8.431115e-25,
  9.436869e-32, 9.436832e-32, 9.436839e-32, 9.436809e-32, 9.436825e-32, 
    9.436806e-32, 9.436862e-32, 9.43683e-32, 9.43685e-32, 9.436866e-32, 
    9.43675e-32, 9.436807e-32, 9.43669e-32, 9.436727e-32, 9.436635e-32, 
    9.436696e-32, 9.436623e-32, 9.436637e-32, 9.436595e-32, 9.436607e-32, 
    9.436553e-32, 9.436589e-32, 9.436525e-32, 9.436561e-32, 9.436556e-32, 
    9.43659e-32, 9.436796e-32, 9.436757e-32, 9.436798e-32, 9.436792e-32, 
    9.436795e-32, 9.436825e-32, 9.43684e-32, 9.436872e-32, 9.436866e-32, 
    9.436843e-32, 9.43679e-32, 9.436808e-32, 9.436763e-32, 9.436763e-32, 
    9.436713e-32, 9.436736e-32, 9.436652e-32, 9.436675e-32, 9.436606e-32, 
    9.436624e-32, 9.436607e-32, 9.436612e-32, 9.436607e-32, 9.436632e-32, 
    9.436622e-32, 9.436644e-32, 9.436732e-32, 9.436706e-32, 9.436783e-32, 
    9.436829e-32, 9.43686e-32, 9.436882e-32, 9.436879e-32, 9.436873e-32, 
    9.436843e-32, 9.436814e-32, 9.436792e-32, 9.436778e-32, 9.436764e-32, 
    9.436721e-32, 9.436698e-32, 9.436646e-32, 9.436656e-32, 9.43664e-32, 
    9.436625e-32, 9.4366e-32, 9.436604e-32, 9.436594e-32, 9.436641e-32, 
    9.436609e-32, 9.436661e-32, 9.436647e-32, 9.43676e-32, 9.436803e-32, 
    9.436822e-32, 9.436837e-32, 9.436876e-32, 9.436849e-32, 9.43686e-32, 
    9.436835e-32, 9.436819e-32, 9.436827e-32, 9.436778e-32, 9.436797e-32, 
    9.436696e-32, 9.436739e-32, 9.436627e-32, 9.436654e-32, 9.436621e-32, 
    9.436638e-32, 9.436608e-32, 9.436635e-32, 9.436589e-32, 9.436579e-32, 
    9.436586e-32, 9.43656e-32, 9.436636e-32, 9.436607e-32, 9.436827e-32, 
    9.436826e-32, 9.43682e-32, 9.436846e-32, 9.436848e-32, 9.436872e-32, 
    9.43685e-32, 9.436841e-32, 9.436818e-32, 9.436804e-32, 9.436791e-32, 
    9.436762e-32, 9.436729e-32, 9.436685e-32, 9.436652e-32, 9.436631e-32, 
    9.436644e-32, 9.436632e-32, 9.436645e-32, 9.436651e-32, 9.436583e-32, 
    9.436621e-32, 9.436564e-32, 9.436567e-32, 9.436593e-32, 9.436567e-32, 
    9.436825e-32, 9.436832e-32, 9.436858e-32, 9.436838e-32, 9.436875e-32, 
    9.436854e-32, 9.436842e-32, 9.436796e-32, 9.436786e-32, 9.436777e-32, 
    9.436759e-32, 9.436735e-32, 9.436693e-32, 9.436657e-32, 9.436625e-32, 
    9.436627e-32, 9.436626e-32, 9.436619e-32, 9.436637e-32, 9.436616e-32, 
    9.436612e-32, 9.436621e-32, 9.436568e-32, 9.436583e-32, 9.436567e-32, 
    9.436577e-32, 9.43683e-32, 9.436817e-32, 9.436824e-32, 9.436811e-32, 
    9.43682e-32, 9.43678e-32, 9.436768e-32, 9.436712e-32, 9.436735e-32, 
    9.436699e-32, 9.436732e-32, 9.436726e-32, 9.436698e-32, 9.43673e-32, 
    9.436659e-32, 9.436707e-32, 9.436618e-32, 9.436666e-32, 9.436615e-32, 
    9.436625e-32, 9.436609e-32, 9.436596e-32, 9.436579e-32, 9.436547e-32, 
    9.436554e-32, 9.436528e-32, 9.436799e-32, 9.436782e-32, 9.436783e-32, 
    9.436766e-32, 9.436754e-32, 9.436727e-32, 9.436683e-32, 9.436699e-32, 
    9.436669e-32, 9.436664e-32, 9.436709e-32, 9.436681e-32, 9.436771e-32, 
    9.436757e-32, 9.436765e-32, 9.436797e-32, 9.436696e-32, 9.436748e-32, 
    9.436652e-32, 9.43668e-32, 9.436598e-32, 9.436638e-32, 9.436558e-32, 
    9.436524e-32, 9.436492e-32, 9.436455e-32, 9.436773e-32, 9.436785e-32, 
    9.436765e-32, 9.436737e-32, 9.436712e-32, 9.436678e-32, 9.436675e-32, 
    9.436668e-32, 9.436652e-32, 9.436638e-32, 9.436666e-32, 9.436635e-32, 
    9.436753e-32, 9.436691e-32, 9.436789e-32, 9.436759e-32, 9.436739e-32, 
    9.436748e-32, 9.436701e-32, 9.436691e-32, 9.436646e-32, 9.436669e-32, 
    9.436532e-32, 9.436593e-32, 9.436426e-32, 9.436473e-32, 9.436788e-32, 
    9.436773e-32, 9.436722e-32, 9.436746e-32, 9.436676e-32, 9.436659e-32, 
    9.436645e-32, 9.436626e-32, 9.436625e-32, 9.436614e-32, 9.436631e-32, 
    9.436615e-32, 9.436678e-32, 9.436649e-32, 9.436728e-32, 9.436709e-32, 
    9.436717e-32, 9.436727e-32, 9.436698e-32, 9.436666e-32, 9.436665e-32, 
    9.436655e-32, 9.436627e-32, 9.436676e-32, 9.436525e-32, 9.436618e-32, 
    9.436757e-32, 9.436729e-32, 9.436725e-32, 9.436735e-32, 9.436661e-32, 
    9.436688e-32, 9.436614e-32, 9.436634e-32, 9.436602e-32, 9.436618e-32, 
    9.43662e-32, 9.436641e-32, 9.436654e-32, 9.436686e-32, 9.436713e-32, 
    9.436734e-32, 9.436729e-32, 9.436706e-32, 9.436664e-32, 9.436625e-32, 
    9.436633e-32, 9.436604e-32, 9.436681e-32, 9.436649e-32, 9.436661e-32, 
    9.436629e-32, 9.4367e-32, 9.436639e-32, 9.436715e-32, 9.436709e-32, 
    9.436688e-32, 9.436646e-32, 9.436637e-32, 9.436628e-32, 9.436634e-32, 
    9.436663e-32, 9.436668e-32, 9.436689e-32, 9.436694e-32, 9.43671e-32, 
    9.436723e-32, 9.436711e-32, 9.436699e-32, 9.436663e-32, 9.436631e-32, 
    9.436595e-32, 9.436587e-32, 9.436546e-32, 9.436579e-32, 9.436524e-32, 
    9.436571e-32, 9.43649e-32, 9.436636e-32, 9.436572e-32, 9.436687e-32, 
    9.436675e-32, 9.436652e-32, 9.436601e-32, 9.436629e-32, 9.436597e-32, 
    9.436668e-32, 9.436705e-32, 9.436715e-32, 9.436733e-32, 9.436714e-32, 
    9.436716e-32, 9.436698e-32, 9.436704e-32, 9.436662e-32, 9.436684e-32, 
    9.43662e-32, 9.436597e-32, 9.436531e-32, 9.43649e-32, 9.43645e-32, 
    9.436431e-32, 9.436425e-32, 9.436424e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.533999e-14, 4.546242e-14, 4.543864e-14, 4.553729e-14, 4.548259e-14, 
    4.554716e-14, 4.536483e-14, 4.546726e-14, 4.540189e-14, 4.535104e-14, 
    4.572844e-14, 4.554169e-14, 4.592225e-14, 4.580336e-14, 4.61018e-14, 
    4.590373e-14, 4.61417e-14, 4.609613e-14, 4.623332e-14, 4.619404e-14, 
    4.636924e-14, 4.625144e-14, 4.646e-14, 4.634114e-14, 4.635973e-14, 
    4.624755e-14, 4.557933e-14, 4.57052e-14, 4.557186e-14, 4.558982e-14, 
    4.558177e-14, 4.54837e-14, 4.543423e-14, 4.533065e-14, 4.534947e-14, 
    4.542555e-14, 4.55979e-14, 4.553945e-14, 4.568677e-14, 4.568344e-14, 
    4.584721e-14, 4.57734e-14, 4.604831e-14, 4.597025e-14, 4.619568e-14, 
    4.613902e-14, 4.619301e-14, 4.617665e-14, 4.619322e-14, 4.611013e-14, 
    4.614573e-14, 4.60726e-14, 4.578722e-14, 4.587116e-14, 4.562061e-14, 
    4.546963e-14, 4.536932e-14, 4.529807e-14, 4.530814e-14, 4.532734e-14, 
    4.5426e-14, 4.551871e-14, 4.55893e-14, 4.563649e-14, 4.568297e-14, 
    4.582345e-14, 4.589781e-14, 4.606406e-14, 4.603411e-14, 4.608487e-14, 
    4.613339e-14, 4.621475e-14, 4.620137e-14, 4.623719e-14, 4.608356e-14, 
    4.618568e-14, 4.601704e-14, 4.606318e-14, 4.569548e-14, 4.555522e-14, 
    4.549545e-14, 4.54432e-14, 4.531589e-14, 4.540382e-14, 4.536916e-14, 
    4.545162e-14, 4.550397e-14, 4.547809e-14, 4.563778e-14, 4.557572e-14, 
    4.590221e-14, 4.57617e-14, 4.612773e-14, 4.604026e-14, 4.614869e-14, 
    4.609338e-14, 4.618812e-14, 4.610286e-14, 4.625053e-14, 4.628265e-14, 
    4.62607e-14, 4.634502e-14, 4.609813e-14, 4.6193e-14, 4.547735e-14, 
    4.548158e-14, 4.550125e-14, 4.541473e-14, 4.540944e-14, 4.533013e-14, 
    4.540072e-14, 4.543075e-14, 4.550701e-14, 4.555207e-14, 4.55949e-14, 
    4.5689e-14, 4.579399e-14, 4.594066e-14, 4.604593e-14, 4.611643e-14, 
    4.607322e-14, 4.611137e-14, 4.606871e-14, 4.604872e-14, 4.62706e-14, 
    4.614606e-14, 4.63329e-14, 4.632257e-14, 4.623804e-14, 4.632373e-14, 
    4.548454e-14, 4.546025e-14, 4.537582e-14, 4.544189e-14, 4.532149e-14, 
    4.538889e-14, 4.542761e-14, 4.557699e-14, 4.560981e-14, 4.56402e-14, 
    4.570021e-14, 4.577718e-14, 4.591205e-14, 4.602929e-14, 4.613621e-14, 
    4.612839e-14, 4.613114e-14, 4.6155e-14, 4.609587e-14, 4.616471e-14, 
    4.617625e-14, 4.614606e-14, 4.632119e-14, 4.627119e-14, 4.632235e-14, 
    4.62898e-14, 4.546815e-14, 4.550903e-14, 4.548694e-14, 4.552846e-14, 
    4.54992e-14, 4.562924e-14, 4.56682e-14, 4.585034e-14, 4.577566e-14, 
    4.589453e-14, 4.578775e-14, 4.580667e-14, 4.589835e-14, 4.579353e-14, 
    4.60228e-14, 4.586737e-14, 4.615593e-14, 4.600086e-14, 4.616564e-14, 
    4.613575e-14, 4.618524e-14, 4.622953e-14, 4.628524e-14, 4.638792e-14, 
    4.636416e-14, 4.644999e-14, 4.556996e-14, 4.562292e-14, 4.561828e-14, 
    4.567369e-14, 4.571465e-14, 4.580341e-14, 4.594558e-14, 4.589215e-14, 
    4.599025e-14, 4.600993e-14, 4.586089e-14, 4.59524e-14, 4.565837e-14, 
    4.57059e-14, 4.567762e-14, 4.557412e-14, 4.590444e-14, 4.573503e-14, 
    4.604767e-14, 4.595605e-14, 4.622321e-14, 4.609041e-14, 4.635107e-14, 
    4.646224e-14, 4.656686e-14, 4.668886e-14, 4.565183e-14, 4.561586e-14, 
    4.568029e-14, 4.576933e-14, 4.585194e-14, 4.596164e-14, 4.597287e-14, 
    4.59934e-14, 4.604658e-14, 4.609127e-14, 4.599987e-14, 4.610247e-14, 
    4.571688e-14, 4.591914e-14, 4.560223e-14, 4.569773e-14, 4.576409e-14, 
    4.573501e-14, 4.588605e-14, 4.592161e-14, 4.606598e-14, 4.599139e-14, 
    4.643479e-14, 4.623885e-14, 4.678173e-14, 4.66303e-14, 4.560328e-14, 
    4.565172e-14, 4.582012e-14, 4.574003e-14, 4.596897e-14, 4.602524e-14, 
    4.607098e-14, 4.612938e-14, 4.61357e-14, 4.617029e-14, 4.61136e-14, 
    4.616806e-14, 4.596187e-14, 4.605407e-14, 4.580091e-14, 4.586257e-14, 
    4.583422e-14, 4.580309e-14, 4.589912e-14, 4.60013e-14, 4.600352e-14, 
    4.603625e-14, 4.612838e-14, 4.59699e-14, 4.645998e-14, 4.615753e-14, 
    4.570452e-14, 4.579767e-14, 4.581101e-14, 4.577493e-14, 4.601959e-14, 
    4.593101e-14, 4.616945e-14, 4.610507e-14, 4.621055e-14, 4.615814e-14, 
    4.615043e-14, 4.608309e-14, 4.604113e-14, 4.593506e-14, 4.584869e-14, 
    4.578017e-14, 4.579611e-14, 4.587137e-14, 4.600755e-14, 4.613625e-14, 
    4.610807e-14, 4.620254e-14, 4.595238e-14, 4.605733e-14, 4.601677e-14, 
    4.612251e-14, 4.589072e-14, 4.608802e-14, 4.584022e-14, 4.586198e-14, 
    4.592925e-14, 4.606442e-14, 4.609436e-14, 4.612625e-14, 4.610658e-14, 
    4.601102e-14, 4.599537e-14, 4.592762e-14, 4.590889e-14, 4.585724e-14, 
    4.581445e-14, 4.585354e-14, 4.589457e-14, 4.601107e-14, 4.611593e-14, 
    4.623015e-14, 4.62581e-14, 4.639127e-14, 4.628283e-14, 4.646166e-14, 
    4.630956e-14, 4.657275e-14, 4.60995e-14, 4.630516e-14, 4.593232e-14, 
    4.597256e-14, 4.604526e-14, 4.62119e-14, 4.612201e-14, 4.622715e-14, 
    4.599476e-14, 4.587395e-14, 4.584271e-14, 4.578433e-14, 4.584404e-14, 
    4.583919e-14, 4.589629e-14, 4.587795e-14, 4.601494e-14, 4.594138e-14, 
    4.615023e-14, 4.622633e-14, 4.644098e-14, 4.657233e-14, 4.670591e-14, 
    4.676481e-14, 4.678273e-14, 4.679022e-14 ;

 LITR1N_vr =
  5.55766e-05, 5.557639e-05, 5.557643e-05, 5.557626e-05, 5.557635e-05, 
    5.557624e-05, 5.557655e-05, 5.557638e-05, 5.557649e-05, 5.557658e-05, 
    5.557592e-05, 5.557625e-05, 5.557558e-05, 5.557579e-05, 5.557527e-05, 
    5.557562e-05, 5.55752e-05, 5.557528e-05, 5.557504e-05, 5.557511e-05, 
    5.55748e-05, 5.557501e-05, 5.557464e-05, 5.557485e-05, 5.557482e-05, 
    5.557502e-05, 5.557618e-05, 5.557596e-05, 5.557619e-05, 5.557616e-05, 
    5.557618e-05, 5.557635e-05, 5.557643e-05, 5.557662e-05, 5.557658e-05, 
    5.557645e-05, 5.557615e-05, 5.557625e-05, 5.557599e-05, 5.5576e-05, 
    5.557571e-05, 5.557584e-05, 5.557536e-05, 5.55755e-05, 5.557511e-05, 
    5.55752e-05, 5.557511e-05, 5.557514e-05, 5.557511e-05, 5.557526e-05, 
    5.557519e-05, 5.557532e-05, 5.557582e-05, 5.557567e-05, 5.557611e-05, 
    5.557637e-05, 5.557655e-05, 5.557667e-05, 5.557666e-05, 5.557662e-05, 
    5.557645e-05, 5.557629e-05, 5.557617e-05, 5.557608e-05, 5.5576e-05, 
    5.557575e-05, 5.557563e-05, 5.557534e-05, 5.557539e-05, 5.55753e-05, 
    5.557521e-05, 5.557507e-05, 5.55751e-05, 5.557503e-05, 5.55753e-05, 
    5.557512e-05, 5.557542e-05, 5.557534e-05, 5.557598e-05, 5.557622e-05, 
    5.557633e-05, 5.557642e-05, 5.557664e-05, 5.557649e-05, 5.557655e-05, 
    5.557641e-05, 5.557631e-05, 5.557636e-05, 5.557608e-05, 5.557619e-05, 
    5.557562e-05, 5.557586e-05, 5.557522e-05, 5.557538e-05, 5.557519e-05, 
    5.557528e-05, 5.557512e-05, 5.557527e-05, 5.557501e-05, 5.557495e-05, 
    5.557499e-05, 5.557484e-05, 5.557527e-05, 5.557511e-05, 5.557636e-05, 
    5.557635e-05, 5.557632e-05, 5.557647e-05, 5.557648e-05, 5.557662e-05, 
    5.557649e-05, 5.557644e-05, 5.557631e-05, 5.557623e-05, 5.557615e-05, 
    5.557599e-05, 5.557581e-05, 5.557555e-05, 5.557536e-05, 5.557524e-05, 
    5.557532e-05, 5.557525e-05, 5.557532e-05, 5.557536e-05, 5.557498e-05, 
    5.557519e-05, 5.557487e-05, 5.557488e-05, 5.557503e-05, 5.557488e-05, 
    5.557635e-05, 5.557639e-05, 5.557654e-05, 5.557642e-05, 5.557663e-05, 
    5.557651e-05, 5.557645e-05, 5.557619e-05, 5.557613e-05, 5.557607e-05, 
    5.557597e-05, 5.557583e-05, 5.55756e-05, 5.557539e-05, 5.557521e-05, 
    5.557522e-05, 5.557522e-05, 5.557518e-05, 5.557528e-05, 5.557516e-05, 
    5.557514e-05, 5.557519e-05, 5.557488e-05, 5.557497e-05, 5.557488e-05, 
    5.557494e-05, 5.557638e-05, 5.55763e-05, 5.557634e-05, 5.557627e-05, 
    5.557632e-05, 5.557609e-05, 5.557603e-05, 5.557571e-05, 5.557584e-05, 
    5.557563e-05, 5.557582e-05, 5.557578e-05, 5.557562e-05, 5.557581e-05, 
    5.557541e-05, 5.557568e-05, 5.557518e-05, 5.557545e-05, 5.557516e-05, 
    5.557521e-05, 5.557512e-05, 5.557504e-05, 5.557495e-05, 5.557477e-05, 
    5.557481e-05, 5.557466e-05, 5.55762e-05, 5.557611e-05, 5.557611e-05, 
    5.557602e-05, 5.557594e-05, 5.557579e-05, 5.557554e-05, 5.557563e-05, 
    5.557546e-05, 5.557543e-05, 5.557569e-05, 5.557553e-05, 5.557605e-05, 
    5.557596e-05, 5.557601e-05, 5.557619e-05, 5.557561e-05, 5.557591e-05, 
    5.557536e-05, 5.557553e-05, 5.557506e-05, 5.557529e-05, 5.557483e-05, 
    5.557464e-05, 5.557446e-05, 5.557424e-05, 5.557606e-05, 5.557612e-05, 
    5.557601e-05, 5.557585e-05, 5.557571e-05, 5.557551e-05, 5.55755e-05, 
    5.557546e-05, 5.557536e-05, 5.557529e-05, 5.557545e-05, 5.557527e-05, 
    5.557594e-05, 5.557559e-05, 5.557614e-05, 5.557598e-05, 5.557586e-05, 
    5.557591e-05, 5.557565e-05, 5.557558e-05, 5.557533e-05, 5.557546e-05, 
    5.557469e-05, 5.557503e-05, 5.557408e-05, 5.557435e-05, 5.557614e-05, 
    5.557606e-05, 5.557576e-05, 5.55759e-05, 5.55755e-05, 5.55754e-05, 
    5.557532e-05, 5.557522e-05, 5.557521e-05, 5.557515e-05, 5.557525e-05, 
    5.557515e-05, 5.557551e-05, 5.557535e-05, 5.557579e-05, 5.557569e-05, 
    5.557574e-05, 5.557579e-05, 5.557562e-05, 5.557545e-05, 5.557544e-05, 
    5.557538e-05, 5.557522e-05, 5.55755e-05, 5.557464e-05, 5.557517e-05, 
    5.557596e-05, 5.55758e-05, 5.557578e-05, 5.557584e-05, 5.557541e-05, 
    5.557557e-05, 5.557515e-05, 5.557526e-05, 5.557508e-05, 5.557517e-05, 
    5.557518e-05, 5.55753e-05, 5.557538e-05, 5.557556e-05, 5.557571e-05, 
    5.557583e-05, 5.55758e-05, 5.557567e-05, 5.557543e-05, 5.557521e-05, 
    5.557526e-05, 5.557509e-05, 5.557553e-05, 5.557535e-05, 5.557542e-05, 
    5.557523e-05, 5.557564e-05, 5.557529e-05, 5.557573e-05, 5.557569e-05, 
    5.557557e-05, 5.557534e-05, 5.557528e-05, 5.557523e-05, 5.557526e-05, 
    5.557543e-05, 5.557546e-05, 5.557557e-05, 5.557561e-05, 5.55757e-05, 
    5.557577e-05, 5.55757e-05, 5.557563e-05, 5.557543e-05, 5.557524e-05, 
    5.557504e-05, 5.5575e-05, 5.557476e-05, 5.557495e-05, 5.557464e-05, 
    5.557491e-05, 5.557444e-05, 5.557527e-05, 5.557491e-05, 5.557557e-05, 
    5.55755e-05, 5.557537e-05, 5.557508e-05, 5.557523e-05, 5.557505e-05, 
    5.557546e-05, 5.557567e-05, 5.557572e-05, 5.557582e-05, 5.557572e-05, 
    5.557573e-05, 5.557563e-05, 5.557566e-05, 5.557542e-05, 5.557555e-05, 
    5.557518e-05, 5.557505e-05, 5.557468e-05, 5.557445e-05, 5.557422e-05, 
    5.557411e-05, 5.557408e-05, 5.557407e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  7.857573e-13, 7.87879e-13, 7.874669e-13, 7.891766e-13, 7.882286e-13, 
    7.893476e-13, 7.86188e-13, 7.87963e-13, 7.868302e-13, 7.859488e-13, 
    7.924893e-13, 7.892529e-13, 7.95848e-13, 7.937878e-13, 7.989598e-13, 
    7.955272e-13, 7.996513e-13, 7.988615e-13, 8.01239e-13, 8.005582e-13, 
    8.035945e-13, 8.015532e-13, 8.051675e-13, 8.031076e-13, 8.034297e-13, 
    8.014857e-13, 7.899053e-13, 7.920865e-13, 7.897758e-13, 7.90087e-13, 
    7.899475e-13, 7.88248e-13, 7.873906e-13, 7.855955e-13, 7.859216e-13, 
    7.872402e-13, 7.90227e-13, 7.89214e-13, 7.917672e-13, 7.917095e-13, 
    7.945476e-13, 7.932685e-13, 7.980327e-13, 7.9668e-13, 8.005867e-13, 
    7.996049e-13, 8.005405e-13, 8.002569e-13, 8.005441e-13, 7.991041e-13, 
    7.997212e-13, 7.984536e-13, 7.93508e-13, 7.949626e-13, 7.906206e-13, 
    7.88004e-13, 7.862657e-13, 7.850308e-13, 7.852054e-13, 7.855381e-13, 
    7.872479e-13, 7.888546e-13, 7.900779e-13, 7.908957e-13, 7.917012e-13, 
    7.941359e-13, 7.954245e-13, 7.983058e-13, 7.977866e-13, 7.986664e-13, 
    7.995072e-13, 8.009173e-13, 8.006853e-13, 8.013062e-13, 7.986436e-13, 
    8.004134e-13, 7.974908e-13, 7.982905e-13, 7.919181e-13, 7.894875e-13, 
    7.884516e-13, 7.875461e-13, 7.853396e-13, 7.868635e-13, 7.862629e-13, 
    7.87692e-13, 7.885992e-13, 7.881506e-13, 7.909181e-13, 7.898425e-13, 
    7.955009e-13, 7.930657e-13, 7.994091e-13, 7.978933e-13, 7.997724e-13, 
    7.988139e-13, 8.004558e-13, 7.989781e-13, 8.015373e-13, 8.020939e-13, 
    8.017135e-13, 8.031749e-13, 7.988962e-13, 8.005402e-13, 7.881379e-13, 
    7.882111e-13, 7.885521e-13, 7.870526e-13, 7.86961e-13, 7.855864e-13, 
    7.868097e-13, 7.873303e-13, 7.886519e-13, 7.894328e-13, 7.90175e-13, 
    7.918059e-13, 7.936253e-13, 7.961672e-13, 7.979916e-13, 7.992133e-13, 
    7.984644e-13, 7.991256e-13, 7.983864e-13, 7.980399e-13, 8.018852e-13, 
    7.997268e-13, 8.029647e-13, 8.027858e-13, 8.013208e-13, 8.02806e-13, 
    7.882625e-13, 7.878414e-13, 7.863782e-13, 7.875234e-13, 7.854367e-13, 
    7.866048e-13, 7.872759e-13, 7.898646e-13, 7.904334e-13, 7.9096e-13, 
    7.920001e-13, 7.933339e-13, 7.956714e-13, 7.977031e-13, 7.995562e-13, 
    7.994205e-13, 7.994683e-13, 7.998818e-13, 7.98857e-13, 8.0005e-13, 
    8.002499e-13, 7.997268e-13, 8.027618e-13, 8.018953e-13, 8.02782e-13, 
    8.022179e-13, 7.879784e-13, 7.886868e-13, 7.88304e-13, 7.890237e-13, 
    7.885166e-13, 7.907701e-13, 7.914453e-13, 7.94602e-13, 7.933076e-13, 
    7.953677e-13, 7.935171e-13, 7.938451e-13, 7.95434e-13, 7.936173e-13, 
    7.975907e-13, 7.94897e-13, 7.998979e-13, 7.972104e-13, 8.000661e-13, 
    7.995482e-13, 8.004058e-13, 8.011733e-13, 8.021388e-13, 8.039183e-13, 
    8.035065e-13, 8.04994e-13, 7.897427e-13, 7.906606e-13, 7.905802e-13, 
    7.915406e-13, 7.922504e-13, 7.937885e-13, 7.962525e-13, 7.953265e-13, 
    7.970266e-13, 7.973676e-13, 7.947848e-13, 7.963706e-13, 7.912749e-13, 
    7.920987e-13, 7.916085e-13, 7.898149e-13, 7.955394e-13, 7.926035e-13, 
    7.980216e-13, 7.964339e-13, 8.010639e-13, 7.987623e-13, 8.032796e-13, 
    8.052063e-13, 8.070194e-13, 8.091338e-13, 7.911617e-13, 7.905382e-13, 
    7.916548e-13, 7.931979e-13, 7.946296e-13, 7.965307e-13, 7.967253e-13, 
    7.970811e-13, 7.980028e-13, 7.987773e-13, 7.971932e-13, 7.989714e-13, 
    7.922889e-13, 7.957941e-13, 7.903021e-13, 7.91957e-13, 7.931071e-13, 
    7.926031e-13, 7.952207e-13, 7.95837e-13, 7.98339e-13, 7.970463e-13, 
    8.047306e-13, 8.013348e-13, 8.107433e-13, 8.081189e-13, 7.903202e-13, 
    7.911598e-13, 7.940781e-13, 7.926902e-13, 7.966578e-13, 7.976329e-13, 
    7.984256e-13, 7.994377e-13, 7.995473e-13, 8.001467e-13, 7.991643e-13, 
    8.001081e-13, 7.965348e-13, 7.981325e-13, 7.937452e-13, 7.948138e-13, 
    7.943225e-13, 7.93783e-13, 7.954473e-13, 7.97218e-13, 7.972565e-13, 
    7.978238e-13, 7.994204e-13, 7.966738e-13, 8.051672e-13, 7.999255e-13, 
    7.920747e-13, 7.936891e-13, 7.939204e-13, 7.932951e-13, 7.975352e-13, 
    7.959998e-13, 8.001322e-13, 7.990165e-13, 8.008444e-13, 7.999362e-13, 
    7.998026e-13, 7.986355e-13, 7.979084e-13, 7.960701e-13, 7.945733e-13, 
    7.933859e-13, 7.936621e-13, 7.949663e-13, 7.973265e-13, 7.995569e-13, 
    7.990684e-13, 8.007056e-13, 7.963703e-13, 7.981891e-13, 7.974862e-13, 
    7.993186e-13, 7.953017e-13, 7.98721e-13, 7.944265e-13, 7.948036e-13, 
    7.959694e-13, 7.983119e-13, 7.988308e-13, 7.993835e-13, 7.990426e-13, 
    7.973865e-13, 7.971153e-13, 7.959412e-13, 7.956166e-13, 7.947215e-13, 
    7.939798e-13, 7.946573e-13, 7.953684e-13, 7.973874e-13, 7.992047e-13, 
    8.011842e-13, 8.016685e-13, 8.039763e-13, 8.02097e-13, 8.051962e-13, 
    8.025603e-13, 8.071215e-13, 7.989198e-13, 8.02484e-13, 7.960226e-13, 
    7.967199e-13, 7.9798e-13, 8.008678e-13, 7.9931e-13, 8.011321e-13, 
    7.971047e-13, 7.95011e-13, 7.944696e-13, 7.93458e-13, 7.944928e-13, 
    7.944086e-13, 7.953983e-13, 7.950804e-13, 7.974544e-13, 7.961796e-13, 
    7.99799e-13, 8.011179e-13, 8.04838e-13, 8.071142e-13, 8.094292e-13, 
    8.1045e-13, 8.107606e-13, 8.108904e-13 ;

 LITR2C =
  1.939607e-05, 1.939605e-05, 1.939605e-05, 1.939604e-05, 1.939605e-05, 
    1.939604e-05, 1.939607e-05, 1.939605e-05, 1.939606e-05, 1.939607e-05, 
    1.939601e-05, 1.939604e-05, 1.939598e-05, 1.939599e-05, 1.939595e-05, 
    1.939598e-05, 1.939594e-05, 1.939595e-05, 1.939593e-05, 1.939593e-05, 
    1.93959e-05, 1.939592e-05, 1.939589e-05, 1.939591e-05, 1.939591e-05, 
    1.939592e-05, 1.939603e-05, 1.939601e-05, 1.939603e-05, 1.939603e-05, 
    1.939603e-05, 1.939605e-05, 1.939605e-05, 1.939607e-05, 1.939607e-05, 
    1.939606e-05, 1.939603e-05, 1.939604e-05, 1.939601e-05, 1.939601e-05, 
    1.939599e-05, 1.9396e-05, 1.939596e-05, 1.939597e-05, 1.939593e-05, 
    1.939594e-05, 1.939593e-05, 1.939593e-05, 1.939593e-05, 1.939595e-05, 
    1.939594e-05, 1.939595e-05, 1.9396e-05, 1.939598e-05, 1.939603e-05, 
    1.939605e-05, 1.939607e-05, 1.939608e-05, 1.939608e-05, 1.939607e-05, 
    1.939606e-05, 1.939604e-05, 1.939603e-05, 1.939602e-05, 1.939601e-05, 
    1.939599e-05, 1.939598e-05, 1.939595e-05, 1.939596e-05, 1.939595e-05, 
    1.939594e-05, 1.939593e-05, 1.939593e-05, 1.939593e-05, 1.939595e-05, 
    1.939593e-05, 1.939596e-05, 1.939595e-05, 1.939601e-05, 1.939603e-05, 
    1.939605e-05, 1.939605e-05, 1.939608e-05, 1.939606e-05, 1.939607e-05, 
    1.939605e-05, 1.939604e-05, 1.939605e-05, 1.939602e-05, 1.939603e-05, 
    1.939598e-05, 1.9396e-05, 1.939594e-05, 1.939596e-05, 1.939594e-05, 
    1.939595e-05, 1.939593e-05, 1.939595e-05, 1.939592e-05, 1.939592e-05, 
    1.939592e-05, 1.939591e-05, 1.939595e-05, 1.939593e-05, 1.939605e-05, 
    1.939605e-05, 1.939604e-05, 1.939606e-05, 1.939606e-05, 1.939607e-05, 
    1.939606e-05, 1.939605e-05, 1.939604e-05, 1.939604e-05, 1.939603e-05, 
    1.939601e-05, 1.9396e-05, 1.939597e-05, 1.939596e-05, 1.939595e-05, 
    1.939595e-05, 1.939595e-05, 1.939595e-05, 1.939596e-05, 1.939592e-05, 
    1.939594e-05, 1.939591e-05, 1.939591e-05, 1.939593e-05, 1.939591e-05, 
    1.939605e-05, 1.939605e-05, 1.939606e-05, 1.939605e-05, 1.939607e-05, 
    1.939606e-05, 1.939606e-05, 1.939603e-05, 1.939603e-05, 1.939602e-05, 
    1.939601e-05, 1.9396e-05, 1.939598e-05, 1.939596e-05, 1.939594e-05, 
    1.939594e-05, 1.939594e-05, 1.939594e-05, 1.939595e-05, 1.939594e-05, 
    1.939593e-05, 1.939594e-05, 1.939591e-05, 1.939592e-05, 1.939591e-05, 
    1.939592e-05, 1.939605e-05, 1.939604e-05, 1.939605e-05, 1.939604e-05, 
    1.939604e-05, 1.939602e-05, 1.939602e-05, 1.939599e-05, 1.9396e-05, 
    1.939598e-05, 1.9396e-05, 1.939599e-05, 1.939598e-05, 1.9396e-05, 
    1.939596e-05, 1.939599e-05, 1.939594e-05, 1.939596e-05, 1.939594e-05, 
    1.939594e-05, 1.939593e-05, 1.939593e-05, 1.939592e-05, 1.93959e-05, 
    1.939591e-05, 1.939589e-05, 1.939603e-05, 1.939602e-05, 1.939603e-05, 
    1.939602e-05, 1.939601e-05, 1.939599e-05, 1.939597e-05, 1.939598e-05, 
    1.939597e-05, 1.939596e-05, 1.939599e-05, 1.939597e-05, 1.939602e-05, 
    1.939601e-05, 1.939602e-05, 1.939603e-05, 1.939598e-05, 1.939601e-05, 
    1.939596e-05, 1.939597e-05, 1.939593e-05, 1.939595e-05, 1.939591e-05, 
    1.939589e-05, 1.939587e-05, 1.939585e-05, 1.939602e-05, 1.939603e-05, 
    1.939601e-05, 1.9396e-05, 1.939599e-05, 1.939597e-05, 1.939597e-05, 
    1.939597e-05, 1.939596e-05, 1.939595e-05, 1.939596e-05, 1.939595e-05, 
    1.939601e-05, 1.939598e-05, 1.939603e-05, 1.939601e-05, 1.9396e-05, 
    1.939601e-05, 1.939598e-05, 1.939598e-05, 1.939595e-05, 1.939597e-05, 
    1.939589e-05, 1.939593e-05, 1.939584e-05, 1.939586e-05, 1.939603e-05, 
    1.939602e-05, 1.939599e-05, 1.939601e-05, 1.939597e-05, 1.939596e-05, 
    1.939595e-05, 1.939594e-05, 1.939594e-05, 1.939594e-05, 1.939595e-05, 
    1.939594e-05, 1.939597e-05, 1.939595e-05, 1.9396e-05, 1.939599e-05, 
    1.939599e-05, 1.939599e-05, 1.939598e-05, 1.939596e-05, 1.939596e-05, 
    1.939596e-05, 1.939594e-05, 1.939597e-05, 1.939589e-05, 1.939594e-05, 
    1.939601e-05, 1.9396e-05, 1.939599e-05, 1.9396e-05, 1.939596e-05, 
    1.939597e-05, 1.939594e-05, 1.939595e-05, 1.939593e-05, 1.939594e-05, 
    1.939594e-05, 1.939595e-05, 1.939596e-05, 1.939597e-05, 1.939599e-05, 
    1.9396e-05, 1.9396e-05, 1.939598e-05, 1.939596e-05, 1.939594e-05, 
    1.939595e-05, 1.939593e-05, 1.939597e-05, 1.939595e-05, 1.939596e-05, 
    1.939594e-05, 1.939598e-05, 1.939595e-05, 1.939599e-05, 1.939599e-05, 
    1.939597e-05, 1.939595e-05, 1.939595e-05, 1.939594e-05, 1.939595e-05, 
    1.939596e-05, 1.939596e-05, 1.939597e-05, 1.939598e-05, 1.939599e-05, 
    1.939599e-05, 1.939599e-05, 1.939598e-05, 1.939596e-05, 1.939595e-05, 
    1.939593e-05, 1.939592e-05, 1.93959e-05, 1.939592e-05, 1.939589e-05, 
    1.939591e-05, 1.939587e-05, 1.939595e-05, 1.939591e-05, 1.939597e-05, 
    1.939597e-05, 1.939596e-05, 1.939593e-05, 1.939594e-05, 1.939593e-05, 
    1.939596e-05, 1.939598e-05, 1.939599e-05, 1.9396e-05, 1.939599e-05, 
    1.939599e-05, 1.939598e-05, 1.939598e-05, 1.939596e-05, 1.939597e-05, 
    1.939594e-05, 1.939593e-05, 1.939589e-05, 1.939587e-05, 1.939585e-05, 
    1.939584e-05, 1.939584e-05, 1.939584e-05 ;

 LITR2C_TO_SOIL1C =
  1.196551e-13, 1.199785e-13, 1.199157e-13, 1.201763e-13, 1.200318e-13, 
    1.202024e-13, 1.197207e-13, 1.199913e-13, 1.198186e-13, 1.196843e-13, 
    1.206813e-13, 1.201879e-13, 1.211933e-13, 1.208792e-13, 1.216676e-13, 
    1.211444e-13, 1.21773e-13, 1.216526e-13, 1.220151e-13, 1.219113e-13, 
    1.223742e-13, 1.22063e-13, 1.226139e-13, 1.222999e-13, 1.22349e-13, 
    1.220527e-13, 1.202874e-13, 1.206199e-13, 1.202676e-13, 1.203151e-13, 
    1.202938e-13, 1.200347e-13, 1.19904e-13, 1.196304e-13, 1.196801e-13, 
    1.198811e-13, 1.203364e-13, 1.20182e-13, 1.205712e-13, 1.205624e-13, 
    1.20995e-13, 1.208e-13, 1.215263e-13, 1.213201e-13, 1.219156e-13, 
    1.21766e-13, 1.219086e-13, 1.218654e-13, 1.219092e-13, 1.216896e-13, 
    1.217837e-13, 1.215905e-13, 1.208366e-13, 1.210583e-13, 1.203964e-13, 
    1.199976e-13, 1.197326e-13, 1.195443e-13, 1.19571e-13, 1.196217e-13, 
    1.198823e-13, 1.201272e-13, 1.203137e-13, 1.204384e-13, 1.205611e-13, 
    1.209323e-13, 1.211287e-13, 1.215679e-13, 1.214888e-13, 1.216229e-13, 
    1.217511e-13, 1.21966e-13, 1.219307e-13, 1.220253e-13, 1.216194e-13, 
    1.218892e-13, 1.214437e-13, 1.215656e-13, 1.205942e-13, 1.202237e-13, 
    1.200658e-13, 1.199277e-13, 1.195914e-13, 1.198237e-13, 1.197321e-13, 
    1.1995e-13, 1.200883e-13, 1.200199e-13, 1.204418e-13, 1.202778e-13, 
    1.211403e-13, 1.207691e-13, 1.217361e-13, 1.21505e-13, 1.217915e-13, 
    1.216454e-13, 1.218957e-13, 1.216704e-13, 1.220606e-13, 1.221454e-13, 
    1.220874e-13, 1.223102e-13, 1.216579e-13, 1.219086e-13, 1.20018e-13, 
    1.200291e-13, 1.200811e-13, 1.198525e-13, 1.198386e-13, 1.19629e-13, 
    1.198155e-13, 1.198948e-13, 1.200963e-13, 1.202153e-13, 1.203285e-13, 
    1.205771e-13, 1.208544e-13, 1.212419e-13, 1.2152e-13, 1.217063e-13, 
    1.215921e-13, 1.216929e-13, 1.215802e-13, 1.215274e-13, 1.221136e-13, 
    1.217846e-13, 1.222782e-13, 1.222509e-13, 1.220276e-13, 1.222539e-13, 
    1.20037e-13, 1.199728e-13, 1.197497e-13, 1.199243e-13, 1.196062e-13, 
    1.197843e-13, 1.198866e-13, 1.202812e-13, 1.203679e-13, 1.204482e-13, 
    1.206067e-13, 1.2081e-13, 1.211663e-13, 1.214761e-13, 1.217585e-13, 
    1.217379e-13, 1.217451e-13, 1.218082e-13, 1.21652e-13, 1.218338e-13, 
    1.218643e-13, 1.217846e-13, 1.222472e-13, 1.221151e-13, 1.222503e-13, 
    1.221643e-13, 1.199936e-13, 1.201016e-13, 1.200433e-13, 1.20153e-13, 
    1.200757e-13, 1.204192e-13, 1.205221e-13, 1.210033e-13, 1.20806e-13, 
    1.211201e-13, 1.20838e-13, 1.208879e-13, 1.211302e-13, 1.208532e-13, 
    1.214589e-13, 1.210483e-13, 1.218106e-13, 1.214009e-13, 1.218363e-13, 
    1.217573e-13, 1.218881e-13, 1.220051e-13, 1.221522e-13, 1.224235e-13, 
    1.223607e-13, 1.225875e-13, 1.202626e-13, 1.204025e-13, 1.203902e-13, 
    1.205367e-13, 1.206449e-13, 1.208793e-13, 1.212549e-13, 1.211138e-13, 
    1.213729e-13, 1.214249e-13, 1.210312e-13, 1.212729e-13, 1.204962e-13, 
    1.206217e-13, 1.20547e-13, 1.202736e-13, 1.211462e-13, 1.206987e-13, 
    1.215246e-13, 1.212826e-13, 1.219884e-13, 1.216375e-13, 1.223262e-13, 
    1.226199e-13, 1.228963e-13, 1.232186e-13, 1.204789e-13, 1.203839e-13, 
    1.205541e-13, 1.207893e-13, 1.210075e-13, 1.212973e-13, 1.21327e-13, 
    1.213812e-13, 1.215218e-13, 1.216398e-13, 1.213983e-13, 1.216694e-13, 
    1.206507e-13, 1.211851e-13, 1.203479e-13, 1.206001e-13, 1.207755e-13, 
    1.206986e-13, 1.210976e-13, 1.211916e-13, 1.21573e-13, 1.213759e-13, 
    1.225473e-13, 1.220297e-13, 1.234639e-13, 1.230639e-13, 1.203506e-13, 
    1.204786e-13, 1.209235e-13, 1.207119e-13, 1.213167e-13, 1.214654e-13, 
    1.215862e-13, 1.217405e-13, 1.217572e-13, 1.218486e-13, 1.216988e-13, 
    1.218427e-13, 1.21298e-13, 1.215415e-13, 1.208727e-13, 1.210356e-13, 
    1.209607e-13, 1.208785e-13, 1.211322e-13, 1.214021e-13, 1.21408e-13, 
    1.214945e-13, 1.217379e-13, 1.213192e-13, 1.226139e-13, 1.218148e-13, 
    1.206181e-13, 1.208642e-13, 1.208994e-13, 1.208041e-13, 1.214505e-13, 
    1.212164e-13, 1.218464e-13, 1.216763e-13, 1.219549e-13, 1.218165e-13, 
    1.217961e-13, 1.216182e-13, 1.215074e-13, 1.212271e-13, 1.20999e-13, 
    1.208179e-13, 1.208601e-13, 1.210589e-13, 1.214186e-13, 1.217587e-13, 
    1.216842e-13, 1.219338e-13, 1.212729e-13, 1.215501e-13, 1.21443e-13, 
    1.217223e-13, 1.2111e-13, 1.216312e-13, 1.209766e-13, 1.210341e-13, 
    1.212118e-13, 1.215689e-13, 1.21648e-13, 1.217322e-13, 1.216802e-13, 
    1.214278e-13, 1.213864e-13, 1.212075e-13, 1.21158e-13, 1.210215e-13, 
    1.209085e-13, 1.210118e-13, 1.211202e-13, 1.214279e-13, 1.21705e-13, 
    1.220067e-13, 1.220805e-13, 1.224324e-13, 1.221459e-13, 1.226183e-13, 
    1.222165e-13, 1.229118e-13, 1.216615e-13, 1.222049e-13, 1.212199e-13, 
    1.213262e-13, 1.215183e-13, 1.219585e-13, 1.21721e-13, 1.219988e-13, 
    1.213848e-13, 1.210657e-13, 1.209832e-13, 1.208289e-13, 1.209867e-13, 
    1.209739e-13, 1.211247e-13, 1.210763e-13, 1.214382e-13, 1.212438e-13, 
    1.217956e-13, 1.219966e-13, 1.225637e-13, 1.229107e-13, 1.232636e-13, 
    1.234192e-13, 1.234666e-13, 1.234864e-13 ;

 LITR2C_vr =
  0.001107536, 0.001107535, 0.001107535, 0.001107534, 0.001107534, 
    0.001107534, 0.001107535, 0.001107535, 0.001107535, 0.001107536, 
    0.001107532, 0.001107534, 0.00110753, 0.001107531, 0.001107529, 
    0.00110753, 0.001107528, 0.001107529, 0.001107527, 0.001107528, 
    0.001107526, 0.001107527, 0.001107525, 0.001107526, 0.001107526, 
    0.001107527, 0.001107533, 0.001107532, 0.001107534, 0.001107533, 
    0.001107533, 0.001107534, 0.001107535, 0.001107536, 0.001107536, 
    0.001107535, 0.001107533, 0.001107534, 0.001107533, 0.001107533, 
    0.001107531, 0.001107532, 0.001107529, 0.00110753, 0.001107528, 
    0.001107528, 0.001107528, 0.001107528, 0.001107528, 0.001107529, 
    0.001107528, 0.001107529, 0.001107532, 0.001107531, 0.001107533, 
    0.001107535, 0.001107535, 0.001107536, 0.001107536, 0.001107536, 
    0.001107535, 0.001107534, 0.001107533, 0.001107533, 0.001107533, 
    0.001107531, 0.001107531, 0.001107529, 0.001107529, 0.001107529, 
    0.001107528, 0.001107528, 0.001107528, 0.001107527, 0.001107529, 
    0.001107528, 0.001107529, 0.001107529, 0.001107532, 0.001107534, 
    0.001107534, 0.001107535, 0.001107536, 0.001107535, 0.001107535, 
    0.001107535, 0.001107534, 0.001107534, 0.001107533, 0.001107533, 
    0.00110753, 0.001107532, 0.001107528, 0.001107529, 0.001107528, 
    0.001107529, 0.001107528, 0.001107529, 0.001107527, 0.001107527, 
    0.001107527, 0.001107526, 0.001107529, 0.001107528, 0.001107534, 
    0.001107534, 0.001107534, 0.001107535, 0.001107535, 0.001107536, 
    0.001107535, 0.001107535, 0.001107534, 0.001107534, 0.001107533, 
    0.001107532, 0.001107531, 0.00110753, 0.001107529, 0.001107529, 
    0.001107529, 0.001107529, 0.001107529, 0.001107529, 0.001107527, 
    0.001107528, 0.001107526, 0.001107527, 0.001107527, 0.001107527, 
    0.001107534, 0.001107535, 0.001107535, 0.001107535, 0.001107536, 
    0.001107535, 0.001107535, 0.001107533, 0.001107533, 0.001107533, 
    0.001107532, 0.001107532, 0.00110753, 0.001107529, 0.001107528, 
    0.001107528, 0.001107528, 0.001107528, 0.001107529, 0.001107528, 
    0.001107528, 0.001107528, 0.001107527, 0.001107527, 0.001107527, 
    0.001107527, 0.001107535, 0.001107534, 0.001107534, 0.001107534, 
    0.001107534, 0.001107533, 0.001107533, 0.001107531, 0.001107532, 
    0.001107531, 0.001107532, 0.001107531, 0.001107531, 0.001107531, 
    0.001107529, 0.001107531, 0.001107528, 0.00110753, 0.001107528, 
    0.001107528, 0.001107528, 0.001107528, 0.001107527, 0.001107526, 
    0.001107526, 0.001107525, 0.001107534, 0.001107533, 0.001107533, 
    0.001107533, 0.001107532, 0.001107531, 0.00110753, 0.001107531, 
    0.00110753, 0.00110753, 0.001107531, 0.00110753, 0.001107533, 
    0.001107532, 0.001107533, 0.001107533, 0.00110753, 0.001107532, 
    0.001107529, 0.00110753, 0.001107528, 0.001107529, 0.001107526, 
    0.001107525, 0.001107524, 0.001107523, 0.001107533, 0.001107533, 
    0.001107533, 0.001107532, 0.001107531, 0.00110753, 0.00110753, 
    0.00110753, 0.001107529, 0.001107529, 0.00110753, 0.001107529, 
    0.001107532, 0.00110753, 0.001107533, 0.001107532, 0.001107532, 
    0.001107532, 0.001107531, 0.00110753, 0.001107529, 0.00110753, 
    0.001107526, 0.001107527, 0.001107522, 0.001107524, 0.001107533, 
    0.001107533, 0.001107531, 0.001107532, 0.00110753, 0.001107529, 
    0.001107529, 0.001107528, 0.001107528, 0.001107528, 0.001107529, 
    0.001107528, 0.00110753, 0.001107529, 0.001107531, 0.001107531, 
    0.001107531, 0.001107531, 0.001107531, 0.00110753, 0.00110753, 
    0.001107529, 0.001107528, 0.00110753, 0.001107525, 0.001107528, 
    0.001107532, 0.001107531, 0.001107531, 0.001107532, 0.001107529, 
    0.00110753, 0.001107528, 0.001107529, 0.001107528, 0.001107528, 
    0.001107528, 0.001107529, 0.001107529, 0.00110753, 0.001107531, 
    0.001107532, 0.001107531, 0.001107531, 0.00110753, 0.001107528, 
    0.001107529, 0.001107528, 0.00110753, 0.001107529, 0.001107529, 
    0.001107528, 0.001107531, 0.001107529, 0.001107531, 0.001107531, 
    0.00110753, 0.001107529, 0.001107529, 0.001107528, 0.001107529, 
    0.00110753, 0.00110753, 0.00110753, 0.00110753, 0.001107531, 0.001107531, 
    0.001107531, 0.001107531, 0.00110753, 0.001107529, 0.001107528, 
    0.001107527, 0.001107526, 0.001107527, 0.001107525, 0.001107527, 
    0.001107524, 0.001107529, 0.001107527, 0.00110753, 0.00110753, 
    0.001107529, 0.001107528, 0.001107528, 0.001107528, 0.00110753, 
    0.001107531, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.001107531, 0.001107531, 0.00110753, 0.00110753, 0.001107528, 
    0.001107528, 0.001107526, 0.001107524, 0.001107523, 0.001107523, 
    0.001107522, 0.001107522,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684274e-07, 2.684271e-07, 2.684271e-07, 2.684269e-07, 2.68427e-07, 
    2.684269e-07, 2.684273e-07, 2.684271e-07, 2.684272e-07, 2.684273e-07, 
    2.684265e-07, 2.684269e-07, 2.68426e-07, 2.684263e-07, 2.684257e-07, 
    2.684261e-07, 2.684256e-07, 2.684257e-07, 2.684254e-07, 2.684255e-07, 
    2.684251e-07, 2.684253e-07, 2.684249e-07, 2.684251e-07, 2.684251e-07, 
    2.684253e-07, 2.684268e-07, 2.684265e-07, 2.684268e-07, 2.684268e-07, 
    2.684268e-07, 2.68427e-07, 2.684272e-07, 2.684274e-07, 2.684273e-07, 
    2.684272e-07, 2.684268e-07, 2.684269e-07, 2.684266e-07, 2.684266e-07, 
    2.684262e-07, 2.684264e-07, 2.684258e-07, 2.684259e-07, 2.684255e-07, 
    2.684256e-07, 2.684255e-07, 2.684255e-07, 2.684255e-07, 2.684256e-07, 
    2.684256e-07, 2.684257e-07, 2.684264e-07, 2.684262e-07, 2.684267e-07, 
    2.684271e-07, 2.684273e-07, 2.684274e-07, 2.684274e-07, 2.684274e-07, 
    2.684272e-07, 2.68427e-07, 2.684268e-07, 2.684267e-07, 2.684266e-07, 
    2.684263e-07, 2.684261e-07, 2.684257e-07, 2.684258e-07, 2.684257e-07, 
    2.684256e-07, 2.684254e-07, 2.684254e-07, 2.684253e-07, 2.684257e-07, 
    2.684255e-07, 2.684259e-07, 2.684257e-07, 2.684266e-07, 2.684269e-07, 
    2.68427e-07, 2.684271e-07, 2.684274e-07, 2.684272e-07, 2.684273e-07, 
    2.684271e-07, 2.68427e-07, 2.68427e-07, 2.684267e-07, 2.684268e-07, 
    2.684261e-07, 2.684264e-07, 2.684256e-07, 2.684258e-07, 2.684255e-07, 
    2.684257e-07, 2.684255e-07, 2.684257e-07, 2.684253e-07, 2.684253e-07, 
    2.684253e-07, 2.684251e-07, 2.684257e-07, 2.684255e-07, 2.68427e-07, 
    2.68427e-07, 2.68427e-07, 2.684272e-07, 2.684272e-07, 2.684274e-07, 
    2.684272e-07, 2.684272e-07, 2.68427e-07, 2.684269e-07, 2.684268e-07, 
    2.684266e-07, 2.684263e-07, 2.68426e-07, 2.684258e-07, 2.684256e-07, 
    2.684257e-07, 2.684256e-07, 2.684257e-07, 2.684258e-07, 2.684253e-07, 
    2.684256e-07, 2.684251e-07, 2.684252e-07, 2.684253e-07, 2.684252e-07, 
    2.68427e-07, 2.684271e-07, 2.684273e-07, 2.684271e-07, 2.684274e-07, 
    2.684272e-07, 2.684272e-07, 2.684268e-07, 2.684268e-07, 2.684267e-07, 
    2.684266e-07, 2.684264e-07, 2.684261e-07, 2.684258e-07, 2.684256e-07, 
    2.684256e-07, 2.684256e-07, 2.684255e-07, 2.684257e-07, 2.684255e-07, 
    2.684255e-07, 2.684256e-07, 2.684252e-07, 2.684253e-07, 2.684252e-07, 
    2.684252e-07, 2.684271e-07, 2.68427e-07, 2.68427e-07, 2.684269e-07, 
    2.68427e-07, 2.684267e-07, 2.684266e-07, 2.684262e-07, 2.684264e-07, 
    2.684261e-07, 2.684264e-07, 2.684263e-07, 2.684261e-07, 2.684263e-07, 
    2.684258e-07, 2.684262e-07, 2.684255e-07, 2.684259e-07, 2.684255e-07, 
    2.684256e-07, 2.684255e-07, 2.684254e-07, 2.684253e-07, 2.68425e-07, 
    2.684251e-07, 2.684249e-07, 2.684268e-07, 2.684267e-07, 2.684267e-07, 
    2.684266e-07, 2.684265e-07, 2.684263e-07, 2.68426e-07, 2.684261e-07, 
    2.684259e-07, 2.684259e-07, 2.684262e-07, 2.68426e-07, 2.684266e-07, 
    2.684265e-07, 2.684266e-07, 2.684268e-07, 2.684261e-07, 2.684265e-07, 
    2.684258e-07, 2.68426e-07, 2.684254e-07, 2.684257e-07, 2.684251e-07, 
    2.684249e-07, 2.684246e-07, 2.684243e-07, 2.684266e-07, 2.684267e-07, 
    2.684266e-07, 2.684264e-07, 2.684262e-07, 2.68426e-07, 2.684259e-07, 
    2.684259e-07, 2.684258e-07, 2.684257e-07, 2.684259e-07, 2.684257e-07, 
    2.684265e-07, 2.68426e-07, 2.684268e-07, 2.684266e-07, 2.684264e-07, 
    2.684265e-07, 2.684261e-07, 2.68426e-07, 2.684257e-07, 2.684259e-07, 
    2.684249e-07, 2.684253e-07, 2.684241e-07, 2.684245e-07, 2.684268e-07, 
    2.684266e-07, 2.684263e-07, 2.684264e-07, 2.684259e-07, 2.684258e-07, 
    2.684257e-07, 2.684256e-07, 2.684256e-07, 2.684255e-07, 2.684256e-07, 
    2.684255e-07, 2.68426e-07, 2.684258e-07, 2.684263e-07, 2.684262e-07, 
    2.684262e-07, 2.684263e-07, 2.684261e-07, 2.684259e-07, 2.684259e-07, 
    2.684258e-07, 2.684256e-07, 2.684259e-07, 2.684249e-07, 2.684255e-07, 
    2.684265e-07, 2.684263e-07, 2.684263e-07, 2.684264e-07, 2.684258e-07, 
    2.68426e-07, 2.684255e-07, 2.684257e-07, 2.684254e-07, 2.684255e-07, 
    2.684255e-07, 2.684257e-07, 2.684258e-07, 2.68426e-07, 2.684262e-07, 
    2.684264e-07, 2.684263e-07, 2.684262e-07, 2.684259e-07, 2.684256e-07, 
    2.684257e-07, 2.684254e-07, 2.68426e-07, 2.684258e-07, 2.684259e-07, 
    2.684256e-07, 2.684261e-07, 2.684257e-07, 2.684262e-07, 2.684262e-07, 
    2.68426e-07, 2.684257e-07, 2.684257e-07, 2.684256e-07, 2.684257e-07, 
    2.684259e-07, 2.684259e-07, 2.68426e-07, 2.684261e-07, 2.684262e-07, 
    2.684263e-07, 2.684262e-07, 2.684261e-07, 2.684259e-07, 2.684256e-07, 
    2.684254e-07, 2.684253e-07, 2.68425e-07, 2.684253e-07, 2.684249e-07, 
    2.684252e-07, 2.684246e-07, 2.684257e-07, 2.684252e-07, 2.68426e-07, 
    2.684259e-07, 2.684258e-07, 2.684254e-07, 2.684256e-07, 2.684254e-07, 
    2.684259e-07, 2.684262e-07, 2.684262e-07, 2.684264e-07, 2.684262e-07, 
    2.684262e-07, 2.684261e-07, 2.684262e-07, 2.684259e-07, 2.68426e-07, 
    2.684255e-07, 2.684254e-07, 2.684249e-07, 2.684246e-07, 2.684243e-07, 
    2.684242e-07, 2.684241e-07, 2.684241e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  -2.058761e-25, -1.617598e-25, 7.352717e-27, 7.842898e-26, -4.65672e-26, 
    -2.205815e-26, -2.450906e-27, -4.65672e-26, 7.842898e-26, 3.186177e-26, 
    -7.352717e-27, 6.617445e-26, -7.352717e-27, -2.450906e-27, -9.068351e-26, 
    -1.225453e-25, 3.676358e-26, 1.862688e-25, 6.617445e-26, 1.715634e-26, 
    -9.313441e-26, -2.695996e-26, 1.519561e-25, -1.862688e-25, 8.333079e-26, 
    -3.89694e-25, -7.842898e-26, 1.862688e-25, 9.803622e-26, 9.313441e-26, 
    1.249962e-25, 2.303851e-25, 4.65672e-26, 1.642107e-25, -3.921449e-26, 
    -2.303851e-25, -1.29898e-25, -9.313441e-26, 2.941087e-26, 1.715634e-25, 
    8.333079e-26, 2.499924e-25, 1.617598e-25, -2.303851e-25, 1.911706e-25, 
    7.352717e-27, -2.132288e-25, -1.446034e-25, -1.960724e-26, -1.960724e-26, 
    6.372354e-26, -1.740143e-25, 1.274471e-25, -2.965596e-25, 1.593089e-25, 
    -1.078398e-25, 2.695996e-26, -1.02938e-25, 7.842898e-26, 9.068351e-26, 
    -7.352717e-27, -1.421525e-25, 1.789161e-25, 1.715634e-26, 8.333079e-26, 
    2.450905e-26, 1.446034e-25, 1.274471e-25, -1.715634e-26, -1.078398e-25, 
    2.695996e-26, 1.862688e-25, 1.02938e-25, -1.397016e-25, 7.352717e-26, 
    9.803622e-27, 1.519561e-25, 7.352717e-26, -3.235195e-25, 4.41163e-26, 
    -1.519561e-25, 2.303851e-25, 1.960724e-26, -1.470543e-25, -7.352717e-26, 
    1.078398e-25, 1.02938e-25, -1.127417e-25, 4.166539e-26, -9.558531e-26, 
    -1.421525e-25, -1.053889e-25, -2.450905e-26, 1.54407e-25, -9.803622e-27, 
    -5.146902e-26, 6.372354e-26, -3.235195e-25, 1.102908e-25, 3.921449e-26, 
    -2.254833e-25, -8.333079e-26, 2.058761e-25, 1.02938e-25, -1.666616e-25, 
    -4.901811e-26, -1.078398e-25, -1.495052e-25, -4.65672e-26, -1.004871e-25, 
    -3.921449e-26, 1.887197e-25, 5.882173e-26, -4.41163e-26, -1.715634e-26, 
    6.617445e-26, -1.225453e-25, -4.166539e-26, -5.146902e-26, -7.352717e-27, 
    -4.166539e-26, -4.65672e-26, -5.637083e-26, 1.715634e-25, 8.087988e-26, 
    4.901811e-27, -2.279342e-25, -7.352717e-27, 2.426396e-25, -1.519561e-25, 
    1.176435e-25, 1.446034e-25, 6.372354e-26, 7.842898e-26, 2.401887e-25, 
    -9.558531e-26, 7.107626e-26, 1.519561e-25, -4.901811e-27, 8.333079e-26, 
    -7.352717e-27, -8.333079e-26, -1.960724e-26, -2.524433e-25, 1.421525e-25, 
    -1.495052e-25, -1.691125e-25, 7.107626e-26, -3.431268e-26, -7.352717e-26, 
    -1.887197e-25, 9.068351e-26, -6.862535e-26, 8.578169e-26, -4.166539e-26, 
    9.803622e-27, -1.519561e-25, 7.597807e-26, -2.181306e-25, -9.558531e-26, 
    6.127264e-26, 7.842898e-26, -1.519561e-25, 1.102908e-25, 3.676358e-26, 
    -9.558531e-26, 1.691125e-25, 2.205815e-26, 3.186177e-26, -4.901811e-27, 
    -7.597807e-26, -1.127417e-25, 1.274471e-25, 1.225453e-26, -9.558531e-26, 
    -2.450905e-26, -6.862535e-26, 1.02938e-25, -1.789161e-25, 8.82326e-26, 
    -6.862535e-26, 3.014614e-25, -1.078398e-25, 4.901811e-26, 9.558531e-26, 
    4.41163e-26, 8.333079e-26, -3.504795e-25, -4.41163e-26, -2.009742e-25, 
    -1.347998e-25, -3.38225e-25, 6.862535e-26, 1.200944e-25, -1.274471e-25, 
    -4.41163e-26, -9.803622e-27, 1.446034e-25, 1.911706e-25, -8.82326e-26, 
    -9.803622e-26, -5.882173e-26, -1.838179e-25, 6.862535e-26, -1.225453e-25, 
    -1.02938e-25, -1.764652e-25, -4.41163e-26, 1.372507e-25, 3.921449e-26, 
    1.127417e-25, -3.676358e-26, 6.127264e-26, -1.519561e-25, -2.205815e-26, 
    5.146902e-26, 7.107626e-26, 7.597807e-26, 3.921449e-26, 1.495052e-25, 
    -2.941087e-26, -1.519561e-25, 2.034252e-25, -2.205815e-26, -7.597807e-26, 
    -8.578169e-26, -1.862688e-25, -9.558531e-26, -8.333079e-26, 
    -8.087988e-26, -2.279342e-25, -2.499924e-25, -2.181306e-25, 
    -1.960724e-26, -1.715634e-26, -1.911706e-25, 8.578169e-26, -1.838179e-25, 
    -5.391992e-26, -5.146902e-26, -6.127264e-26, 1.470543e-26, 4.41163e-26, 
    -2.450906e-27, -1.56858e-25, -1.127417e-25, 7.107626e-26, -1.249962e-25, 
    -8.333079e-26, 2.450906e-25, -1.960724e-25, -3.186177e-26, -3.431268e-26, 
    2.352869e-25, -3.431268e-26, 5.391992e-26, -9.313441e-26, 7.842898e-26, 
    -1.715634e-26, -2.450906e-27, 3.186177e-25, -1.862688e-25, -5.882173e-26, 
    -1.715634e-25, -9.803622e-27, 1.274471e-25, 4.901811e-27, -2.205815e-26, 
    2.867559e-25, 1.960724e-26, 1.372507e-25, -1.078398e-25, -1.666616e-25, 
    -1.347998e-25, -2.941087e-26, -7.842898e-26, -1.151926e-25, 4.65672e-26, 
    -7.597807e-26, 3.921449e-26, -9.803622e-27, -1.053889e-25, -1.887197e-25, 
    -1.519561e-25, 3.259704e-25, -8.087988e-26, 1.078398e-25, -1.02938e-25, 
    -1.715634e-26, 1.053889e-25, -9.068351e-26, -5.882173e-26, 2.990105e-25, 
    -9.803622e-26, 3.333231e-25, -1.470543e-25, -1.519561e-25, 3.431268e-26, 
    -2.524433e-25, 3.921449e-26, 7.352717e-27, 8.087988e-26, -2.450905e-26, 
    1.078398e-25, 1.715634e-26, -2.450906e-27, 6.617445e-26, -1.642107e-25, 
    -2.08327e-25, 8.578169e-26, -2.205815e-26, -2.181306e-25, -1.530638e-41, 
    -7.597807e-26, 7.352717e-27, -1.789161e-25, -1.372507e-25, 4.117521e-25, 
    -8.578169e-26, -5.146902e-26, 5.882173e-26, -3.186177e-26, -6.127264e-26, 
    -1.691125e-25, -1.053889e-25, 1.397016e-25, 5.146902e-26, 9.558531e-26, 
    2.548942e-25, -1.078398e-25, -1.151926e-25, -1.470543e-26, -8.333079e-26, 
    -5.882173e-26, 3.921449e-26, -5.146902e-26, -1.200944e-25, 2.450905e-26,
  2.67626e-32, 2.676257e-32, 2.676258e-32, 2.676255e-32, 2.676257e-32, 
    2.676255e-32, 2.676259e-32, 2.676257e-32, 2.676258e-32, 2.676259e-32, 
    2.676251e-32, 2.676255e-32, 2.676247e-32, 2.676249e-32, 2.676243e-32, 
    2.676247e-32, 2.676242e-32, 2.676243e-32, 2.67624e-32, 2.676241e-32, 
    2.676237e-32, 2.676239e-32, 2.676235e-32, 2.676237e-32, 2.676237e-32, 
    2.676239e-32, 2.676254e-32, 2.676252e-32, 2.676255e-32, 2.676254e-32, 
    2.676254e-32, 2.676257e-32, 2.676258e-32, 2.67626e-32, 2.676259e-32, 
    2.676258e-32, 2.676254e-32, 2.676255e-32, 2.676252e-32, 2.676252e-32, 
    2.676248e-32, 2.67625e-32, 2.676244e-32, 2.676246e-32, 2.676241e-32, 
    2.676242e-32, 2.676241e-32, 2.676241e-32, 2.676241e-32, 2.676242e-32, 
    2.676242e-32, 2.676243e-32, 2.67625e-32, 2.676248e-32, 2.676254e-32, 
    2.676257e-32, 2.676259e-32, 2.676261e-32, 2.676261e-32, 2.67626e-32, 
    2.676258e-32, 2.676256e-32, 2.676254e-32, 2.676253e-32, 2.676252e-32, 
    2.676249e-32, 2.676247e-32, 2.676244e-32, 2.676244e-32, 2.676243e-32, 
    2.676242e-32, 2.67624e-32, 2.67624e-32, 2.67624e-32, 2.676243e-32, 
    2.676241e-32, 2.676244e-32, 2.676244e-32, 2.676252e-32, 2.676255e-32, 
    2.676256e-32, 2.676257e-32, 2.67626e-32, 2.676258e-32, 2.676259e-32, 
    2.676257e-32, 2.676256e-32, 2.676257e-32, 2.676253e-32, 2.676254e-32, 
    2.676247e-32, 2.67625e-32, 2.676242e-32, 2.676244e-32, 2.676242e-32, 
    2.676243e-32, 2.676241e-32, 2.676243e-32, 2.676239e-32, 2.676239e-32, 
    2.676239e-32, 2.676237e-32, 2.676243e-32, 2.676241e-32, 2.676257e-32, 
    2.676257e-32, 2.676256e-32, 2.676258e-32, 2.676258e-32, 2.67626e-32, 
    2.676259e-32, 2.676258e-32, 2.676256e-32, 2.676255e-32, 2.676254e-32, 
    2.676252e-32, 2.67625e-32, 2.676246e-32, 2.676244e-32, 2.676242e-32, 
    2.676243e-32, 2.676242e-32, 2.676244e-32, 2.676244e-32, 2.676239e-32, 
    2.676242e-32, 2.676237e-32, 2.676238e-32, 2.67624e-32, 2.676238e-32, 
    2.676257e-32, 2.676257e-32, 2.676259e-32, 2.676257e-32, 2.67626e-32, 
    2.676259e-32, 2.676258e-32, 2.676254e-32, 2.676254e-32, 2.676253e-32, 
    2.676252e-32, 2.67625e-32, 2.676247e-32, 2.676244e-32, 2.676242e-32, 
    2.676242e-32, 2.676242e-32, 2.676242e-32, 2.676243e-32, 2.676241e-32, 
    2.676241e-32, 2.676242e-32, 2.676238e-32, 2.676239e-32, 2.676238e-32, 
    2.676239e-32, 2.676257e-32, 2.676256e-32, 2.676257e-32, 2.676256e-32, 
    2.676256e-32, 2.676253e-32, 2.676252e-32, 2.676248e-32, 2.67625e-32, 
    2.676247e-32, 2.67625e-32, 2.676249e-32, 2.676247e-32, 2.67625e-32, 
    2.676244e-32, 2.676248e-32, 2.676242e-32, 2.676245e-32, 2.676241e-32, 
    2.676242e-32, 2.676241e-32, 2.67624e-32, 2.676239e-32, 2.676236e-32, 
    2.676237e-32, 2.676235e-32, 2.676255e-32, 2.676254e-32, 2.676254e-32, 
    2.676252e-32, 2.676252e-32, 2.676249e-32, 2.676246e-32, 2.676247e-32, 
    2.676245e-32, 2.676245e-32, 2.676248e-32, 2.676246e-32, 2.676253e-32, 
    2.676252e-32, 2.676252e-32, 2.676254e-32, 2.676247e-32, 2.676251e-32, 
    2.676244e-32, 2.676246e-32, 2.67624e-32, 2.676243e-32, 2.676237e-32, 
    2.676234e-32, 2.676232e-32, 2.676229e-32, 2.676253e-32, 2.676254e-32, 
    2.676252e-32, 2.67625e-32, 2.676248e-32, 2.676246e-32, 2.676246e-32, 
    2.676245e-32, 2.676244e-32, 2.676243e-32, 2.676245e-32, 2.676243e-32, 
    2.676251e-32, 2.676247e-32, 2.676254e-32, 2.676252e-32, 2.67625e-32, 
    2.676251e-32, 2.676248e-32, 2.676247e-32, 2.676244e-32, 2.676245e-32, 
    2.676235e-32, 2.67624e-32, 2.676227e-32, 2.676231e-32, 2.676254e-32, 
    2.676253e-32, 2.676249e-32, 2.676251e-32, 2.676246e-32, 2.676244e-32, 
    2.676243e-32, 2.676242e-32, 2.676242e-32, 2.676241e-32, 2.676242e-32, 
    2.676241e-32, 2.676246e-32, 2.676244e-32, 2.676249e-32, 2.676248e-32, 
    2.676249e-32, 2.676249e-32, 2.676247e-32, 2.676245e-32, 2.676245e-32, 
    2.676244e-32, 2.676242e-32, 2.676246e-32, 2.676235e-32, 2.676242e-32, 
    2.676252e-32, 2.676249e-32, 2.676249e-32, 2.67625e-32, 2.676244e-32, 
    2.676247e-32, 2.676241e-32, 2.676243e-32, 2.67624e-32, 2.676242e-32, 
    2.676242e-32, 2.676243e-32, 2.676244e-32, 2.676247e-32, 2.676248e-32, 
    2.67625e-32, 2.676249e-32, 2.676248e-32, 2.676245e-32, 2.676242e-32, 
    2.676243e-32, 2.67624e-32, 2.676246e-32, 2.676244e-32, 2.676245e-32, 
    2.676242e-32, 2.676247e-32, 2.676243e-32, 2.676249e-32, 2.676248e-32, 
    2.676247e-32, 2.676244e-32, 2.676243e-32, 2.676242e-32, 2.676243e-32, 
    2.676245e-32, 2.676245e-32, 2.676247e-32, 2.676247e-32, 2.676248e-32, 
    2.676249e-32, 2.676248e-32, 2.676247e-32, 2.676245e-32, 2.676242e-32, 
    2.67624e-32, 2.676239e-32, 2.676236e-32, 2.676239e-32, 2.676235e-32, 
    2.676238e-32, 2.676232e-32, 2.676243e-32, 2.676238e-32, 2.676247e-32, 
    2.676246e-32, 2.676244e-32, 2.67624e-32, 2.676242e-32, 2.67624e-32, 
    2.676245e-32, 2.676248e-32, 2.676249e-32, 2.67625e-32, 2.676249e-32, 
    2.676249e-32, 2.676247e-32, 2.676248e-32, 2.676245e-32, 2.676246e-32, 
    2.676242e-32, 2.67624e-32, 2.676235e-32, 2.676232e-32, 2.676229e-32, 
    2.676228e-32, 2.676227e-32, 2.676227e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.311877e-15, 3.320829e-15, 3.31909e-15, 3.326303e-15, 3.322303e-15, 
    3.327025e-15, 3.313693e-15, 3.321183e-15, 3.316403e-15, 3.312684e-15, 
    3.340281e-15, 3.326625e-15, 3.354452e-15, 3.345759e-15, 3.367581e-15, 
    3.353098e-15, 3.370498e-15, 3.367166e-15, 3.377198e-15, 3.374326e-15, 
    3.387137e-15, 3.378523e-15, 3.393773e-15, 3.385082e-15, 3.386441e-15, 
    3.378238e-15, 3.329378e-15, 3.338581e-15, 3.328831e-15, 3.330145e-15, 
    3.329556e-15, 3.322385e-15, 3.318767e-15, 3.311194e-15, 3.31257e-15, 
    3.318133e-15, 3.330735e-15, 3.326461e-15, 3.337233e-15, 3.33699e-15, 
    3.348965e-15, 3.343568e-15, 3.363669e-15, 3.357962e-15, 3.374445e-15, 
    3.370303e-15, 3.37425e-15, 3.373054e-15, 3.374266e-15, 3.36819e-15, 
    3.370794e-15, 3.365445e-15, 3.344578e-15, 3.350716e-15, 3.332396e-15, 
    3.321356e-15, 3.314022e-15, 3.308811e-15, 3.309548e-15, 3.310952e-15, 
    3.318166e-15, 3.324945e-15, 3.330106e-15, 3.333557e-15, 3.336955e-15, 
    3.347228e-15, 3.352665e-15, 3.364822e-15, 3.362631e-15, 3.366343e-15, 
    3.369891e-15, 3.37584e-15, 3.374862e-15, 3.377481e-15, 3.366247e-15, 
    3.373714e-15, 3.361383e-15, 3.364757e-15, 3.33787e-15, 3.327615e-15, 
    3.323244e-15, 3.319424e-15, 3.310114e-15, 3.316544e-15, 3.31401e-15, 
    3.320039e-15, 3.323867e-15, 3.321974e-15, 3.333651e-15, 3.329113e-15, 
    3.352987e-15, 3.342712e-15, 3.369477e-15, 3.363081e-15, 3.37101e-15, 
    3.366965e-15, 3.373893e-15, 3.367659e-15, 3.378457e-15, 3.380805e-15, 
    3.3792e-15, 3.385366e-15, 3.367313e-15, 3.37425e-15, 3.321921e-15, 
    3.322229e-15, 3.323668e-15, 3.317342e-15, 3.316955e-15, 3.311156e-15, 
    3.316317e-15, 3.318513e-15, 3.324089e-15, 3.327384e-15, 3.330516e-15, 
    3.337397e-15, 3.345074e-15, 3.355798e-15, 3.363496e-15, 3.368651e-15, 
    3.365491e-15, 3.368281e-15, 3.365162e-15, 3.3637e-15, 3.379924e-15, 
    3.370817e-15, 3.384479e-15, 3.383724e-15, 3.377543e-15, 3.383809e-15, 
    3.322446e-15, 3.32067e-15, 3.314496e-15, 3.319328e-15, 3.310524e-15, 
    3.315452e-15, 3.318284e-15, 3.329206e-15, 3.331606e-15, 3.333828e-15, 
    3.338216e-15, 3.343844e-15, 3.353706e-15, 3.362279e-15, 3.370098e-15, 
    3.369525e-15, 3.369727e-15, 3.371471e-15, 3.367148e-15, 3.372181e-15, 
    3.373025e-15, 3.370817e-15, 3.383623e-15, 3.379967e-15, 3.383708e-15, 
    3.381328e-15, 3.321248e-15, 3.324237e-15, 3.322622e-15, 3.325658e-15, 
    3.323518e-15, 3.333027e-15, 3.335875e-15, 3.349194e-15, 3.343733e-15, 
    3.352425e-15, 3.344617e-15, 3.346001e-15, 3.352705e-15, 3.34504e-15, 
    3.361805e-15, 3.350439e-15, 3.371539e-15, 3.3602e-15, 3.372249e-15, 
    3.370064e-15, 3.373682e-15, 3.376921e-15, 3.380994e-15, 3.388503e-15, 
    3.386765e-15, 3.393042e-15, 3.328692e-15, 3.332564e-15, 3.332225e-15, 
    3.336277e-15, 3.339272e-15, 3.345762e-15, 3.356158e-15, 3.352251e-15, 
    3.359425e-15, 3.360863e-15, 3.349965e-15, 3.356657e-15, 3.335156e-15, 
    3.338632e-15, 3.336564e-15, 3.328996e-15, 3.353149e-15, 3.340762e-15, 
    3.363623e-15, 3.356923e-15, 3.376459e-15, 3.366748e-15, 3.385808e-15, 
    3.393937e-15, 3.401588e-15, 3.410509e-15, 3.334679e-15, 3.332048e-15, 
    3.336759e-15, 3.34327e-15, 3.349311e-15, 3.357332e-15, 3.358153e-15, 
    3.359654e-15, 3.363543e-15, 3.366811e-15, 3.360127e-15, 3.36763e-15, 
    3.339435e-15, 3.354224e-15, 3.331052e-15, 3.338034e-15, 3.342887e-15, 
    3.34076e-15, 3.351805e-15, 3.354405e-15, 3.364962e-15, 3.359507e-15, 
    3.39193e-15, 3.377602e-15, 3.4173e-15, 3.406227e-15, 3.331129e-15, 
    3.334671e-15, 3.346984e-15, 3.341128e-15, 3.357868e-15, 3.361983e-15, 
    3.365327e-15, 3.369598e-15, 3.37006e-15, 3.372589e-15, 3.368444e-15, 
    3.372426e-15, 3.357349e-15, 3.36409e-15, 3.345579e-15, 3.350088e-15, 
    3.348015e-15, 3.345739e-15, 3.352761e-15, 3.360232e-15, 3.360394e-15, 
    3.362788e-15, 3.369525e-15, 3.357936e-15, 3.393772e-15, 3.371656e-15, 
    3.338531e-15, 3.345343e-15, 3.346318e-15, 3.34368e-15, 3.36157e-15, 
    3.355092e-15, 3.372528e-15, 3.36782e-15, 3.375533e-15, 3.371701e-15, 
    3.371137e-15, 3.366213e-15, 3.363145e-15, 3.355389e-15, 3.349073e-15, 
    3.344063e-15, 3.345229e-15, 3.350731e-15, 3.36069e-15, 3.370101e-15, 
    3.36804e-15, 3.374947e-15, 3.356655e-15, 3.364329e-15, 3.361363e-15, 
    3.369095e-15, 3.352147e-15, 3.366573e-15, 3.348454e-15, 3.350045e-15, 
    3.354964e-15, 3.364848e-15, 3.367037e-15, 3.369369e-15, 3.36793e-15, 
    3.360943e-15, 3.359799e-15, 3.354845e-15, 3.353475e-15, 3.349699e-15, 
    3.346569e-15, 3.349428e-15, 3.352428e-15, 3.360947e-15, 3.368614e-15, 
    3.376966e-15, 3.37901e-15, 3.388747e-15, 3.380818e-15, 3.393895e-15, 
    3.382773e-15, 3.402018e-15, 3.367413e-15, 3.382451e-15, 3.355188e-15, 
    3.358131e-15, 3.363447e-15, 3.375632e-15, 3.369059e-15, 3.376747e-15, 
    3.359754e-15, 3.35092e-15, 3.348636e-15, 3.344367e-15, 3.348733e-15, 
    3.348378e-15, 3.352554e-15, 3.351213e-15, 3.361229e-15, 3.355851e-15, 
    3.371122e-15, 3.376687e-15, 3.392383e-15, 3.401987e-15, 3.411756e-15, 
    3.416062e-15, 3.417373e-15, 3.417921e-15 ;

 LITR2N_vr =
  1.532748e-05, 1.532746e-05, 1.532747e-05, 1.532745e-05, 1.532746e-05, 
    1.532745e-05, 1.532748e-05, 1.532746e-05, 1.532747e-05, 1.532748e-05, 
    1.532743e-05, 1.532745e-05, 1.53274e-05, 1.532742e-05, 1.532738e-05, 
    1.532741e-05, 1.532738e-05, 1.532738e-05, 1.532736e-05, 1.532737e-05, 
    1.532735e-05, 1.532736e-05, 1.532734e-05, 1.532735e-05, 1.532735e-05, 
    1.532736e-05, 1.532745e-05, 1.532743e-05, 1.532745e-05, 1.532745e-05, 
    1.532745e-05, 1.532746e-05, 1.532747e-05, 1.532748e-05, 1.532748e-05, 
    1.532747e-05, 1.532745e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532741e-05, 1.532742e-05, 1.532739e-05, 1.53274e-05, 1.532737e-05, 
    1.532738e-05, 1.532737e-05, 1.532737e-05, 1.532737e-05, 1.532738e-05, 
    1.532738e-05, 1.532738e-05, 1.532742e-05, 1.532741e-05, 1.532744e-05, 
    1.532746e-05, 1.532748e-05, 1.532749e-05, 1.532748e-05, 1.532748e-05, 
    1.532747e-05, 1.532746e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532737e-05, 1.532737e-05, 1.532736e-05, 1.532738e-05, 
    1.532737e-05, 1.532739e-05, 1.532739e-05, 1.532743e-05, 1.532745e-05, 
    1.532746e-05, 1.532747e-05, 1.532748e-05, 1.532747e-05, 1.532748e-05, 
    1.532747e-05, 1.532746e-05, 1.532746e-05, 1.532744e-05, 1.532745e-05, 
    1.532741e-05, 1.532742e-05, 1.532738e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532737e-05, 1.532738e-05, 1.532736e-05, 1.532736e-05, 
    1.532736e-05, 1.532735e-05, 1.532738e-05, 1.532737e-05, 1.532746e-05, 
    1.532746e-05, 1.532746e-05, 1.532747e-05, 1.532747e-05, 1.532748e-05, 
    1.532747e-05, 1.532747e-05, 1.532746e-05, 1.532745e-05, 1.532745e-05, 
    1.532743e-05, 1.532742e-05, 1.53274e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532738e-05, 1.532739e-05, 1.532739e-05, 1.532736e-05, 
    1.532738e-05, 1.532735e-05, 1.532735e-05, 1.532736e-05, 1.532735e-05, 
    1.532746e-05, 1.532746e-05, 1.532747e-05, 1.532747e-05, 1.532748e-05, 
    1.532747e-05, 1.532747e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532743e-05, 1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532738e-05, 1.532738e-05, 1.532738e-05, 1.532737e-05, 
    1.532737e-05, 1.532738e-05, 1.532735e-05, 1.532736e-05, 1.532735e-05, 
    1.532736e-05, 1.532746e-05, 1.532746e-05, 1.532746e-05, 1.532746e-05, 
    1.532746e-05, 1.532744e-05, 1.532744e-05, 1.532741e-05, 1.532742e-05, 
    1.532741e-05, 1.532742e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 
    1.532739e-05, 1.532741e-05, 1.532738e-05, 1.53274e-05, 1.532737e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532736e-05, 1.532734e-05, 
    1.532735e-05, 1.532734e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532744e-05, 1.532743e-05, 1.532742e-05, 1.53274e-05, 1.532741e-05, 
    1.53274e-05, 1.532739e-05, 1.532741e-05, 1.53274e-05, 1.532744e-05, 
    1.532743e-05, 1.532744e-05, 1.532745e-05, 1.532741e-05, 1.532743e-05, 
    1.532739e-05, 1.53274e-05, 1.532737e-05, 1.532738e-05, 1.532735e-05, 
    1.532734e-05, 1.532732e-05, 1.532731e-05, 1.532744e-05, 1.532744e-05, 
    1.532744e-05, 1.532742e-05, 1.532741e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532739e-05, 1.532738e-05, 1.53274e-05, 1.532738e-05, 
    1.532743e-05, 1.53274e-05, 1.532744e-05, 1.532743e-05, 1.532742e-05, 
    1.532743e-05, 1.532741e-05, 1.53274e-05, 1.532739e-05, 1.53274e-05, 
    1.532734e-05, 1.532736e-05, 1.53273e-05, 1.532731e-05, 1.532744e-05, 
    1.532744e-05, 1.532742e-05, 1.532743e-05, 1.53274e-05, 1.532739e-05, 
    1.532739e-05, 1.532738e-05, 1.532738e-05, 1.532737e-05, 1.532738e-05, 
    1.532737e-05, 1.53274e-05, 1.532739e-05, 1.532742e-05, 1.532741e-05, 
    1.532742e-05, 1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532739e-05, 
    1.532739e-05, 1.532738e-05, 1.53274e-05, 1.532734e-05, 1.532738e-05, 
    1.532743e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 1.532739e-05, 
    1.53274e-05, 1.532737e-05, 1.532738e-05, 1.532737e-05, 1.532737e-05, 
    1.532738e-05, 1.532738e-05, 1.532739e-05, 1.53274e-05, 1.532741e-05, 
    1.532742e-05, 1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532737e-05, 1.53274e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532741e-05, 1.532738e-05, 1.532742e-05, 1.532741e-05, 
    1.53274e-05, 1.532739e-05, 1.532738e-05, 1.532738e-05, 1.532738e-05, 
    1.532739e-05, 1.53274e-05, 1.53274e-05, 1.532741e-05, 1.532741e-05, 
    1.532742e-05, 1.532741e-05, 1.532741e-05, 1.532739e-05, 1.532738e-05, 
    1.532736e-05, 1.532736e-05, 1.532734e-05, 1.532736e-05, 1.532734e-05, 
    1.532736e-05, 1.532732e-05, 1.532738e-05, 1.532736e-05, 1.53274e-05, 
    1.53274e-05, 1.532739e-05, 1.532737e-05, 1.532738e-05, 1.532737e-05, 
    1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 
    1.532742e-05, 1.532741e-05, 1.532741e-05, 1.532739e-05, 1.53274e-05, 
    1.532738e-05, 1.532737e-05, 1.532734e-05, 1.532732e-05, 1.53273e-05, 
    1.53273e-05, 1.53273e-05, 1.532729e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.196551e-13, 1.199785e-13, 1.199157e-13, 1.201763e-13, 1.200318e-13, 
    1.202024e-13, 1.197207e-13, 1.199913e-13, 1.198186e-13, 1.196843e-13, 
    1.206813e-13, 1.201879e-13, 1.211933e-13, 1.208792e-13, 1.216676e-13, 
    1.211444e-13, 1.21773e-13, 1.216526e-13, 1.220151e-13, 1.219113e-13, 
    1.223742e-13, 1.22063e-13, 1.226139e-13, 1.222999e-13, 1.22349e-13, 
    1.220527e-13, 1.202874e-13, 1.206199e-13, 1.202676e-13, 1.203151e-13, 
    1.202938e-13, 1.200347e-13, 1.19904e-13, 1.196304e-13, 1.196801e-13, 
    1.198811e-13, 1.203364e-13, 1.20182e-13, 1.205712e-13, 1.205624e-13, 
    1.20995e-13, 1.208e-13, 1.215263e-13, 1.213201e-13, 1.219156e-13, 
    1.21766e-13, 1.219086e-13, 1.218654e-13, 1.219092e-13, 1.216896e-13, 
    1.217837e-13, 1.215905e-13, 1.208366e-13, 1.210583e-13, 1.203964e-13, 
    1.199976e-13, 1.197326e-13, 1.195443e-13, 1.19571e-13, 1.196217e-13, 
    1.198823e-13, 1.201272e-13, 1.203137e-13, 1.204384e-13, 1.205611e-13, 
    1.209323e-13, 1.211287e-13, 1.215679e-13, 1.214888e-13, 1.216229e-13, 
    1.217511e-13, 1.21966e-13, 1.219307e-13, 1.220253e-13, 1.216194e-13, 
    1.218892e-13, 1.214437e-13, 1.215656e-13, 1.205942e-13, 1.202237e-13, 
    1.200658e-13, 1.199277e-13, 1.195914e-13, 1.198237e-13, 1.197321e-13, 
    1.1995e-13, 1.200883e-13, 1.200199e-13, 1.204418e-13, 1.202778e-13, 
    1.211403e-13, 1.207691e-13, 1.217361e-13, 1.21505e-13, 1.217915e-13, 
    1.216454e-13, 1.218957e-13, 1.216704e-13, 1.220606e-13, 1.221454e-13, 
    1.220874e-13, 1.223102e-13, 1.216579e-13, 1.219086e-13, 1.20018e-13, 
    1.200291e-13, 1.200811e-13, 1.198525e-13, 1.198386e-13, 1.19629e-13, 
    1.198155e-13, 1.198948e-13, 1.200963e-13, 1.202153e-13, 1.203285e-13, 
    1.205771e-13, 1.208544e-13, 1.212419e-13, 1.2152e-13, 1.217063e-13, 
    1.215921e-13, 1.216929e-13, 1.215802e-13, 1.215274e-13, 1.221136e-13, 
    1.217846e-13, 1.222782e-13, 1.222509e-13, 1.220276e-13, 1.222539e-13, 
    1.20037e-13, 1.199728e-13, 1.197497e-13, 1.199243e-13, 1.196062e-13, 
    1.197843e-13, 1.198866e-13, 1.202812e-13, 1.203679e-13, 1.204482e-13, 
    1.206067e-13, 1.2081e-13, 1.211663e-13, 1.214761e-13, 1.217585e-13, 
    1.217379e-13, 1.217451e-13, 1.218082e-13, 1.21652e-13, 1.218338e-13, 
    1.218643e-13, 1.217846e-13, 1.222472e-13, 1.221151e-13, 1.222503e-13, 
    1.221643e-13, 1.199936e-13, 1.201016e-13, 1.200433e-13, 1.20153e-13, 
    1.200757e-13, 1.204192e-13, 1.205221e-13, 1.210033e-13, 1.20806e-13, 
    1.211201e-13, 1.20838e-13, 1.208879e-13, 1.211302e-13, 1.208532e-13, 
    1.214589e-13, 1.210483e-13, 1.218106e-13, 1.214009e-13, 1.218363e-13, 
    1.217573e-13, 1.218881e-13, 1.220051e-13, 1.221522e-13, 1.224235e-13, 
    1.223607e-13, 1.225875e-13, 1.202626e-13, 1.204025e-13, 1.203902e-13, 
    1.205367e-13, 1.206449e-13, 1.208793e-13, 1.212549e-13, 1.211138e-13, 
    1.213729e-13, 1.214249e-13, 1.210312e-13, 1.212729e-13, 1.204962e-13, 
    1.206217e-13, 1.20547e-13, 1.202736e-13, 1.211462e-13, 1.206987e-13, 
    1.215246e-13, 1.212826e-13, 1.219884e-13, 1.216375e-13, 1.223262e-13, 
    1.226199e-13, 1.228963e-13, 1.232186e-13, 1.204789e-13, 1.203839e-13, 
    1.205541e-13, 1.207893e-13, 1.210075e-13, 1.212973e-13, 1.21327e-13, 
    1.213812e-13, 1.215218e-13, 1.216398e-13, 1.213983e-13, 1.216694e-13, 
    1.206507e-13, 1.211851e-13, 1.203479e-13, 1.206001e-13, 1.207755e-13, 
    1.206986e-13, 1.210976e-13, 1.211916e-13, 1.21573e-13, 1.213759e-13, 
    1.225473e-13, 1.220297e-13, 1.234639e-13, 1.230639e-13, 1.203506e-13, 
    1.204786e-13, 1.209235e-13, 1.207119e-13, 1.213167e-13, 1.214654e-13, 
    1.215862e-13, 1.217405e-13, 1.217572e-13, 1.218486e-13, 1.216988e-13, 
    1.218427e-13, 1.21298e-13, 1.215415e-13, 1.208727e-13, 1.210356e-13, 
    1.209607e-13, 1.208785e-13, 1.211322e-13, 1.214021e-13, 1.21408e-13, 
    1.214945e-13, 1.217379e-13, 1.213192e-13, 1.226139e-13, 1.218148e-13, 
    1.206181e-13, 1.208642e-13, 1.208994e-13, 1.208041e-13, 1.214505e-13, 
    1.212164e-13, 1.218464e-13, 1.216763e-13, 1.219549e-13, 1.218165e-13, 
    1.217961e-13, 1.216182e-13, 1.215074e-13, 1.212271e-13, 1.20999e-13, 
    1.208179e-13, 1.208601e-13, 1.210589e-13, 1.214186e-13, 1.217587e-13, 
    1.216842e-13, 1.219338e-13, 1.212729e-13, 1.215501e-13, 1.21443e-13, 
    1.217223e-13, 1.2111e-13, 1.216312e-13, 1.209766e-13, 1.210341e-13, 
    1.212118e-13, 1.215689e-13, 1.21648e-13, 1.217322e-13, 1.216802e-13, 
    1.214278e-13, 1.213864e-13, 1.212075e-13, 1.21158e-13, 1.210215e-13, 
    1.209085e-13, 1.210118e-13, 1.211202e-13, 1.214279e-13, 1.21705e-13, 
    1.220067e-13, 1.220805e-13, 1.224324e-13, 1.221459e-13, 1.226183e-13, 
    1.222165e-13, 1.229118e-13, 1.216615e-13, 1.222049e-13, 1.212199e-13, 
    1.213262e-13, 1.215183e-13, 1.219585e-13, 1.21721e-13, 1.219988e-13, 
    1.213848e-13, 1.210657e-13, 1.209832e-13, 1.208289e-13, 1.209867e-13, 
    1.209739e-13, 1.211247e-13, 1.210763e-13, 1.214382e-13, 1.212438e-13, 
    1.217956e-13, 1.219966e-13, 1.225637e-13, 1.229107e-13, 1.232636e-13, 
    1.234192e-13, 1.234666e-13, 1.234864e-13 ;

 LITR3C =
  9.698032e-06, 9.698022e-06, 9.698025e-06, 9.698017e-06, 9.698021e-06, 
    9.698016e-06, 9.69803e-06, 9.698022e-06, 9.698027e-06, 9.698031e-06, 
    9.698001e-06, 9.698016e-06, 9.697986e-06, 9.697995e-06, 9.697971e-06, 
    9.697987e-06, 9.697967e-06, 9.697971e-06, 9.69796e-06, 9.697964e-06, 
    9.697949e-06, 9.697958e-06, 9.697942e-06, 9.697952e-06, 9.69795e-06, 
    9.697959e-06, 9.698013e-06, 9.698003e-06, 9.698014e-06, 9.698012e-06, 
    9.698013e-06, 9.698021e-06, 9.698025e-06, 9.698033e-06, 9.698031e-06, 
    9.698026e-06, 9.698011e-06, 9.698017e-06, 9.698005e-06, 9.698005e-06, 
    9.697991e-06, 9.697997e-06, 9.697976e-06, 9.697981e-06, 9.697963e-06, 
    9.697967e-06, 9.697964e-06, 9.697965e-06, 9.697964e-06, 9.69797e-06, 
    9.697967e-06, 9.697973e-06, 9.697997e-06, 9.697989e-06, 9.698009e-06, 
    9.698022e-06, 9.69803e-06, 9.698036e-06, 9.698035e-06, 9.698033e-06, 
    9.698026e-06, 9.698017e-06, 9.698012e-06, 9.698008e-06, 9.698005e-06, 
    9.697993e-06, 9.697987e-06, 9.697974e-06, 9.697977e-06, 9.697972e-06, 
    9.697968e-06, 9.697962e-06, 9.697963e-06, 9.69796e-06, 9.697972e-06, 
    9.697964e-06, 9.697977e-06, 9.697974e-06, 9.698004e-06, 9.698015e-06, 
    9.69802e-06, 9.698024e-06, 9.698034e-06, 9.698027e-06, 9.69803e-06, 
    9.698023e-06, 9.698019e-06, 9.698021e-06, 9.698008e-06, 9.698013e-06, 
    9.697987e-06, 9.697998e-06, 9.697968e-06, 9.697976e-06, 9.697967e-06, 
    9.697972e-06, 9.697964e-06, 9.697971e-06, 9.697959e-06, 9.697957e-06, 
    9.697958e-06, 9.697951e-06, 9.697971e-06, 9.697964e-06, 9.698021e-06, 
    9.698021e-06, 9.698019e-06, 9.698027e-06, 9.698027e-06, 9.698033e-06, 
    9.698027e-06, 9.698025e-06, 9.698019e-06, 9.698016e-06, 9.698012e-06, 
    9.698004e-06, 9.697996e-06, 9.697984e-06, 9.697976e-06, 9.697969e-06, 
    9.697973e-06, 9.69797e-06, 9.697974e-06, 9.697975e-06, 9.697957e-06, 
    9.697967e-06, 9.697952e-06, 9.697953e-06, 9.69796e-06, 9.697953e-06, 
    9.698021e-06, 9.698023e-06, 9.698029e-06, 9.698024e-06, 9.698034e-06, 
    9.698028e-06, 9.698026e-06, 9.698013e-06, 9.69801e-06, 9.698008e-06, 
    9.698003e-06, 9.697997e-06, 9.697987e-06, 9.697977e-06, 9.697968e-06, 
    9.697968e-06, 9.697968e-06, 9.697967e-06, 9.697971e-06, 9.697966e-06, 
    9.697965e-06, 9.697967e-06, 9.697953e-06, 9.697957e-06, 9.697953e-06, 
    9.697956e-06, 9.698022e-06, 9.698018e-06, 9.69802e-06, 9.698017e-06, 
    9.698019e-06, 9.698009e-06, 9.698006e-06, 9.697991e-06, 9.697997e-06, 
    9.697987e-06, 9.697997e-06, 9.697995e-06, 9.697987e-06, 9.697996e-06, 
    9.697977e-06, 9.69799e-06, 9.697967e-06, 9.697979e-06, 9.697966e-06, 
    9.697968e-06, 9.697964e-06, 9.69796e-06, 9.697956e-06, 9.697947e-06, 
    9.697949e-06, 9.697943e-06, 9.698014e-06, 9.698009e-06, 9.69801e-06, 
    9.698006e-06, 9.698002e-06, 9.697995e-06, 9.697984e-06, 9.697987e-06, 
    9.69798e-06, 9.697978e-06, 9.69799e-06, 9.697983e-06, 9.698007e-06, 
    9.698003e-06, 9.698005e-06, 9.698014e-06, 9.697987e-06, 9.698e-06, 
    9.697976e-06, 9.697983e-06, 9.697961e-06, 9.697972e-06, 9.697951e-06, 
    9.697942e-06, 9.697934e-06, 9.697924e-06, 9.698007e-06, 9.69801e-06, 
    9.698005e-06, 9.697997e-06, 9.697991e-06, 9.697982e-06, 9.697981e-06, 
    9.697979e-06, 9.697976e-06, 9.697972e-06, 9.697979e-06, 9.697971e-06, 
    9.698002e-06, 9.697986e-06, 9.698011e-06, 9.698004e-06, 9.697998e-06, 
    9.698e-06, 9.697988e-06, 9.697986e-06, 9.697974e-06, 9.69798e-06, 
    9.697944e-06, 9.69796e-06, 9.697916e-06, 9.697928e-06, 9.698011e-06, 
    9.698007e-06, 9.697994e-06, 9.698e-06, 9.697982e-06, 9.697977e-06, 
    9.697973e-06, 9.697968e-06, 9.697968e-06, 9.697966e-06, 9.69797e-06, 
    9.697966e-06, 9.697982e-06, 9.697975e-06, 9.697995e-06, 9.69799e-06, 
    9.697992e-06, 9.697995e-06, 9.697987e-06, 9.697979e-06, 9.697978e-06, 
    9.697977e-06, 9.697968e-06, 9.697981e-06, 9.697942e-06, 9.697967e-06, 
    9.698003e-06, 9.697996e-06, 9.697995e-06, 9.697997e-06, 9.697977e-06, 
    9.697985e-06, 9.697966e-06, 9.69797e-06, 9.697962e-06, 9.697967e-06, 
    9.697967e-06, 9.697972e-06, 9.697976e-06, 9.697985e-06, 9.697991e-06, 
    9.697997e-06, 9.697996e-06, 9.697989e-06, 9.697978e-06, 9.697968e-06, 
    9.69797e-06, 9.697963e-06, 9.697983e-06, 9.697975e-06, 9.697977e-06, 
    9.697969e-06, 9.697987e-06, 9.697972e-06, 9.697992e-06, 9.69799e-06, 
    9.697985e-06, 9.697974e-06, 9.697971e-06, 9.697969e-06, 9.69797e-06, 
    9.697978e-06, 9.697979e-06, 9.697985e-06, 9.697987e-06, 9.69799e-06, 
    9.697994e-06, 9.697991e-06, 9.697987e-06, 9.697978e-06, 9.69797e-06, 
    9.69796e-06, 9.697958e-06, 9.697947e-06, 9.697957e-06, 9.697942e-06, 
    9.697954e-06, 9.697933e-06, 9.697971e-06, 9.697955e-06, 9.697985e-06, 
    9.697981e-06, 9.697976e-06, 9.697962e-06, 9.697969e-06, 9.697961e-06, 
    9.697979e-06, 9.697989e-06, 9.697992e-06, 9.697997e-06, 9.697992e-06, 
    9.697992e-06, 9.697987e-06, 9.697989e-06, 9.697977e-06, 9.697984e-06, 
    9.697967e-06, 9.697961e-06, 9.697944e-06, 9.697933e-06, 9.697922e-06, 
    9.697917e-06, 9.697916e-06, 9.697916e-06 ;

 LITR3C_TO_SOIL2C =
  5.982752e-14, 5.998923e-14, 5.995782e-14, 6.008813e-14, 6.001588e-14, 
    6.010117e-14, 5.986034e-14, 5.999564e-14, 5.990929e-14, 5.984211e-14, 
    6.034062e-14, 6.009395e-14, 6.059662e-14, 6.043959e-14, 6.08338e-14, 
    6.057217e-14, 6.08865e-14, 6.08263e-14, 6.100752e-14, 6.095563e-14, 
    6.118706e-14, 6.103146e-14, 6.130695e-14, 6.114994e-14, 6.117449e-14, 
    6.102632e-14, 6.014367e-14, 6.030992e-14, 6.01338e-14, 6.015752e-14, 
    6.014689e-14, 6.001735e-14, 5.9952e-14, 5.981518e-14, 5.984005e-14, 
    5.994054e-14, 6.016819e-14, 6.009098e-14, 6.028558e-14, 6.028119e-14, 
    6.04975e-14, 6.040001e-14, 6.076313e-14, 6.066003e-14, 6.09578e-14, 
    6.088297e-14, 6.095427e-14, 6.093266e-14, 6.095456e-14, 6.08448e-14, 
    6.089183e-14, 6.079522e-14, 6.041826e-14, 6.052914e-14, 6.019818e-14, 
    5.999876e-14, 5.986627e-14, 5.977215e-14, 5.978546e-14, 5.981082e-14, 
    5.994113e-14, 6.006359e-14, 6.015683e-14, 6.021916e-14, 6.028056e-14, 
    6.046612e-14, 6.056434e-14, 6.078394e-14, 6.074438e-14, 6.081144e-14, 
    6.087552e-14, 6.0983e-14, 6.096532e-14, 6.101264e-14, 6.080969e-14, 
    6.094459e-14, 6.072183e-14, 6.078279e-14, 6.029708e-14, 6.011182e-14, 
    6.003287e-14, 5.996385e-14, 5.979569e-14, 5.991183e-14, 5.986605e-14, 
    5.997497e-14, 6.004412e-14, 6.000993e-14, 6.022086e-14, 6.013889e-14, 
    6.057016e-14, 6.038455e-14, 6.086805e-14, 6.07525e-14, 6.089573e-14, 
    6.082267e-14, 6.094782e-14, 6.083519e-14, 6.103026e-14, 6.107267e-14, 
    6.104369e-14, 6.115507e-14, 6.082895e-14, 6.095426e-14, 6.000896e-14, 
    6.001454e-14, 6.004053e-14, 5.992625e-14, 5.991926e-14, 5.98145e-14, 
    5.990773e-14, 5.994741e-14, 6.004814e-14, 6.010766e-14, 6.016423e-14, 
    6.028853e-14, 6.042721e-14, 6.062095e-14, 6.076e-14, 6.085312e-14, 
    6.079603e-14, 6.084644e-14, 6.079009e-14, 6.076368e-14, 6.105677e-14, 
    6.089226e-14, 6.113905e-14, 6.112541e-14, 6.101376e-14, 6.112695e-14, 
    6.001846e-14, 5.998637e-14, 5.987484e-14, 5.996213e-14, 5.980309e-14, 
    5.989211e-14, 5.994326e-14, 6.014057e-14, 6.018392e-14, 6.022406e-14, 
    6.030334e-14, 6.0405e-14, 6.058316e-14, 6.073802e-14, 6.087925e-14, 
    6.086891e-14, 6.087255e-14, 6.090407e-14, 6.082596e-14, 6.091689e-14, 
    6.093213e-14, 6.089226e-14, 6.112358e-14, 6.105754e-14, 6.112512e-14, 
    6.108213e-14, 5.99968e-14, 6.00508e-14, 6.002162e-14, 6.007648e-14, 
    6.003782e-14, 6.020959e-14, 6.026105e-14, 6.050164e-14, 6.040299e-14, 
    6.056001e-14, 6.041896e-14, 6.044395e-14, 6.056506e-14, 6.04266e-14, 
    6.072945e-14, 6.052413e-14, 6.090529e-14, 6.070045e-14, 6.091812e-14, 
    6.087864e-14, 6.094401e-14, 6.100251e-14, 6.10761e-14, 6.121174e-14, 
    6.118035e-14, 6.129373e-14, 6.013128e-14, 6.020123e-14, 6.019511e-14, 
    6.026831e-14, 6.032241e-14, 6.043965e-14, 6.062745e-14, 6.055687e-14, 
    6.068645e-14, 6.071244e-14, 6.051558e-14, 6.063645e-14, 6.024806e-14, 
    6.031085e-14, 6.027349e-14, 6.013678e-14, 6.057309e-14, 6.034932e-14, 
    6.076229e-14, 6.064127e-14, 6.099416e-14, 6.081875e-14, 6.116306e-14, 
    6.13099e-14, 6.144811e-14, 6.160927e-14, 6.023943e-14, 6.019191e-14, 
    6.027702e-14, 6.039463e-14, 6.050375e-14, 6.064865e-14, 6.066348e-14, 
    6.06906e-14, 6.076086e-14, 6.081989e-14, 6.069915e-14, 6.083469e-14, 
    6.032535e-14, 6.059252e-14, 6.017391e-14, 6.030005e-14, 6.038771e-14, 
    6.03493e-14, 6.05488e-14, 6.059577e-14, 6.078648e-14, 6.068795e-14, 
    6.127365e-14, 6.101482e-14, 6.173194e-14, 6.153191e-14, 6.017529e-14, 
    6.023928e-14, 6.046172e-14, 6.035593e-14, 6.065833e-14, 6.073266e-14, 
    6.079308e-14, 6.087023e-14, 6.087858e-14, 6.092426e-14, 6.084938e-14, 
    6.092132e-14, 6.064896e-14, 6.077074e-14, 6.043635e-14, 6.051779e-14, 
    6.048034e-14, 6.043922e-14, 6.056607e-14, 6.070104e-14, 6.070397e-14, 
    6.074721e-14, 6.086891e-14, 6.065956e-14, 6.130693e-14, 6.09074e-14, 
    6.030902e-14, 6.043207e-14, 6.044969e-14, 6.040203e-14, 6.072521e-14, 
    6.060819e-14, 6.092316e-14, 6.083811e-14, 6.097744e-14, 6.090822e-14, 
    6.089803e-14, 6.080908e-14, 6.075365e-14, 6.061355e-14, 6.049946e-14, 
    6.040895e-14, 6.043001e-14, 6.052941e-14, 6.07093e-14, 6.087931e-14, 
    6.084208e-14, 6.096686e-14, 6.063643e-14, 6.077505e-14, 6.072147e-14, 
    6.086115e-14, 6.055498e-14, 6.081559e-14, 6.048827e-14, 6.051701e-14, 
    6.060586e-14, 6.078442e-14, 6.082397e-14, 6.086609e-14, 6.084011e-14, 
    6.071388e-14, 6.069321e-14, 6.060372e-14, 6.057898e-14, 6.051076e-14, 
    6.045423e-14, 6.050587e-14, 6.056006e-14, 6.071395e-14, 6.085246e-14, 
    6.100333e-14, 6.104025e-14, 6.121616e-14, 6.107291e-14, 6.130914e-14, 
    6.110823e-14, 6.145589e-14, 6.083075e-14, 6.110242e-14, 6.060992e-14, 
    6.066308e-14, 6.075911e-14, 6.097923e-14, 6.086049e-14, 6.099937e-14, 
    6.06924e-14, 6.053282e-14, 6.049156e-14, 6.041445e-14, 6.049332e-14, 
    6.048691e-14, 6.056234e-14, 6.053811e-14, 6.071906e-14, 6.062189e-14, 
    6.089776e-14, 6.099828e-14, 6.128183e-14, 6.145533e-14, 6.163179e-14, 
    6.170959e-14, 6.173327e-14, 6.174316e-14 ;

 LITR3C_vr =
  0.0005537677, 0.0005537671, 0.0005537672, 0.0005537667, 0.000553767, 
    0.0005537667, 0.0005537675, 0.0005537671, 0.0005537674, 0.0005537676, 
    0.0005537659, 0.0005537667, 0.000553765, 0.0005537655, 0.0005537642, 
    0.000553765, 0.000553764, 0.0005537642, 0.0005537635, 0.0005537638, 
    0.0005537629, 0.0005537635, 0.0005537625, 0.0005537631, 0.0005537629, 
    0.0005537635, 0.0005537666, 0.000553766, 0.0005537666, 0.0005537665, 
    0.0005537666, 0.000553767, 0.0005537673, 0.0005537677, 0.0005537676, 
    0.0005537673, 0.0005537665, 0.0005537667, 0.0005537661, 0.0005537661, 
    0.0005537653, 0.0005537657, 0.0005537644, 0.0005537648, 0.0005537637, 
    0.000553764, 0.0005537638, 0.0005537638, 0.0005537638, 0.0005537641, 
    0.0005537639, 0.0005537643, 0.0005537656, 0.0005537652, 0.0005537664, 
    0.0005537671, 0.0005537675, 0.0005537678, 0.0005537678, 0.0005537677, 
    0.0005537673, 0.0005537668, 0.0005537665, 0.0005537663, 0.0005537661, 
    0.0005537655, 0.0005537651, 0.0005537643, 0.0005537645, 0.0005537642, 
    0.000553764, 0.0005537636, 0.0005537637, 0.0005537635, 0.0005537642, 
    0.0005537638, 0.0005537646, 0.0005537643, 0.000553766, 0.0005537667, 
    0.000553767, 0.0005537672, 0.0005537678, 0.0005537674, 0.0005537675, 
    0.0005537671, 0.0005537669, 0.000553767, 0.0005537663, 0.0005537666, 
    0.0005537651, 0.0005537657, 0.0005537641, 0.0005537645, 0.0005537639, 
    0.0005537642, 0.0005537638, 0.0005537642, 0.0005537635, 0.0005537634, 
    0.0005537634, 0.0005537631, 0.0005537642, 0.0005537638, 0.000553767, 
    0.000553767, 0.0005537669, 0.0005537673, 0.0005537674, 0.0005537677, 
    0.0005537674, 0.0005537673, 0.0005537669, 0.0005537667, 0.0005537665, 
    0.000553766, 0.0005537656, 0.0005537649, 0.0005537644, 0.0005537641, 
    0.0005537643, 0.0005537641, 0.0005537643, 0.0005537644, 0.0005537634, 
    0.0005537639, 0.0005537631, 0.0005537631, 0.0005537635, 0.0005537631, 
    0.000553767, 0.0005537671, 0.0005537675, 0.0005537672, 0.0005537678, 
    0.0005537674, 0.0005537673, 0.0005537666, 0.0005537664, 0.0005537663, 
    0.000553766, 0.0005537657, 0.000553765, 0.0005537645, 0.000553764, 
    0.0005537641, 0.000553764, 0.0005537639, 0.0005537642, 0.0005537639, 
    0.0005537638, 0.0005537639, 0.0005537631, 0.0005537634, 0.0005537631, 
    0.0005537633, 0.0005537671, 0.0005537669, 0.000553767, 0.0005537668, 
    0.0005537669, 0.0005537663, 0.0005537661, 0.0005537653, 0.0005537657, 
    0.0005537651, 0.0005537656, 0.0005537655, 0.0005537651, 0.0005537656, 
    0.0005537645, 0.0005537652, 0.0005537639, 0.0005537646, 0.0005537639, 
    0.000553764, 0.0005537638, 0.0005537636, 0.0005537633, 0.0005537628, 
    0.0005537629, 0.0005537625, 0.0005537666, 0.0005537664, 0.0005537664, 
    0.0005537661, 0.0005537659, 0.0005537655, 0.0005537649, 0.0005537651, 
    0.0005537647, 0.0005537646, 0.0005537653, 0.0005537649, 0.0005537662, 
    0.000553766, 0.0005537661, 0.0005537666, 0.000553765, 0.0005537659, 
    0.0005537644, 0.0005537648, 0.0005537636, 0.0005537642, 0.000553763, 
    0.0005537625, 0.000553762, 0.0005537614, 0.0005537662, 0.0005537664, 
    0.0005537661, 0.0005537657, 0.0005537653, 0.0005537648, 0.0005537648, 
    0.0005537646, 0.0005537644, 0.0005537642, 0.0005537646, 0.0005537642, 
    0.0005537659, 0.000553765, 0.0005537664, 0.000553766, 0.0005537657, 
    0.0005537659, 0.0005537652, 0.000553765, 0.0005537643, 0.0005537647, 
    0.0005537626, 0.0005537635, 0.000553761, 0.0005537617, 0.0005537664, 
    0.0005537662, 0.0005537655, 0.0005537658, 0.0005537648, 0.0005537645, 
    0.0005537643, 0.0005537641, 0.000553764, 0.0005537638, 0.0005537641, 
    0.0005537639, 0.0005537648, 0.0005537644, 0.0005537656, 0.0005537653, 
    0.0005537654, 0.0005537655, 0.0005537651, 0.0005537646, 0.0005537646, 
    0.0005537645, 0.0005537641, 0.0005537648, 0.0005537625, 0.0005537639, 
    0.000553766, 0.0005537656, 0.0005537655, 0.0005537657, 0.0005537645, 
    0.0005537649, 0.0005537638, 0.0005537642, 0.0005537636, 0.0005537639, 
    0.0005537639, 0.0005537642, 0.0005537645, 0.0005537649, 0.0005537653, 
    0.0005537656, 0.0005537656, 0.0005537652, 0.0005537646, 0.000553764, 
    0.0005537641, 0.0005537637, 0.0005537649, 0.0005537643, 0.0005537646, 
    0.0005537641, 0.0005537652, 0.0005537642, 0.0005537654, 0.0005537653, 
    0.0005537649, 0.0005537643, 0.0005537642, 0.0005537641, 0.0005537641, 
    0.0005537646, 0.0005537646, 0.000553765, 0.000553765, 0.0005537653, 
    0.0005537655, 0.0005537653, 0.0005537651, 0.0005537646, 0.0005537641, 
    0.0005537636, 0.0005537634, 0.0005537628, 0.0005537633, 0.0005537625, 
    0.0005537632, 0.000553762, 0.0005537642, 0.0005537632, 0.0005537649, 
    0.0005537648, 0.0005537644, 0.0005537636, 0.0005537641, 0.0005537636, 
    0.0005537646, 0.0005537652, 0.0005537653, 0.0005537656, 0.0005537653, 
    0.0005537654, 0.0005537651, 0.0005537652, 0.0005537646, 0.0005537649, 
    0.0005537639, 0.0005537636, 0.0005537626, 0.000553762, 0.0005537614, 
    0.0005537611, 0.000553761, 0.000553761,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342137e-07, 1.342135e-07, 1.342136e-07, 1.342135e-07, 1.342135e-07, 
    1.342134e-07, 1.342136e-07, 1.342135e-07, 1.342136e-07, 1.342137e-07, 
    1.342132e-07, 1.342135e-07, 1.34213e-07, 1.342132e-07, 1.342128e-07, 
    1.34213e-07, 1.342128e-07, 1.342128e-07, 1.342127e-07, 1.342127e-07, 
    1.342125e-07, 1.342127e-07, 1.342124e-07, 1.342126e-07, 1.342125e-07, 
    1.342127e-07, 1.342134e-07, 1.342133e-07, 1.342134e-07, 1.342134e-07, 
    1.342134e-07, 1.342135e-07, 1.342136e-07, 1.342137e-07, 1.342137e-07, 
    1.342136e-07, 1.342134e-07, 1.342135e-07, 1.342133e-07, 1.342133e-07, 
    1.342131e-07, 1.342132e-07, 1.342129e-07, 1.34213e-07, 1.342127e-07, 
    1.342128e-07, 1.342127e-07, 1.342127e-07, 1.342127e-07, 1.342128e-07, 
    1.342128e-07, 1.342129e-07, 1.342132e-07, 1.342131e-07, 1.342134e-07, 
    1.342135e-07, 1.342136e-07, 1.342137e-07, 1.342137e-07, 1.342137e-07, 
    1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 
    1.342131e-07, 1.342131e-07, 1.342129e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.342127e-07, 1.342127e-07, 1.342128e-07, 
    1.342127e-07, 1.342129e-07, 1.342129e-07, 1.342133e-07, 1.342134e-07, 
    1.342135e-07, 1.342136e-07, 1.342137e-07, 1.342136e-07, 1.342136e-07, 
    1.342136e-07, 1.342135e-07, 1.342135e-07, 1.342133e-07, 1.342134e-07, 
    1.34213e-07, 1.342132e-07, 1.342128e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.342128e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342125e-07, 1.342128e-07, 1.342127e-07, 1.342135e-07, 
    1.342135e-07, 1.342135e-07, 1.342136e-07, 1.342136e-07, 1.342137e-07, 
    1.342136e-07, 1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342134e-07, 
    1.342133e-07, 1.342132e-07, 1.34213e-07, 1.342129e-07, 1.342128e-07, 
    1.342129e-07, 1.342128e-07, 1.342129e-07, 1.342129e-07, 1.342126e-07, 
    1.342128e-07, 1.342126e-07, 1.342126e-07, 1.342127e-07, 1.342126e-07, 
    1.342135e-07, 1.342135e-07, 1.342136e-07, 1.342136e-07, 1.342137e-07, 
    1.342136e-07, 1.342136e-07, 1.342134e-07, 1.342134e-07, 1.342133e-07, 
    1.342133e-07, 1.342132e-07, 1.34213e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342128e-07, 1.342128e-07, 1.342128e-07, 1.342128e-07, 
    1.342127e-07, 1.342128e-07, 1.342126e-07, 1.342126e-07, 1.342126e-07, 
    1.342126e-07, 1.342135e-07, 1.342135e-07, 1.342135e-07, 1.342135e-07, 
    1.342135e-07, 1.342134e-07, 1.342133e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 
    1.342129e-07, 1.342131e-07, 1.342128e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 
    1.342125e-07, 1.342124e-07, 1.342134e-07, 1.342134e-07, 1.342134e-07, 
    1.342133e-07, 1.342133e-07, 1.342132e-07, 1.34213e-07, 1.342131e-07, 
    1.342129e-07, 1.342129e-07, 1.342131e-07, 1.34213e-07, 1.342133e-07, 
    1.342133e-07, 1.342133e-07, 1.342134e-07, 1.34213e-07, 1.342132e-07, 
    1.342129e-07, 1.34213e-07, 1.342127e-07, 1.342128e-07, 1.342125e-07, 
    1.342124e-07, 1.342123e-07, 1.342122e-07, 1.342133e-07, 1.342134e-07, 
    1.342133e-07, 1.342132e-07, 1.342131e-07, 1.34213e-07, 1.34213e-07, 
    1.342129e-07, 1.342129e-07, 1.342128e-07, 1.342129e-07, 1.342128e-07, 
    1.342133e-07, 1.34213e-07, 1.342134e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342124e-07, 1.342127e-07, 1.342121e-07, 1.342122e-07, 1.342134e-07, 
    1.342133e-07, 1.342131e-07, 1.342132e-07, 1.34213e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.342128e-07, 1.342127e-07, 1.342128e-07, 
    1.342127e-07, 1.34213e-07, 1.342129e-07, 1.342132e-07, 1.342131e-07, 
    1.342131e-07, 1.342132e-07, 1.342131e-07, 1.342129e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.34213e-07, 1.342124e-07, 1.342128e-07, 
    1.342133e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 1.342129e-07, 
    1.34213e-07, 1.342127e-07, 1.342128e-07, 1.342127e-07, 1.342128e-07, 
    1.342128e-07, 1.342128e-07, 1.342129e-07, 1.34213e-07, 1.342131e-07, 
    1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342131e-07, 1.342128e-07, 1.342131e-07, 1.342131e-07, 
    1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342128e-07, 1.342128e-07, 
    1.342129e-07, 1.342129e-07, 1.34213e-07, 1.34213e-07, 1.342131e-07, 
    1.342131e-07, 1.342131e-07, 1.342131e-07, 1.342129e-07, 1.342128e-07, 
    1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342126e-07, 1.342124e-07, 
    1.342126e-07, 1.342123e-07, 1.342128e-07, 1.342126e-07, 1.34213e-07, 
    1.34213e-07, 1.342129e-07, 1.342127e-07, 1.342128e-07, 1.342127e-07, 
    1.342129e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 
    1.342131e-07, 1.342131e-07, 1.342131e-07, 1.342129e-07, 1.34213e-07, 
    1.342128e-07, 1.342127e-07, 1.342124e-07, 1.342123e-07, 1.342121e-07, 
    1.342121e-07, 1.342121e-07, 1.34212e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  -1.446034e-25, -7.652491e-42, 2.450906e-27, -4.65672e-26, 3.431268e-26, 
    6.98508e-26, 7.652491e-42, -4.65672e-26, -5.269447e-26, 2.08327e-26, 
    4.41163e-26, 1.225453e-27, 1.225453e-26, 7.352717e-26, -2.695996e-26, 
    -1.593089e-26, 9.926167e-26, -4.289085e-26, -2.695996e-26, 1.225453e-27, 
    -7.652491e-42, 4.043994e-26, -4.41163e-26, -3.186177e-26, 2.941087e-26, 
    -1.715634e-26, 4.41163e-26, -5.882173e-26, -7.965443e-26, -1.593089e-26, 
    2.695996e-26, 1.225453e-25, -1.225453e-26, 4.41163e-26, 6.249809e-26, 
    -7.230172e-26, -7.475262e-26, 9.803622e-27, 2.450905e-26, -4.289085e-26, 
    -6.4949e-26, 5.759628e-26, 1.249962e-25, -4.65672e-26, 2.450906e-27, 
    -8.333079e-26, 7.475262e-26, 9.068351e-26, -5.637083e-26, -7.965443e-26, 
    -7.352717e-27, 3.553813e-26, -6.127264e-27, -1.200944e-25, 5.637083e-26, 
    7.720352e-26, -3.063632e-26, -6.73999e-26, 7.352717e-27, -4.534175e-26, 
    -1.225453e-26, -4.901811e-26, 5.146902e-26, 3.676358e-26, 7.352717e-26, 
    9.313441e-26, 6.249809e-26, 1.017126e-25, 3.798904e-26, 1.519561e-25, 
    -1.642107e-25, -3.553813e-26, -1.225453e-26, -2.205815e-26, 
    -6.372354e-26, 2.941087e-26, -6.127264e-26, -1.838179e-26, -7.597807e-26, 
    -9.803622e-26, -6.73999e-26, 9.313441e-26, 8.210533e-26, 1.102908e-26, 
    -4.289085e-26, 8.210533e-26, -1.02938e-25, -4.65672e-26, -7.720352e-26, 
    -7.107626e-26, -9.803622e-27, -1.225453e-26, 1.225453e-27, -3.431268e-26, 
    -8.333079e-26, -1.225453e-27, -3.431268e-26, -3.308722e-26, 
    -5.024356e-26, 6.127264e-26, -9.068351e-26, -8.087988e-26, 1.372507e-25, 
    3.676358e-26, -1.02938e-25, -2.08327e-26, -1.102908e-26, -6.4949e-26, 
    -7.597807e-26, -2.205815e-26, -6.862535e-26, 8.82326e-26, 1.838179e-26, 
    3.553813e-26, 3.676358e-27, -1.311234e-25, -3.798904e-26, 6.617445e-26, 
    6.127264e-27, -1.347998e-26, 2.08327e-26, -6.4949e-26, -1.225453e-26, 
    -1.593089e-26, 5.882173e-26, -6.372354e-26, -1.004871e-25, -4.779266e-26, 
    -1.960724e-26, 5.146902e-26, -7.720352e-26, -8.700715e-26, 1.838179e-26, 
    -1.225453e-27, 4.65672e-26, 1.102908e-26, -7.475262e-26, 8.700715e-26, 
    1.225453e-27, 3.798904e-26, -8.087988e-26, -6.249809e-26, -9.435986e-26, 
    -1.115162e-25, 1.470543e-26, 6.004719e-26, 2.08327e-26, 6.127264e-27, 
    -5.269447e-26, 2.695996e-26, -6.617445e-26, -6.372354e-26, -2.450906e-27, 
    8.333079e-26, -4.65672e-26, 1.715634e-26, 6.127264e-27, -2.818541e-26, 
    -2.32836e-26, 1.507307e-25, -4.901811e-27, 1.102908e-26, -1.225453e-27, 
    5.882173e-26, -1.715634e-26, -3.921449e-26, -1.176435e-25, -2.695996e-26, 
    -2.695996e-26, -2.695996e-26, -3.063632e-26, 7.352717e-27, -3.431268e-26, 
    9.681077e-26, 1.470543e-26, 1.225453e-27, 6.4949e-26, -7.475262e-26, 
    -8.700715e-26, -7.352717e-27, 4.901811e-27, 3.676358e-27, 8.578169e-26, 
    -9.803622e-26, 1.593089e-26, -8.82326e-26, 9.803622e-27, -5.024356e-26, 
    -5.024356e-26, 1.02938e-25, -1.960724e-26, 3.676358e-27, 2.08327e-26, 
    4.41163e-26, -6.617445e-26, 1.225453e-27, 2.450905e-26, -3.553813e-26, 
    -4.534175e-26, 1.066144e-25, 7.230172e-26, 6.98508e-26, -1.127417e-25, 
    2.818541e-26, 3.063632e-26, -3.186177e-26, 2.205815e-26, 1.347998e-26, 
    -8.210533e-26, -8.578169e-27, -4.41163e-26, 3.676358e-26, -1.066144e-25, 
    -3.186177e-26, -2.695996e-26, 1.225453e-27, 8.578169e-27, 7.597807e-26, 
    -1.997488e-25, -3.676358e-27, 3.431268e-26, 1.102908e-26, -2.818541e-26, 
    4.779266e-26, -6.127264e-27, 2.941087e-26, -3.431268e-26, 2.205815e-26, 
    4.65672e-26, 5.882173e-26, -3.431268e-26, 4.534175e-26, -6.4949e-26, 
    6.617445e-26, -1.225453e-27, 8.455624e-26, 4.534175e-26, -5.759628e-26, 
    1.43378e-25, 2.205815e-26, 6.372354e-26, -5.637083e-26, 1.213198e-25, 
    -4.901811e-26, -1.850434e-25, -1.715634e-26, -7.720352e-26, 3.063632e-26, 
    -8.945805e-26, 4.41163e-26, -2.536687e-25, 5.146902e-26, -8.700715e-26, 
    7.965443e-26, 5.391992e-26, 2.205815e-26, -4.166539e-26, -1.347998e-26, 
    1.200944e-25, 1.960724e-26, -6.249809e-26, 7.720352e-26, -3.676358e-27, 
    1.593089e-26, -6.98508e-26, -3.431268e-26, -1.225453e-27, -5.637083e-26, 
    6.73999e-26, 1.715634e-25, 1.225453e-27, -7.842898e-26, 5.024356e-26, 
    1.838179e-26, 6.4949e-26, 7.352717e-26, -2.205815e-26, 1.262216e-25, 
    -1.16418e-25, -1.188689e-25, 3.553813e-26, 1.482798e-25, 9.803622e-27, 
    4.534175e-26, -4.043994e-26, 5.146902e-26, 9.803622e-27, 3.553813e-26, 
    -7.842898e-26, -1.249962e-25, 8.945805e-26, -2.32836e-26, -9.558531e-26, 
    4.534175e-26, 6.372354e-26, -3.798904e-26, 1.347998e-25, 2.941087e-26, 
    -3.431268e-26, 1.519561e-25, 7.652491e-42, 4.166539e-26, 2.205815e-26, 
    7.720352e-26, 2.695996e-26, 1.004871e-25, 6.4949e-26, 5.391992e-26, 
    -8.087988e-26, -6.249809e-26, 2.438651e-25, -6.372354e-26, 1.139671e-25, 
    7.965443e-26, 8.700715e-26, 1.347998e-26, -3.676358e-26, 5.269447e-26, 
    -5.024356e-26, 1.666616e-25, -8.578169e-27, 1.593089e-26, -4.901811e-26, 
    1.053889e-25, 1.593089e-26, 1.225453e-26, 7.352717e-27, -6.004719e-26, 
    -3.676358e-27, -9.681077e-26, 4.901811e-26, 4.779266e-26, -3.186177e-26, 
    1.066144e-25, -7.230172e-26, -1.960724e-26, -8.333079e-26, 7.352717e-27,
  1.33813e-32, 1.338128e-32, 1.338129e-32, 1.338128e-32, 1.338128e-32, 
    1.338128e-32, 1.33813e-32, 1.338128e-32, 1.338129e-32, 1.33813e-32, 
    1.338125e-32, 1.338128e-32, 1.338123e-32, 1.338125e-32, 1.338121e-32, 
    1.338124e-32, 1.338121e-32, 1.338121e-32, 1.33812e-32, 1.33812e-32, 
    1.338118e-32, 1.33812e-32, 1.338117e-32, 1.338119e-32, 1.338118e-32, 
    1.33812e-32, 1.338127e-32, 1.338126e-32, 1.338127e-32, 1.338127e-32, 
    1.338127e-32, 1.338128e-32, 1.338129e-32, 1.33813e-32, 1.33813e-32, 
    1.338129e-32, 1.338127e-32, 1.338128e-32, 1.338126e-32, 1.338126e-32, 
    1.338124e-32, 1.338125e-32, 1.338122e-32, 1.338123e-32, 1.33812e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 1.338121e-32, 
    1.338121e-32, 1.338122e-32, 1.338125e-32, 1.338124e-32, 1.338127e-32, 
    1.338128e-32, 1.33813e-32, 1.33813e-32, 1.33813e-32, 1.33813e-32, 
    1.338129e-32, 1.338128e-32, 1.338127e-32, 1.338126e-32, 1.338126e-32, 
    1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 1.338121e-32, 
    1.33812e-32, 1.338122e-32, 1.338122e-32, 1.338126e-32, 1.338127e-32, 
    1.338128e-32, 1.338129e-32, 1.33813e-32, 1.338129e-32, 1.33813e-32, 
    1.338129e-32, 1.338128e-32, 1.338128e-32, 1.338126e-32, 1.338127e-32, 
    1.338124e-32, 1.338125e-32, 1.338121e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.338121e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338119e-32, 1.338121e-32, 1.33812e-32, 1.338128e-32, 
    1.338128e-32, 1.338128e-32, 1.338129e-32, 1.338129e-32, 1.33813e-32, 
    1.338129e-32, 1.338129e-32, 1.338128e-32, 1.338128e-32, 1.338127e-32, 
    1.338126e-32, 1.338125e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 
    1.338122e-32, 1.338121e-32, 1.338122e-32, 1.338122e-32, 1.338119e-32, 
    1.338121e-32, 1.338119e-32, 1.338119e-32, 1.33812e-32, 1.338119e-32, 
    1.338128e-32, 1.338129e-32, 1.338129e-32, 1.338129e-32, 1.33813e-32, 
    1.338129e-32, 1.338129e-32, 1.338127e-32, 1.338127e-32, 1.338126e-32, 
    1.338126e-32, 1.338125e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.338121e-32, 1.338121e-32, 1.338121e-32, 1.338121e-32, 
    1.33812e-32, 1.338121e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 
    1.338119e-32, 1.338128e-32, 1.338128e-32, 1.338128e-32, 1.338128e-32, 
    1.338128e-32, 1.338127e-32, 1.338126e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 
    1.338122e-32, 1.338124e-32, 1.338121e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 
    1.338118e-32, 1.338117e-32, 1.338127e-32, 1.338127e-32, 1.338127e-32, 
    1.338126e-32, 1.338126e-32, 1.338125e-32, 1.338123e-32, 1.338124e-32, 
    1.338123e-32, 1.338122e-32, 1.338124e-32, 1.338123e-32, 1.338126e-32, 
    1.338126e-32, 1.338126e-32, 1.338127e-32, 1.338124e-32, 1.338125e-32, 
    1.338122e-32, 1.338123e-32, 1.33812e-32, 1.338121e-32, 1.338119e-32, 
    1.338117e-32, 1.338116e-32, 1.338115e-32, 1.338126e-32, 1.338127e-32, 
    1.338126e-32, 1.338125e-32, 1.338124e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338122e-32, 1.338121e-32, 1.338122e-32, 1.338121e-32, 
    1.338126e-32, 1.338123e-32, 1.338127e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338123e-32, 
    1.338118e-32, 1.33812e-32, 1.338114e-32, 1.338115e-32, 1.338127e-32, 
    1.338126e-32, 1.338124e-32, 1.338125e-32, 1.338123e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.338121e-32, 1.33812e-32, 1.338121e-32, 
    1.338121e-32, 1.338123e-32, 1.338122e-32, 1.338125e-32, 1.338124e-32, 
    1.338124e-32, 1.338125e-32, 1.338124e-32, 1.338122e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.338123e-32, 1.338117e-32, 1.338121e-32, 
    1.338126e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 1.338122e-32, 
    1.338123e-32, 1.33812e-32, 1.338121e-32, 1.33812e-32, 1.338121e-32, 
    1.338121e-32, 1.338121e-32, 1.338122e-32, 1.338123e-32, 1.338124e-32, 
    1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.338123e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.338124e-32, 1.338121e-32, 1.338124e-32, 1.338124e-32, 
    1.338123e-32, 1.338122e-32, 1.338121e-32, 1.338121e-32, 1.338121e-32, 
    1.338122e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 1.338124e-32, 
    1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338121e-32, 
    1.33812e-32, 1.33812e-32, 1.338118e-32, 1.338119e-32, 1.338117e-32, 
    1.338119e-32, 1.338116e-32, 1.338121e-32, 1.338119e-32, 1.338123e-32, 
    1.338123e-32, 1.338122e-32, 1.33812e-32, 1.338121e-32, 1.33812e-32, 
    1.338123e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 
    1.338124e-32, 1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338123e-32, 
    1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338116e-32, 1.338114e-32, 
    1.338114e-32, 1.338114e-32, 1.338114e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.655938e-15, 1.660414e-15, 1.659545e-15, 1.663152e-15, 1.661152e-15, 
    1.663512e-15, 1.656847e-15, 1.660591e-15, 1.658202e-15, 1.656342e-15, 
    1.67014e-15, 1.663312e-15, 1.677226e-15, 1.672879e-15, 1.68379e-15, 
    1.676549e-15, 1.685249e-15, 1.683583e-15, 1.688599e-15, 1.687163e-15, 
    1.693568e-15, 1.689262e-15, 1.696887e-15, 1.692541e-15, 1.693221e-15, 
    1.689119e-15, 1.664689e-15, 1.66929e-15, 1.664416e-15, 1.665072e-15, 
    1.664778e-15, 1.661193e-15, 1.659384e-15, 1.655597e-15, 1.656285e-15, 
    1.659066e-15, 1.665367e-15, 1.663231e-15, 1.668617e-15, 1.668495e-15, 
    1.674482e-15, 1.671784e-15, 1.681835e-15, 1.678981e-15, 1.687223e-15, 
    1.685151e-15, 1.687125e-15, 1.686527e-15, 1.687133e-15, 1.684095e-15, 
    1.685397e-15, 1.682723e-15, 1.672289e-15, 1.675358e-15, 1.666198e-15, 
    1.660678e-15, 1.657011e-15, 1.654406e-15, 1.654774e-15, 1.655476e-15, 
    1.659083e-15, 1.662472e-15, 1.665053e-15, 1.666778e-15, 1.668478e-15, 
    1.673614e-15, 1.676332e-15, 1.682411e-15, 1.681316e-15, 1.683171e-15, 
    1.684945e-15, 1.68792e-15, 1.687431e-15, 1.68874e-15, 1.683123e-15, 
    1.686857e-15, 1.680691e-15, 1.682379e-15, 1.668935e-15, 1.663807e-15, 
    1.661622e-15, 1.659712e-15, 1.655057e-15, 1.658272e-15, 1.657005e-15, 
    1.66002e-15, 1.661933e-15, 1.660987e-15, 1.666825e-15, 1.664556e-15, 
    1.676493e-15, 1.671356e-15, 1.684738e-15, 1.681541e-15, 1.685505e-15, 
    1.683483e-15, 1.686946e-15, 1.683829e-15, 1.689228e-15, 1.690402e-15, 
    1.6896e-15, 1.692683e-15, 1.683656e-15, 1.687125e-15, 1.66096e-15, 
    1.661115e-15, 1.661834e-15, 1.658671e-15, 1.658477e-15, 1.655578e-15, 
    1.658158e-15, 1.659257e-15, 1.662045e-15, 1.663692e-15, 1.665258e-15, 
    1.668698e-15, 1.672537e-15, 1.677899e-15, 1.681748e-15, 1.684325e-15, 
    1.682745e-15, 1.68414e-15, 1.682581e-15, 1.68185e-15, 1.689962e-15, 
    1.685409e-15, 1.69224e-15, 1.691862e-15, 1.688772e-15, 1.691905e-15, 
    1.661223e-15, 1.660335e-15, 1.657248e-15, 1.659664e-15, 1.655262e-15, 
    1.657726e-15, 1.659142e-15, 1.664603e-15, 1.665803e-15, 1.666914e-15, 
    1.669108e-15, 1.671922e-15, 1.676853e-15, 1.681139e-15, 1.685049e-15, 
    1.684763e-15, 1.684863e-15, 1.685736e-15, 1.683574e-15, 1.68609e-15, 
    1.686512e-15, 1.685409e-15, 1.691811e-15, 1.689983e-15, 1.691854e-15, 
    1.690664e-15, 1.660624e-15, 1.662118e-15, 1.661311e-15, 1.662829e-15, 
    1.661759e-15, 1.666513e-15, 1.667938e-15, 1.674597e-15, 1.671866e-15, 
    1.676212e-15, 1.672308e-15, 1.673e-15, 1.676352e-15, 1.67252e-15, 
    1.680902e-15, 1.675219e-15, 1.685769e-15, 1.6801e-15, 1.686124e-15, 
    1.685032e-15, 1.686841e-15, 1.68846e-15, 1.690497e-15, 1.694251e-15, 
    1.693383e-15, 1.696521e-15, 1.664346e-15, 1.666282e-15, 1.666112e-15, 
    1.668139e-15, 1.669636e-15, 1.672881e-15, 1.678079e-15, 1.676125e-15, 
    1.679712e-15, 1.680432e-15, 1.674983e-15, 1.678328e-15, 1.667578e-15, 
    1.669316e-15, 1.668282e-15, 1.664498e-15, 1.676575e-15, 1.670381e-15, 
    1.681811e-15, 1.678462e-15, 1.688229e-15, 1.683374e-15, 1.692904e-15, 
    1.696968e-15, 1.700794e-15, 1.705254e-15, 1.667339e-15, 1.666024e-15, 
    1.66838e-15, 1.671635e-15, 1.674655e-15, 1.678666e-15, 1.679076e-15, 
    1.679827e-15, 1.681772e-15, 1.683405e-15, 1.680064e-15, 1.683815e-15, 
    1.669717e-15, 1.677112e-15, 1.665526e-15, 1.669017e-15, 1.671443e-15, 
    1.67038e-15, 1.675902e-15, 1.677202e-15, 1.682481e-15, 1.679754e-15, 
    1.695965e-15, 1.688801e-15, 1.70865e-15, 1.703113e-15, 1.665564e-15, 
    1.667335e-15, 1.673492e-15, 1.670564e-15, 1.678934e-15, 1.680991e-15, 
    1.682663e-15, 1.684799e-15, 1.68503e-15, 1.686294e-15, 1.684222e-15, 
    1.686213e-15, 1.678674e-15, 1.682045e-15, 1.67279e-15, 1.675044e-15, 
    1.674007e-15, 1.672869e-15, 1.67638e-15, 1.680116e-15, 1.680197e-15, 
    1.681394e-15, 1.684762e-15, 1.678968e-15, 1.696886e-15, 1.685828e-15, 
    1.669266e-15, 1.672671e-15, 1.673159e-15, 1.67184e-15, 1.680785e-15, 
    1.677546e-15, 1.686264e-15, 1.68391e-15, 1.687766e-15, 1.68585e-15, 
    1.685568e-15, 1.683106e-15, 1.681572e-15, 1.677694e-15, 1.674537e-15, 
    1.672031e-15, 1.672614e-15, 1.675366e-15, 1.680345e-15, 1.68505e-15, 
    1.68402e-15, 1.687473e-15, 1.678328e-15, 1.682165e-15, 1.680682e-15, 
    1.684547e-15, 1.676073e-15, 1.683287e-15, 1.674227e-15, 1.675022e-15, 
    1.677482e-15, 1.682424e-15, 1.683518e-15, 1.684684e-15, 1.683965e-15, 
    1.680471e-15, 1.679899e-15, 1.677422e-15, 1.676738e-15, 1.674849e-15, 
    1.673285e-15, 1.674714e-15, 1.676214e-15, 1.680473e-15, 1.684307e-15, 
    1.688483e-15, 1.689505e-15, 1.694374e-15, 1.690409e-15, 1.696947e-15, 
    1.691386e-15, 1.701009e-15, 1.683706e-15, 1.691225e-15, 1.677594e-15, 
    1.679065e-15, 1.681723e-15, 1.687816e-15, 1.684529e-15, 1.688373e-15, 
    1.679877e-15, 1.67546e-15, 1.674318e-15, 1.672184e-15, 1.674367e-15, 
    1.674189e-15, 1.676277e-15, 1.675606e-15, 1.680615e-15, 1.677925e-15, 
    1.685561e-15, 1.688343e-15, 1.696191e-15, 1.700994e-15, 1.705878e-15, 
    1.708031e-15, 1.708686e-15, 1.70896e-15 ;

 LITR3N_vr =
  7.66374e-06, 7.663732e-06, 7.663733e-06, 7.663727e-06, 7.663731e-06, 
    7.663726e-06, 7.663738e-06, 7.663732e-06, 7.663735e-06, 7.663739e-06, 
    7.663714e-06, 7.663726e-06, 7.663702e-06, 7.66371e-06, 7.663691e-06, 
    7.663703e-06, 7.663688e-06, 7.663691e-06, 7.663682e-06, 7.663685e-06, 
    7.663673e-06, 7.663682e-06, 7.663668e-06, 7.663675e-06, 7.663674e-06, 
    7.663682e-06, 7.663724e-06, 7.663716e-06, 7.663724e-06, 7.663723e-06, 
    7.663724e-06, 7.66373e-06, 7.663733e-06, 7.66374e-06, 7.663739e-06, 
    7.663734e-06, 7.663722e-06, 7.663727e-06, 7.663717e-06, 7.663717e-06, 
    7.663707e-06, 7.663712e-06, 7.663694e-06, 7.663699e-06, 7.663684e-06, 
    7.663688e-06, 7.663685e-06, 7.663686e-06, 7.663685e-06, 7.66369e-06, 
    7.663688e-06, 7.663692e-06, 7.663711e-06, 7.663705e-06, 7.663722e-06, 
    7.663731e-06, 7.663737e-06, 7.663742e-06, 7.663742e-06, 7.66374e-06, 
    7.663733e-06, 7.663728e-06, 7.663723e-06, 7.663721e-06, 7.663717e-06, 
    7.663709e-06, 7.663703e-06, 7.663693e-06, 7.663695e-06, 7.663692e-06, 
    7.663689e-06, 7.663683e-06, 7.663684e-06, 7.663682e-06, 7.663692e-06, 
    7.663685e-06, 7.663696e-06, 7.663693e-06, 7.663717e-06, 7.663725e-06, 
    7.66373e-06, 7.663733e-06, 7.663741e-06, 7.663735e-06, 7.663737e-06, 
    7.663733e-06, 7.663729e-06, 7.663731e-06, 7.663721e-06, 7.663724e-06, 
    7.663703e-06, 7.663712e-06, 7.663689e-06, 7.663694e-06, 7.663688e-06, 
    7.663692e-06, 7.663685e-06, 7.663691e-06, 7.663682e-06, 7.663679e-06, 
    7.663681e-06, 7.663675e-06, 7.663691e-06, 7.663685e-06, 7.663731e-06, 
    7.663731e-06, 7.663729e-06, 7.663734e-06, 7.663735e-06, 7.66374e-06, 
    7.663735e-06, 7.663733e-06, 7.663729e-06, 7.663726e-06, 7.663723e-06, 
    7.663717e-06, 7.663711e-06, 7.663701e-06, 7.663694e-06, 7.66369e-06, 
    7.663692e-06, 7.66369e-06, 7.663692e-06, 7.663694e-06, 7.66368e-06, 
    7.663688e-06, 7.663676e-06, 7.663677e-06, 7.663682e-06, 7.663676e-06, 
    7.66373e-06, 7.663732e-06, 7.663737e-06, 7.663733e-06, 7.663741e-06, 
    7.663736e-06, 7.663733e-06, 7.663724e-06, 7.663722e-06, 7.66372e-06, 
    7.663716e-06, 7.663712e-06, 7.663702e-06, 7.663695e-06, 7.663689e-06, 
    7.663689e-06, 7.663689e-06, 7.663687e-06, 7.663691e-06, 7.663687e-06, 
    7.663686e-06, 7.663688e-06, 7.663677e-06, 7.66368e-06, 7.663677e-06, 
    7.663679e-06, 7.663732e-06, 7.663729e-06, 7.66373e-06, 7.663727e-06, 
    7.663729e-06, 7.663721e-06, 7.663718e-06, 7.663707e-06, 7.663712e-06, 
    7.663704e-06, 7.663711e-06, 7.66371e-06, 7.663703e-06, 7.663711e-06, 
    7.663696e-06, 7.663706e-06, 7.663687e-06, 7.663697e-06, 7.663687e-06, 
    7.663689e-06, 7.663685e-06, 7.663682e-06, 7.663679e-06, 7.663672e-06, 
    7.663674e-06, 7.663669e-06, 7.663724e-06, 7.663722e-06, 7.663722e-06, 
    7.663718e-06, 7.663715e-06, 7.66371e-06, 7.663701e-06, 7.663704e-06, 
    7.663698e-06, 7.663697e-06, 7.663706e-06, 7.663701e-06, 7.663719e-06, 
    7.663716e-06, 7.663718e-06, 7.663724e-06, 7.663703e-06, 7.663714e-06, 
    7.663694e-06, 7.6637e-06, 7.663683e-06, 7.663692e-06, 7.663675e-06, 
    7.663668e-06, 7.663661e-06, 7.663653e-06, 7.66372e-06, 7.663722e-06, 
    7.663718e-06, 7.663712e-06, 7.663707e-06, 7.6637e-06, 7.663699e-06, 
    7.663698e-06, 7.663694e-06, 7.663692e-06, 7.663697e-06, 7.663691e-06, 
    7.663715e-06, 7.663702e-06, 7.663722e-06, 7.663716e-06, 7.663712e-06, 
    7.663714e-06, 7.663704e-06, 7.663702e-06, 7.663693e-06, 7.663698e-06, 
    7.66367e-06, 7.663682e-06, 7.663647e-06, 7.663657e-06, 7.663722e-06, 
    7.66372e-06, 7.663709e-06, 7.663713e-06, 7.663699e-06, 7.663695e-06, 
    7.663692e-06, 7.663689e-06, 7.663689e-06, 7.663686e-06, 7.66369e-06, 
    7.663686e-06, 7.6637e-06, 7.663693e-06, 7.66371e-06, 7.663706e-06, 
    7.663708e-06, 7.66371e-06, 7.663703e-06, 7.663697e-06, 7.663697e-06, 
    7.663695e-06, 7.663689e-06, 7.663699e-06, 7.663668e-06, 7.663687e-06, 
    7.663716e-06, 7.66371e-06, 7.663709e-06, 7.663712e-06, 7.663696e-06, 
    7.663702e-06, 7.663686e-06, 7.663691e-06, 7.663683e-06, 7.663687e-06, 
    7.663688e-06, 7.663692e-06, 7.663694e-06, 7.663702e-06, 7.663707e-06, 
    7.663712e-06, 7.663711e-06, 7.663705e-06, 7.663697e-06, 7.663689e-06, 
    7.663691e-06, 7.663684e-06, 7.663701e-06, 7.663693e-06, 7.663696e-06, 
    7.66369e-06, 7.663704e-06, 7.663692e-06, 7.663707e-06, 7.663706e-06, 
    7.663702e-06, 7.663693e-06, 7.663692e-06, 7.663689e-06, 7.663691e-06, 
    7.663696e-06, 7.663698e-06, 7.663702e-06, 7.663703e-06, 7.663706e-06, 
    7.663709e-06, 7.663706e-06, 7.663704e-06, 7.663696e-06, 7.66369e-06, 
    7.663682e-06, 7.663681e-06, 7.663672e-06, 7.663679e-06, 7.663668e-06, 
    7.663677e-06, 7.663661e-06, 7.663691e-06, 7.663678e-06, 7.663702e-06, 
    7.663699e-06, 7.663694e-06, 7.663683e-06, 7.66369e-06, 7.663682e-06, 
    7.663698e-06, 7.663705e-06, 7.663707e-06, 7.663711e-06, 7.663707e-06, 
    7.663708e-06, 7.663703e-06, 7.663705e-06, 7.663696e-06, 7.663701e-06, 
    7.663688e-06, 7.663682e-06, 7.663669e-06, 7.663661e-06, 7.663652e-06, 
    7.663649e-06, 7.663647e-06, 7.663647e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.982752e-14, 5.998923e-14, 5.995782e-14, 6.008813e-14, 6.001588e-14, 
    6.010117e-14, 5.986034e-14, 5.999564e-14, 5.990929e-14, 5.984211e-14, 
    6.034062e-14, 6.009395e-14, 6.059662e-14, 6.043959e-14, 6.08338e-14, 
    6.057217e-14, 6.08865e-14, 6.08263e-14, 6.100752e-14, 6.095563e-14, 
    6.118706e-14, 6.103146e-14, 6.130695e-14, 6.114994e-14, 6.117449e-14, 
    6.102632e-14, 6.014367e-14, 6.030992e-14, 6.01338e-14, 6.015752e-14, 
    6.014689e-14, 6.001735e-14, 5.9952e-14, 5.981518e-14, 5.984005e-14, 
    5.994054e-14, 6.016819e-14, 6.009098e-14, 6.028558e-14, 6.028119e-14, 
    6.04975e-14, 6.040001e-14, 6.076313e-14, 6.066003e-14, 6.09578e-14, 
    6.088297e-14, 6.095427e-14, 6.093266e-14, 6.095456e-14, 6.08448e-14, 
    6.089183e-14, 6.079522e-14, 6.041826e-14, 6.052914e-14, 6.019818e-14, 
    5.999876e-14, 5.986627e-14, 5.977215e-14, 5.978546e-14, 5.981082e-14, 
    5.994113e-14, 6.006359e-14, 6.015683e-14, 6.021916e-14, 6.028056e-14, 
    6.046612e-14, 6.056434e-14, 6.078394e-14, 6.074438e-14, 6.081144e-14, 
    6.087552e-14, 6.0983e-14, 6.096532e-14, 6.101264e-14, 6.080969e-14, 
    6.094459e-14, 6.072183e-14, 6.078279e-14, 6.029708e-14, 6.011182e-14, 
    6.003287e-14, 5.996385e-14, 5.979569e-14, 5.991183e-14, 5.986605e-14, 
    5.997497e-14, 6.004412e-14, 6.000993e-14, 6.022086e-14, 6.013889e-14, 
    6.057016e-14, 6.038455e-14, 6.086805e-14, 6.07525e-14, 6.089573e-14, 
    6.082267e-14, 6.094782e-14, 6.083519e-14, 6.103026e-14, 6.107267e-14, 
    6.104369e-14, 6.115507e-14, 6.082895e-14, 6.095426e-14, 6.000896e-14, 
    6.001454e-14, 6.004053e-14, 5.992625e-14, 5.991926e-14, 5.98145e-14, 
    5.990773e-14, 5.994741e-14, 6.004814e-14, 6.010766e-14, 6.016423e-14, 
    6.028853e-14, 6.042721e-14, 6.062095e-14, 6.076e-14, 6.085312e-14, 
    6.079603e-14, 6.084644e-14, 6.079009e-14, 6.076368e-14, 6.105677e-14, 
    6.089226e-14, 6.113905e-14, 6.112541e-14, 6.101376e-14, 6.112695e-14, 
    6.001846e-14, 5.998637e-14, 5.987484e-14, 5.996213e-14, 5.980309e-14, 
    5.989211e-14, 5.994326e-14, 6.014057e-14, 6.018392e-14, 6.022406e-14, 
    6.030334e-14, 6.0405e-14, 6.058316e-14, 6.073802e-14, 6.087925e-14, 
    6.086891e-14, 6.087255e-14, 6.090407e-14, 6.082596e-14, 6.091689e-14, 
    6.093213e-14, 6.089226e-14, 6.112358e-14, 6.105754e-14, 6.112512e-14, 
    6.108213e-14, 5.99968e-14, 6.00508e-14, 6.002162e-14, 6.007648e-14, 
    6.003782e-14, 6.020959e-14, 6.026105e-14, 6.050164e-14, 6.040299e-14, 
    6.056001e-14, 6.041896e-14, 6.044395e-14, 6.056506e-14, 6.04266e-14, 
    6.072945e-14, 6.052413e-14, 6.090529e-14, 6.070045e-14, 6.091812e-14, 
    6.087864e-14, 6.094401e-14, 6.100251e-14, 6.10761e-14, 6.121174e-14, 
    6.118035e-14, 6.129373e-14, 6.013128e-14, 6.020123e-14, 6.019511e-14, 
    6.026831e-14, 6.032241e-14, 6.043965e-14, 6.062745e-14, 6.055687e-14, 
    6.068645e-14, 6.071244e-14, 6.051558e-14, 6.063645e-14, 6.024806e-14, 
    6.031085e-14, 6.027349e-14, 6.013678e-14, 6.057309e-14, 6.034932e-14, 
    6.076229e-14, 6.064127e-14, 6.099416e-14, 6.081875e-14, 6.116306e-14, 
    6.13099e-14, 6.144811e-14, 6.160927e-14, 6.023943e-14, 6.019191e-14, 
    6.027702e-14, 6.039463e-14, 6.050375e-14, 6.064865e-14, 6.066348e-14, 
    6.06906e-14, 6.076086e-14, 6.081989e-14, 6.069915e-14, 6.083469e-14, 
    6.032535e-14, 6.059252e-14, 6.017391e-14, 6.030005e-14, 6.038771e-14, 
    6.03493e-14, 6.05488e-14, 6.059577e-14, 6.078648e-14, 6.068795e-14, 
    6.127365e-14, 6.101482e-14, 6.173194e-14, 6.153191e-14, 6.017529e-14, 
    6.023928e-14, 6.046172e-14, 6.035593e-14, 6.065833e-14, 6.073266e-14, 
    6.079308e-14, 6.087023e-14, 6.087858e-14, 6.092426e-14, 6.084938e-14, 
    6.092132e-14, 6.064896e-14, 6.077074e-14, 6.043635e-14, 6.051779e-14, 
    6.048034e-14, 6.043922e-14, 6.056607e-14, 6.070104e-14, 6.070397e-14, 
    6.074721e-14, 6.086891e-14, 6.065956e-14, 6.130693e-14, 6.09074e-14, 
    6.030902e-14, 6.043207e-14, 6.044969e-14, 6.040203e-14, 6.072521e-14, 
    6.060819e-14, 6.092316e-14, 6.083811e-14, 6.097744e-14, 6.090822e-14, 
    6.089803e-14, 6.080908e-14, 6.075365e-14, 6.061355e-14, 6.049946e-14, 
    6.040895e-14, 6.043001e-14, 6.052941e-14, 6.07093e-14, 6.087931e-14, 
    6.084208e-14, 6.096686e-14, 6.063643e-14, 6.077505e-14, 6.072147e-14, 
    6.086115e-14, 6.055498e-14, 6.081559e-14, 6.048827e-14, 6.051701e-14, 
    6.060586e-14, 6.078442e-14, 6.082397e-14, 6.086609e-14, 6.084011e-14, 
    6.071388e-14, 6.069321e-14, 6.060372e-14, 6.057898e-14, 6.051076e-14, 
    6.045423e-14, 6.050587e-14, 6.056006e-14, 6.071395e-14, 6.085246e-14, 
    6.100333e-14, 6.104025e-14, 6.121616e-14, 6.107291e-14, 6.130914e-14, 
    6.110823e-14, 6.145589e-14, 6.083075e-14, 6.110242e-14, 6.060992e-14, 
    6.066308e-14, 6.075911e-14, 6.097923e-14, 6.086049e-14, 6.099937e-14, 
    6.06924e-14, 6.053282e-14, 6.049156e-14, 6.041445e-14, 6.049332e-14, 
    6.048691e-14, 6.056234e-14, 6.053811e-14, 6.071906e-14, 6.062189e-14, 
    6.089776e-14, 6.099828e-14, 6.128183e-14, 6.145533e-14, 6.163179e-14, 
    6.170959e-14, 6.173327e-14, 6.174316e-14 ;

 LITTERC =
  5.976256e-05, 5.976241e-05, 5.976244e-05, 5.976232e-05, 5.976239e-05, 
    5.976231e-05, 5.976253e-05, 5.976241e-05, 5.976249e-05, 5.976254e-05, 
    5.976209e-05, 5.976231e-05, 5.976186e-05, 5.9762e-05, 5.976164e-05, 
    5.976188e-05, 5.976159e-05, 5.976165e-05, 5.976148e-05, 5.976153e-05, 
    5.976132e-05, 5.976146e-05, 5.976121e-05, 5.976135e-05, 5.976133e-05, 
    5.976146e-05, 5.976227e-05, 5.976212e-05, 5.976228e-05, 5.976226e-05, 
    5.976227e-05, 5.976238e-05, 5.976245e-05, 5.976257e-05, 5.976255e-05, 
    5.976246e-05, 5.976225e-05, 5.976232e-05, 5.976214e-05, 5.976214e-05, 
    5.976195e-05, 5.976203e-05, 5.97617e-05, 5.97618e-05, 5.976153e-05, 
    5.976159e-05, 5.976153e-05, 5.976155e-05, 5.976153e-05, 5.976163e-05, 
    5.976159e-05, 5.976167e-05, 5.976202e-05, 5.976192e-05, 5.976222e-05, 
    5.97624e-05, 5.976252e-05, 5.976261e-05, 5.97626e-05, 5.976257e-05, 
    5.976246e-05, 5.976234e-05, 5.976226e-05, 5.97622e-05, 5.976214e-05, 
    5.976198e-05, 5.976189e-05, 5.976169e-05, 5.976172e-05, 5.976166e-05, 
    5.97616e-05, 5.97615e-05, 5.976152e-05, 5.976148e-05, 5.976166e-05, 
    5.976154e-05, 5.976174e-05, 5.976169e-05, 5.976213e-05, 5.97623e-05, 
    5.976237e-05, 5.976243e-05, 5.976259e-05, 5.976248e-05, 5.976252e-05, 
    5.976242e-05, 5.976236e-05, 5.976239e-05, 5.97622e-05, 5.976227e-05, 
    5.976188e-05, 5.976205e-05, 5.976161e-05, 5.976171e-05, 5.976158e-05, 
    5.976165e-05, 5.976154e-05, 5.976164e-05, 5.976146e-05, 5.976142e-05, 
    5.976145e-05, 5.976135e-05, 5.976165e-05, 5.976153e-05, 5.976239e-05, 
    5.976239e-05, 5.976237e-05, 5.976247e-05, 5.976247e-05, 5.976257e-05, 
    5.976249e-05, 5.976245e-05, 5.976236e-05, 5.97623e-05, 5.976225e-05, 
    5.976214e-05, 5.976201e-05, 5.976183e-05, 5.976171e-05, 5.976162e-05, 
    5.976167e-05, 5.976163e-05, 5.976168e-05, 5.97617e-05, 5.976144e-05, 
    5.976159e-05, 5.976136e-05, 5.976137e-05, 5.976147e-05, 5.976137e-05, 
    5.976238e-05, 5.976241e-05, 5.976251e-05, 5.976243e-05, 5.976258e-05, 
    5.97625e-05, 5.976245e-05, 5.976227e-05, 5.976223e-05, 5.97622e-05, 
    5.976213e-05, 5.976203e-05, 5.976187e-05, 5.976173e-05, 5.97616e-05, 
    5.976161e-05, 5.976161e-05, 5.976158e-05, 5.976165e-05, 5.976157e-05, 
    5.976155e-05, 5.976159e-05, 5.976138e-05, 5.976143e-05, 5.976137e-05, 
    5.976141e-05, 5.976241e-05, 5.976235e-05, 5.976238e-05, 5.976233e-05, 
    5.976237e-05, 5.976221e-05, 5.976216e-05, 5.976194e-05, 5.976203e-05, 
    5.976189e-05, 5.976202e-05, 5.976199e-05, 5.976189e-05, 5.976201e-05, 
    5.976174e-05, 5.976192e-05, 5.976158e-05, 5.976176e-05, 5.976156e-05, 
    5.97616e-05, 5.976154e-05, 5.976149e-05, 5.976142e-05, 5.97613e-05, 
    5.976133e-05, 5.976122e-05, 5.976228e-05, 5.976222e-05, 5.976222e-05, 
    5.976215e-05, 5.976211e-05, 5.9762e-05, 5.976183e-05, 5.976189e-05, 
    5.976178e-05, 5.976175e-05, 5.976193e-05, 5.976182e-05, 5.976218e-05, 
    5.976212e-05, 5.976215e-05, 5.976227e-05, 5.976188e-05, 5.976208e-05, 
    5.976171e-05, 5.976182e-05, 5.976149e-05, 5.976165e-05, 5.976134e-05, 
    5.976121e-05, 5.976108e-05, 5.976093e-05, 5.976218e-05, 5.976223e-05, 
    5.976215e-05, 5.976204e-05, 5.976194e-05, 5.976181e-05, 5.976179e-05, 
    5.976177e-05, 5.976171e-05, 5.976165e-05, 5.976176e-05, 5.976164e-05, 
    5.97621e-05, 5.976186e-05, 5.976224e-05, 5.976213e-05, 5.976205e-05, 
    5.976208e-05, 5.97619e-05, 5.976186e-05, 5.976168e-05, 5.976177e-05, 
    5.976124e-05, 5.976147e-05, 5.976082e-05, 5.9761e-05, 5.976224e-05, 
    5.976218e-05, 5.976198e-05, 5.976207e-05, 5.97618e-05, 5.976173e-05, 
    5.976168e-05, 5.976161e-05, 5.97616e-05, 5.976156e-05, 5.976163e-05, 
    5.976156e-05, 5.976181e-05, 5.97617e-05, 5.9762e-05, 5.976193e-05, 
    5.976196e-05, 5.9762e-05, 5.976189e-05, 5.976176e-05, 5.976176e-05, 
    5.976172e-05, 5.976161e-05, 5.97618e-05, 5.976121e-05, 5.976157e-05, 
    5.976212e-05, 5.976201e-05, 5.976199e-05, 5.976203e-05, 5.976174e-05, 
    5.976185e-05, 5.976156e-05, 5.976163e-05, 5.976151e-05, 5.976157e-05, 
    5.976158e-05, 5.976166e-05, 5.976171e-05, 5.976184e-05, 5.976194e-05, 
    5.976203e-05, 5.976201e-05, 5.976192e-05, 5.976175e-05, 5.97616e-05, 
    5.976163e-05, 5.976152e-05, 5.976182e-05, 5.976169e-05, 5.976174e-05, 
    5.976162e-05, 5.97619e-05, 5.976166e-05, 5.976195e-05, 5.976193e-05, 
    5.976185e-05, 5.976169e-05, 5.976165e-05, 5.976161e-05, 5.976163e-05, 
    5.976175e-05, 5.976177e-05, 5.976185e-05, 5.976187e-05, 5.976194e-05, 
    5.976199e-05, 5.976194e-05, 5.976189e-05, 5.976175e-05, 5.976162e-05, 
    5.976149e-05, 5.976145e-05, 5.976129e-05, 5.976142e-05, 5.976121e-05, 
    5.976139e-05, 5.976107e-05, 5.976164e-05, 5.976139e-05, 5.976185e-05, 
    5.976179e-05, 5.976171e-05, 5.976151e-05, 5.976162e-05, 5.976149e-05, 
    5.976177e-05, 5.976191e-05, 5.976195e-05, 5.976202e-05, 5.976195e-05, 
    5.976196e-05, 5.976189e-05, 5.976191e-05, 5.976174e-05, 5.976183e-05, 
    5.976158e-05, 5.976149e-05, 5.976123e-05, 5.976107e-05, 5.976091e-05, 
    5.976084e-05, 5.976082e-05, 5.976081e-05 ;

 LITTERC_HR =
  9.652399e-13, 9.678468e-13, 9.673404e-13, 9.69441e-13, 9.682762e-13, 
    9.696512e-13, 9.65769e-13, 9.679499e-13, 9.665581e-13, 9.654752e-13, 
    9.735113e-13, 9.695348e-13, 9.776379e-13, 9.751066e-13, 9.814612e-13, 
    9.772438e-13, 9.823108e-13, 9.813404e-13, 9.842616e-13, 9.834251e-13, 
    9.871558e-13, 9.846476e-13, 9.890884e-13, 9.865574e-13, 9.869532e-13, 
    9.845646e-13, 9.703362e-13, 9.730164e-13, 9.701772e-13, 9.705597e-13, 
    9.703883e-13, 9.683001e-13, 9.672466e-13, 9.650411e-13, 9.654418e-13, 
    9.670618e-13, 9.707316e-13, 9.69487e-13, 9.726239e-13, 9.725531e-13, 
    9.760401e-13, 9.744686e-13, 9.803222e-13, 9.786601e-13, 9.834602e-13, 
    9.822538e-13, 9.834034e-13, 9.830549e-13, 9.834079e-13, 9.816385e-13, 
    9.823967e-13, 9.808393e-13, 9.747628e-13, 9.765501e-13, 9.712151e-13, 
    9.680003e-13, 9.658645e-13, 9.643473e-13, 9.645619e-13, 9.649706e-13, 
    9.670714e-13, 9.690454e-13, 9.705484e-13, 9.715532e-13, 9.725429e-13, 
    9.755342e-13, 9.771176e-13, 9.806576e-13, 9.800199e-13, 9.811007e-13, 
    9.821338e-13, 9.838663e-13, 9.835813e-13, 9.843441e-13, 9.810728e-13, 
    9.832472e-13, 9.796564e-13, 9.80639e-13, 9.728094e-13, 9.69823e-13, 
    9.685502e-13, 9.674376e-13, 9.647268e-13, 9.66599e-13, 9.658611e-13, 
    9.676169e-13, 9.687315e-13, 9.681804e-13, 9.715807e-13, 9.702592e-13, 
    9.772114e-13, 9.742194e-13, 9.820133e-13, 9.801509e-13, 9.824597e-13, 
    9.812819e-13, 9.832993e-13, 9.814838e-13, 9.846282e-13, 9.85312e-13, 
    9.848446e-13, 9.866401e-13, 9.813831e-13, 9.83403e-13, 9.681649e-13, 
    9.682548e-13, 9.686737e-13, 9.668314e-13, 9.667188e-13, 9.650299e-13, 
    9.66533e-13, 9.671725e-13, 9.687963e-13, 9.697559e-13, 9.706678e-13, 
    9.726715e-13, 9.74907e-13, 9.7803e-13, 9.802715e-13, 9.817727e-13, 
    9.808526e-13, 9.816649e-13, 9.807566e-13, 9.803309e-13, 9.850556e-13, 
    9.824036e-13, 9.86382e-13, 9.861621e-13, 9.843621e-13, 9.861868e-13, 
    9.683179e-13, 9.678006e-13, 9.660028e-13, 9.674099e-13, 9.64846e-13, 
    9.662811e-13, 9.671057e-13, 9.702864e-13, 9.709851e-13, 9.716322e-13, 
    9.729102e-13, 9.74549e-13, 9.774209e-13, 9.799172e-13, 9.82194e-13, 
    9.820273e-13, 9.820859e-13, 9.82594e-13, 9.813349e-13, 9.828006e-13, 
    9.830463e-13, 9.824036e-13, 9.861326e-13, 9.850679e-13, 9.861574e-13, 
    9.854643e-13, 9.679688e-13, 9.688393e-13, 9.683689e-13, 9.692532e-13, 
    9.6863e-13, 9.71399e-13, 9.722285e-13, 9.761069e-13, 9.745166e-13, 
    9.770478e-13, 9.747741e-13, 9.75177e-13, 9.771292e-13, 9.748971e-13, 
    9.797791e-13, 9.764694e-13, 9.826137e-13, 9.793118e-13, 9.828205e-13, 
    9.821842e-13, 9.832379e-13, 9.841808e-13, 9.853672e-13, 9.875536e-13, 
    9.870476e-13, 9.888752e-13, 9.701366e-13, 9.712643e-13, 9.711655e-13, 
    9.723455e-13, 9.732176e-13, 9.751076e-13, 9.781349e-13, 9.769971e-13, 
    9.790861e-13, 9.79505e-13, 9.763315e-13, 9.782801e-13, 9.720191e-13, 
    9.730312e-13, 9.724291e-13, 9.702253e-13, 9.772586e-13, 9.736515e-13, 
    9.803085e-13, 9.783578e-13, 9.840464e-13, 9.812186e-13, 9.867688e-13, 
    9.891361e-13, 9.913638e-13, 9.939616e-13, 9.7188e-13, 9.71114e-13, 
    9.724859e-13, 9.743818e-13, 9.761409e-13, 9.784767e-13, 9.787158e-13, 
    9.79153e-13, 9.802855e-13, 9.81237e-13, 9.792907e-13, 9.814755e-13, 
    9.73265e-13, 9.775718e-13, 9.708239e-13, 9.728572e-13, 9.742703e-13, 
    9.73651e-13, 9.768671e-13, 9.776243e-13, 9.806985e-13, 9.791101e-13, 
    9.885516e-13, 9.843794e-13, 9.959391e-13, 9.927146e-13, 9.708461e-13, 
    9.718776e-13, 9.754633e-13, 9.73758e-13, 9.786328e-13, 9.798309e-13, 
    9.808048e-13, 9.820484e-13, 9.821831e-13, 9.829196e-13, 9.817124e-13, 
    9.828721e-13, 9.784816e-13, 9.804448e-13, 9.750543e-13, 9.763672e-13, 
    9.757635e-13, 9.751008e-13, 9.771456e-13, 9.793212e-13, 9.793685e-13, 
    9.800655e-13, 9.820272e-13, 9.786526e-13, 9.89088e-13, 9.826478e-13, 
    9.730018e-13, 9.749854e-13, 9.752695e-13, 9.745013e-13, 9.797108e-13, 
    9.778245e-13, 9.829017e-13, 9.815308e-13, 9.837768e-13, 9.826609e-13, 
    9.824966e-13, 9.810628e-13, 9.801694e-13, 9.779108e-13, 9.760718e-13, 
    9.746128e-13, 9.749522e-13, 9.765546e-13, 9.794544e-13, 9.821949e-13, 
    9.815947e-13, 9.836062e-13, 9.782796e-13, 9.805143e-13, 9.796506e-13, 
    9.819021e-13, 9.769667e-13, 9.811677e-13, 9.758914e-13, 9.763546e-13, 
    9.77787e-13, 9.806652e-13, 9.813027e-13, 9.819817e-13, 9.815629e-13, 
    9.795281e-13, 9.791949e-13, 9.777524e-13, 9.773535e-13, 9.762538e-13, 
    9.753425e-13, 9.76175e-13, 9.770486e-13, 9.795293e-13, 9.817621e-13, 
    9.841942e-13, 9.847893e-13, 9.876248e-13, 9.853158e-13, 9.891237e-13, 
    9.85885e-13, 9.914891e-13, 9.814121e-13, 9.857913e-13, 9.778525e-13, 
    9.787092e-13, 9.802573e-13, 9.838056e-13, 9.818915e-13, 9.841302e-13, 
    9.791819e-13, 9.766094e-13, 9.759444e-13, 9.747013e-13, 9.759728e-13, 
    9.758695e-13, 9.770854e-13, 9.766947e-13, 9.796117e-13, 9.780453e-13, 
    9.824923e-13, 9.841127e-13, 9.886835e-13, 9.914802e-13, 9.943246e-13, 
    9.955787e-13, 9.959604e-13, 9.961199e-13 ;

 LITTERC_LOSS =
  1.787615e-12, 1.792443e-12, 1.791505e-12, 1.795395e-12, 1.793238e-12, 
    1.795785e-12, 1.788595e-12, 1.792634e-12, 1.790056e-12, 1.788051e-12, 
    1.802934e-12, 1.795569e-12, 1.810576e-12, 1.805888e-12, 1.817657e-12, 
    1.809846e-12, 1.819231e-12, 1.817433e-12, 1.822843e-12, 1.821294e-12, 
    1.828203e-12, 1.823558e-12, 1.831783e-12, 1.827095e-12, 1.827828e-12, 
    1.823405e-12, 1.797053e-12, 1.802017e-12, 1.796759e-12, 1.797467e-12, 
    1.79715e-12, 1.793282e-12, 1.791331e-12, 1.787247e-12, 1.787989e-12, 
    1.790989e-12, 1.797786e-12, 1.795481e-12, 1.80129e-12, 1.801159e-12, 
    1.807617e-12, 1.804706e-12, 1.815547e-12, 1.812469e-12, 1.821359e-12, 
    1.819125e-12, 1.821254e-12, 1.820609e-12, 1.821262e-12, 1.817985e-12, 
    1.819389e-12, 1.816505e-12, 1.805251e-12, 1.808562e-12, 1.798681e-12, 
    1.792727e-12, 1.788772e-12, 1.785962e-12, 1.786359e-12, 1.787116e-12, 
    1.791007e-12, 1.794663e-12, 1.797446e-12, 1.799307e-12, 1.80114e-12, 
    1.80668e-12, 1.809613e-12, 1.816169e-12, 1.814988e-12, 1.816989e-12, 
    1.818903e-12, 1.822111e-12, 1.821583e-12, 1.822996e-12, 1.816937e-12, 
    1.820965e-12, 1.814314e-12, 1.816134e-12, 1.801634e-12, 1.796103e-12, 
    1.793746e-12, 1.791685e-12, 1.786664e-12, 1.790132e-12, 1.788765e-12, 
    1.792017e-12, 1.794081e-12, 1.793061e-12, 1.799358e-12, 1.796911e-12, 
    1.809786e-12, 1.804245e-12, 1.81868e-12, 1.81523e-12, 1.819506e-12, 
    1.817325e-12, 1.821061e-12, 1.817699e-12, 1.823522e-12, 1.824789e-12, 
    1.823923e-12, 1.827248e-12, 1.817512e-12, 1.821253e-12, 1.793032e-12, 
    1.793198e-12, 1.793974e-12, 1.790562e-12, 1.790354e-12, 1.787226e-12, 
    1.79001e-12, 1.791194e-12, 1.794201e-12, 1.795978e-12, 1.797667e-12, 
    1.801378e-12, 1.805519e-12, 1.811303e-12, 1.815454e-12, 1.818234e-12, 
    1.81653e-12, 1.818034e-12, 1.816352e-12, 1.815564e-12, 1.824314e-12, 
    1.819402e-12, 1.82677e-12, 1.826363e-12, 1.82303e-12, 1.826409e-12, 
    1.793315e-12, 1.792357e-12, 1.789028e-12, 1.791634e-12, 1.786885e-12, 
    1.789543e-12, 1.79107e-12, 1.796961e-12, 1.798255e-12, 1.799453e-12, 
    1.80182e-12, 1.804855e-12, 1.810174e-12, 1.814797e-12, 1.819014e-12, 
    1.818705e-12, 1.818814e-12, 1.819755e-12, 1.817423e-12, 1.820138e-12, 
    1.820593e-12, 1.819402e-12, 1.826309e-12, 1.824337e-12, 1.826354e-12, 
    1.825071e-12, 1.792669e-12, 1.794281e-12, 1.79341e-12, 1.795048e-12, 
    1.793893e-12, 1.799021e-12, 1.800558e-12, 1.807741e-12, 1.804795e-12, 
    1.809483e-12, 1.805272e-12, 1.806018e-12, 1.809634e-12, 1.8055e-12, 
    1.814542e-12, 1.808412e-12, 1.819791e-12, 1.813676e-12, 1.820174e-12, 
    1.818996e-12, 1.820947e-12, 1.822694e-12, 1.824891e-12, 1.82894e-12, 
    1.828003e-12, 1.831388e-12, 1.796684e-12, 1.798772e-12, 1.798589e-12, 
    1.800774e-12, 1.80239e-12, 1.80589e-12, 1.811497e-12, 1.809389e-12, 
    1.813258e-12, 1.814034e-12, 1.808157e-12, 1.811765e-12, 1.80017e-12, 
    1.802045e-12, 1.800929e-12, 1.796848e-12, 1.809874e-12, 1.803193e-12, 
    1.815522e-12, 1.811909e-12, 1.822445e-12, 1.817208e-12, 1.827487e-12, 
    1.831871e-12, 1.835997e-12, 1.840808e-12, 1.799913e-12, 1.798494e-12, 
    1.801035e-12, 1.804546e-12, 1.807804e-12, 1.81213e-12, 1.812572e-12, 
    1.813382e-12, 1.81548e-12, 1.817242e-12, 1.813637e-12, 1.817683e-12, 
    1.802477e-12, 1.810454e-12, 1.797956e-12, 1.801722e-12, 1.804339e-12, 
    1.803192e-12, 1.809149e-12, 1.810551e-12, 1.816245e-12, 1.813303e-12, 
    1.830789e-12, 1.823061e-12, 1.844471e-12, 1.838499e-12, 1.797998e-12, 
    1.799908e-12, 1.806549e-12, 1.803391e-12, 1.812419e-12, 1.814638e-12, 
    1.816441e-12, 1.818745e-12, 1.818994e-12, 1.820358e-12, 1.818122e-12, 
    1.82027e-12, 1.812139e-12, 1.815775e-12, 1.805791e-12, 1.808223e-12, 
    1.807105e-12, 1.805877e-12, 1.809664e-12, 1.813694e-12, 1.813781e-12, 
    1.815072e-12, 1.818705e-12, 1.812455e-12, 1.831782e-12, 1.819855e-12, 
    1.80199e-12, 1.805664e-12, 1.80619e-12, 1.804767e-12, 1.814415e-12, 
    1.810922e-12, 1.820325e-12, 1.817786e-12, 1.821945e-12, 1.819879e-12, 
    1.819575e-12, 1.816919e-12, 1.815265e-12, 1.811082e-12, 1.807676e-12, 
    1.804974e-12, 1.805602e-12, 1.80857e-12, 1.81394e-12, 1.819016e-12, 
    1.817904e-12, 1.821629e-12, 1.811765e-12, 1.815903e-12, 1.814304e-12, 
    1.818474e-12, 1.809333e-12, 1.817114e-12, 1.807341e-12, 1.8082e-12, 
    1.810852e-12, 1.816183e-12, 1.817363e-12, 1.818621e-12, 1.817845e-12, 
    1.814077e-12, 1.81346e-12, 1.810788e-12, 1.81005e-12, 1.808013e-12, 
    1.806325e-12, 1.807867e-12, 1.809485e-12, 1.814079e-12, 1.818214e-12, 
    1.822719e-12, 1.823821e-12, 1.829072e-12, 1.824796e-12, 1.831848e-12, 
    1.82585e-12, 1.836229e-12, 1.817566e-12, 1.825676e-12, 1.810973e-12, 
    1.81256e-12, 1.815427e-12, 1.821999e-12, 1.818454e-12, 1.8226e-12, 
    1.813436e-12, 1.808671e-12, 1.80744e-12, 1.805138e-12, 1.807492e-12, 
    1.807301e-12, 1.809553e-12, 1.808829e-12, 1.814232e-12, 1.811331e-12, 
    1.819567e-12, 1.822568e-12, 1.831033e-12, 1.836212e-12, 1.84148e-12, 
    1.843803e-12, 1.84451e-12, 1.844805e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  1.676328e-18, 1.676591e-18, 1.676541e-18, 1.676751e-18, 1.676636e-18, 
    1.676772e-18, 1.676384e-18, 1.676599e-18, 1.676463e-18, 1.676355e-18, 
    1.677151e-18, 1.676761e-18, 1.67758e-18, 1.677327e-18, 1.677971e-18, 
    1.677538e-18, 1.67806e-18, 1.677964e-18, 1.678265e-18, 1.678179e-18, 
    1.678554e-18, 1.678305e-18, 1.678757e-18, 1.678497e-18, 1.678536e-18, 
    1.678296e-18, 1.676844e-18, 1.677101e-18, 1.676828e-18, 1.676865e-18, 
    1.676849e-18, 1.676637e-18, 1.676527e-18, 1.676311e-18, 1.676351e-18, 
    1.676511e-18, 1.676881e-18, 1.676759e-18, 1.677077e-18, 1.67707e-18, 
    1.677422e-18, 1.677263e-18, 1.677859e-18, 1.677691e-18, 1.678183e-18, 
    1.678058e-18, 1.678176e-18, 1.678141e-18, 1.678176e-18, 1.677994e-18, 
    1.678072e-18, 1.677913e-18, 1.677292e-18, 1.677473e-18, 1.676932e-18, 
    1.6766e-18, 1.676392e-18, 1.676241e-18, 1.676262e-18, 1.676302e-18, 
    1.676512e-18, 1.676714e-18, 1.676867e-18, 1.676968e-18, 1.677069e-18, 
    1.677361e-18, 1.677527e-18, 1.677891e-18, 1.67783e-18, 1.677937e-18, 
    1.678046e-18, 1.678223e-18, 1.678194e-18, 1.678271e-18, 1.677937e-18, 
    1.678158e-18, 1.677794e-18, 1.677893e-18, 1.677079e-18, 1.676793e-18, 
    1.676656e-18, 1.67655e-18, 1.676279e-18, 1.676465e-18, 1.676391e-18, 
    1.676571e-18, 1.676682e-18, 1.676628e-18, 1.676971e-18, 1.676837e-18, 
    1.677537e-18, 1.677235e-18, 1.678033e-18, 1.677843e-18, 1.678079e-18, 
    1.677959e-18, 1.678164e-18, 1.67798e-18, 1.678301e-18, 1.67837e-18, 
    1.678323e-18, 1.678509e-18, 1.677969e-18, 1.678174e-18, 1.676626e-18, 
    1.676634e-18, 1.676677e-18, 1.676488e-18, 1.676478e-18, 1.676309e-18, 
    1.676461e-18, 1.676524e-18, 1.67669e-18, 1.676786e-18, 1.676878e-18, 
    1.677081e-18, 1.677304e-18, 1.677623e-18, 1.677855e-18, 1.67801e-18, 
    1.677916e-18, 1.677998e-18, 1.677905e-18, 1.677862e-18, 1.678343e-18, 
    1.678071e-18, 1.678482e-18, 1.67846e-18, 1.678273e-18, 1.678462e-18, 
    1.676641e-18, 1.67659e-18, 1.676407e-18, 1.67655e-18, 1.676291e-18, 
    1.676434e-18, 1.676515e-18, 1.676836e-18, 1.676911e-18, 1.676975e-18, 
    1.677106e-18, 1.677271e-18, 1.677561e-18, 1.677817e-18, 1.678053e-18, 
    1.678036e-18, 1.678042e-18, 1.678093e-18, 1.677964e-18, 1.678114e-18, 
    1.678137e-18, 1.678073e-18, 1.678457e-18, 1.678347e-18, 1.678459e-18, 
    1.678389e-18, 1.676607e-18, 1.676694e-18, 1.676646e-18, 1.676734e-18, 
    1.676671e-18, 1.676948e-18, 1.677031e-18, 1.677424e-18, 1.677267e-18, 
    1.677522e-18, 1.677294e-18, 1.677334e-18, 1.677523e-18, 1.677308e-18, 
    1.677799e-18, 1.677459e-18, 1.678095e-18, 1.677748e-18, 1.678116e-18, 
    1.678052e-18, 1.67816e-18, 1.678255e-18, 1.678378e-18, 1.6786e-18, 
    1.678549e-18, 1.678738e-18, 1.676825e-18, 1.676936e-18, 1.67693e-18, 
    1.677048e-18, 1.677136e-18, 1.677329e-18, 1.677636e-18, 1.677521e-18, 
    1.677735e-18, 1.677777e-18, 1.677454e-18, 1.677649e-18, 1.677013e-18, 
    1.677112e-18, 1.677056e-18, 1.676832e-18, 1.677543e-18, 1.677176e-18, 
    1.677858e-18, 1.677659e-18, 1.678241e-18, 1.677948e-18, 1.67852e-18, 
    1.678757e-18, 1.678996e-18, 1.679258e-18, 1.677e-18, 1.676924e-18, 
    1.677064e-18, 1.67725e-18, 1.677433e-18, 1.677671e-18, 1.677697e-18, 
    1.67774e-18, 1.677858e-18, 1.677954e-18, 1.677751e-18, 1.677979e-18, 
    1.677129e-18, 1.677576e-18, 1.676893e-18, 1.677094e-18, 1.677241e-18, 
    1.67718e-18, 1.677509e-18, 1.677586e-18, 1.677896e-18, 1.677737e-18, 
    1.678696e-18, 1.67827e-18, 1.679468e-18, 1.67913e-18, 1.676897e-18, 
    1.677002e-18, 1.677362e-18, 1.677191e-18, 1.677688e-18, 1.677809e-18, 
    1.677911e-18, 1.678035e-18, 1.678051e-18, 1.678125e-18, 1.678003e-18, 
    1.678122e-18, 1.677671e-18, 1.677873e-18, 1.677324e-18, 1.677456e-18, 
    1.677396e-18, 1.677329e-18, 1.677537e-18, 1.677753e-18, 1.677763e-18, 
    1.677832e-18, 1.678016e-18, 1.67769e-18, 1.678741e-18, 1.678082e-18, 
    1.677116e-18, 1.67731e-18, 1.677344e-18, 1.677268e-18, 1.677797e-18, 
    1.677604e-18, 1.678124e-18, 1.677985e-18, 1.678215e-18, 1.6781e-18, 
    1.678083e-18, 1.677937e-18, 1.677844e-18, 1.677612e-18, 1.677425e-18, 
    1.67728e-18, 1.677314e-18, 1.677474e-18, 1.677768e-18, 1.67805e-18, 
    1.677988e-18, 1.678197e-18, 1.677652e-18, 1.677878e-18, 1.677789e-18, 
    1.678022e-18, 1.677517e-18, 1.677931e-18, 1.677409e-18, 1.677456e-18, 
    1.677601e-18, 1.677889e-18, 1.677961e-18, 1.678029e-18, 1.677988e-18, 
    1.677776e-18, 1.677744e-18, 1.677598e-18, 1.677556e-18, 1.677446e-18, 
    1.677354e-18, 1.677437e-18, 1.677524e-18, 1.677779e-18, 1.678006e-18, 
    1.678256e-18, 1.678319e-18, 1.678598e-18, 1.678364e-18, 1.678744e-18, 
    1.678409e-18, 1.678994e-18, 1.677963e-18, 1.67841e-18, 1.677609e-18, 
    1.677696e-18, 1.677849e-18, 1.678211e-18, 1.678021e-18, 1.678246e-18, 
    1.677743e-18, 1.677477e-18, 1.677414e-18, 1.677287e-18, 1.677417e-18, 
    1.677407e-18, 1.677531e-18, 1.677492e-18, 1.677787e-18, 1.677628e-18, 
    1.678081e-18, 1.678245e-18, 1.678716e-18, 1.679002e-18, 1.679303e-18, 
    1.679433e-18, 1.679473e-18, 1.679489e-18 ;

 MEG_acetic_acid =
  2.514492e-19, 2.514887e-19, 2.514812e-19, 2.515126e-19, 2.514954e-19, 
    2.515158e-19, 2.514575e-19, 2.514899e-19, 2.514694e-19, 2.514532e-19, 
    2.515727e-19, 2.515141e-19, 2.51637e-19, 2.51599e-19, 2.516957e-19, 
    2.516306e-19, 2.517089e-19, 2.516945e-19, 2.517397e-19, 2.517268e-19, 
    2.517831e-19, 2.517457e-19, 2.518136e-19, 2.517746e-19, 2.517804e-19, 
    2.517443e-19, 2.515266e-19, 2.515652e-19, 2.515241e-19, 2.515297e-19, 
    2.515274e-19, 2.514955e-19, 2.51479e-19, 2.514467e-19, 2.514527e-19, 
    2.514767e-19, 2.515322e-19, 2.515139e-19, 2.515616e-19, 2.515605e-19, 
    2.516133e-19, 2.515895e-19, 2.516789e-19, 2.516536e-19, 2.517274e-19, 
    2.517087e-19, 2.517264e-19, 2.517211e-19, 2.517264e-19, 2.516991e-19, 
    2.517108e-19, 2.516869e-19, 2.515938e-19, 2.516209e-19, 2.515398e-19, 
    2.514899e-19, 2.514588e-19, 2.514362e-19, 2.514394e-19, 2.514453e-19, 
    2.514768e-19, 2.515072e-19, 2.515301e-19, 2.515453e-19, 2.515604e-19, 
    2.516042e-19, 2.516291e-19, 2.516836e-19, 2.516744e-19, 2.516905e-19, 
    2.517069e-19, 2.517334e-19, 2.517292e-19, 2.517407e-19, 2.516906e-19, 
    2.517236e-19, 2.51669e-19, 2.516839e-19, 2.515619e-19, 2.515189e-19, 
    2.514984e-19, 2.514825e-19, 2.514418e-19, 2.514698e-19, 2.514586e-19, 
    2.514856e-19, 2.515024e-19, 2.514942e-19, 2.515457e-19, 2.515256e-19, 
    2.516305e-19, 2.515853e-19, 2.51705e-19, 2.516764e-19, 2.517119e-19, 
    2.516939e-19, 2.517246e-19, 2.51697e-19, 2.517452e-19, 2.517554e-19, 
    2.517484e-19, 2.517763e-19, 2.516954e-19, 2.517261e-19, 2.514938e-19, 
    2.514951e-19, 2.515016e-19, 2.514732e-19, 2.514716e-19, 2.514464e-19, 
    2.514691e-19, 2.514785e-19, 2.515035e-19, 2.515179e-19, 2.515317e-19, 
    2.515621e-19, 2.515956e-19, 2.516434e-19, 2.516782e-19, 2.517014e-19, 
    2.516874e-19, 2.516998e-19, 2.516858e-19, 2.516794e-19, 2.517514e-19, 
    2.517107e-19, 2.517723e-19, 2.51769e-19, 2.517409e-19, 2.517694e-19, 
    2.514961e-19, 2.514884e-19, 2.51461e-19, 2.514825e-19, 2.514437e-19, 
    2.514651e-19, 2.514772e-19, 2.515254e-19, 2.515366e-19, 2.515462e-19, 
    2.515658e-19, 2.515907e-19, 2.516342e-19, 2.516725e-19, 2.517079e-19, 
    2.517054e-19, 2.517063e-19, 2.517139e-19, 2.516946e-19, 2.517171e-19, 
    2.517206e-19, 2.51711e-19, 2.517685e-19, 2.517521e-19, 2.517689e-19, 
    2.517583e-19, 2.51491e-19, 2.51504e-19, 2.514969e-19, 2.515101e-19, 
    2.515006e-19, 2.515421e-19, 2.515546e-19, 2.516137e-19, 2.515901e-19, 
    2.516284e-19, 2.515941e-19, 2.516001e-19, 2.516285e-19, 2.515962e-19, 
    2.516699e-19, 2.516189e-19, 2.517142e-19, 2.516621e-19, 2.517174e-19, 
    2.517078e-19, 2.51724e-19, 2.517383e-19, 2.517567e-19, 2.5179e-19, 
    2.517824e-19, 2.518107e-19, 2.515237e-19, 2.515404e-19, 2.515394e-19, 
    2.515573e-19, 2.515703e-19, 2.515993e-19, 2.516453e-19, 2.516282e-19, 
    2.516602e-19, 2.516665e-19, 2.516181e-19, 2.516473e-19, 2.51552e-19, 
    2.515668e-19, 2.515583e-19, 2.515248e-19, 2.516314e-19, 2.515763e-19, 
    2.516787e-19, 2.516488e-19, 2.517361e-19, 2.516922e-19, 2.517781e-19, 
    2.518136e-19, 2.518494e-19, 2.518886e-19, 2.515501e-19, 2.515387e-19, 
    2.515595e-19, 2.515875e-19, 2.516149e-19, 2.516506e-19, 2.516545e-19, 
    2.51661e-19, 2.516786e-19, 2.516932e-19, 2.516626e-19, 2.516969e-19, 
    2.515693e-19, 2.516365e-19, 2.515339e-19, 2.515641e-19, 2.515861e-19, 
    2.515769e-19, 2.516263e-19, 2.516378e-19, 2.516844e-19, 2.516606e-19, 
    2.518044e-19, 2.517406e-19, 2.519202e-19, 2.518695e-19, 2.515346e-19, 
    2.515503e-19, 2.516042e-19, 2.515786e-19, 2.516532e-19, 2.516714e-19, 
    2.516866e-19, 2.517053e-19, 2.517077e-19, 2.517188e-19, 2.517005e-19, 
    2.517183e-19, 2.516507e-19, 2.516809e-19, 2.515986e-19, 2.516183e-19, 
    2.516094e-19, 2.515993e-19, 2.516305e-19, 2.51663e-19, 2.516645e-19, 
    2.516748e-19, 2.517024e-19, 2.516535e-19, 2.518112e-19, 2.517123e-19, 
    2.515673e-19, 2.515965e-19, 2.516017e-19, 2.515902e-19, 2.516695e-19, 
    2.516406e-19, 2.517186e-19, 2.516977e-19, 2.517322e-19, 2.51715e-19, 
    2.517124e-19, 2.516905e-19, 2.516767e-19, 2.516418e-19, 2.516138e-19, 
    2.515919e-19, 2.515971e-19, 2.516211e-19, 2.516652e-19, 2.517075e-19, 
    2.516981e-19, 2.517296e-19, 2.516478e-19, 2.516816e-19, 2.516683e-19, 
    2.517033e-19, 2.516275e-19, 2.516896e-19, 2.516114e-19, 2.516184e-19, 
    2.516401e-19, 2.516834e-19, 2.516942e-19, 2.517043e-19, 2.516982e-19, 
    2.516664e-19, 2.516616e-19, 2.516397e-19, 2.516333e-19, 2.51617e-19, 
    2.51603e-19, 2.516156e-19, 2.516285e-19, 2.516668e-19, 2.517008e-19, 
    2.517383e-19, 2.517478e-19, 2.517897e-19, 2.517545e-19, 2.518116e-19, 
    2.517614e-19, 2.518491e-19, 2.516944e-19, 2.517615e-19, 2.516413e-19, 
    2.516545e-19, 2.516773e-19, 2.517316e-19, 2.517031e-19, 2.517368e-19, 
    2.516615e-19, 2.516215e-19, 2.516122e-19, 2.515931e-19, 2.516126e-19, 
    2.51611e-19, 2.516297e-19, 2.516237e-19, 2.51668e-19, 2.516443e-19, 
    2.517121e-19, 2.517368e-19, 2.518074e-19, 2.518503e-19, 2.518954e-19, 
    2.519149e-19, 2.519209e-19, 2.519234e-19 ;

 MEG_acetone =
  8.435572e-17, 8.436433e-17, 8.436269e-17, 8.436956e-17, 8.436581e-17, 
    8.437026e-17, 8.435754e-17, 8.436461e-17, 8.436014e-17, 8.43566e-17, 
    8.438267e-17, 8.436988e-17, 8.43967e-17, 8.43884e-17, 8.44095e-17, 
    8.439531e-17, 8.44124e-17, 8.440926e-17, 8.441913e-17, 8.441631e-17, 
    8.442859e-17, 8.442043e-17, 8.443525e-17, 8.442673e-17, 8.4428e-17, 
    8.442013e-17, 8.437261e-17, 8.438103e-17, 8.437208e-17, 8.437328e-17, 
    8.437278e-17, 8.436583e-17, 8.436222e-17, 8.435518e-17, 8.435649e-17, 
    8.436172e-17, 8.437383e-17, 8.436983e-17, 8.438025e-17, 8.438002e-17, 
    8.439153e-17, 8.438633e-17, 8.440585e-17, 8.440033e-17, 8.441643e-17, 
    8.441235e-17, 8.441621e-17, 8.441506e-17, 8.441622e-17, 8.441025e-17, 
    8.44128e-17, 8.440761e-17, 8.438727e-17, 8.439319e-17, 8.437548e-17, 
    8.436461e-17, 8.435782e-17, 8.435288e-17, 8.435358e-17, 8.435487e-17, 
    8.436175e-17, 8.436837e-17, 8.437337e-17, 8.437668e-17, 8.437999e-17, 
    8.438954e-17, 8.439497e-17, 8.440688e-17, 8.440487e-17, 8.440839e-17, 
    8.441196e-17, 8.441775e-17, 8.441682e-17, 8.441934e-17, 8.44084e-17, 
    8.441561e-17, 8.44037e-17, 8.440693e-17, 8.43803e-17, 8.437093e-17, 
    8.436647e-17, 8.436299e-17, 8.43541e-17, 8.436021e-17, 8.435778e-17, 
    8.436367e-17, 8.436733e-17, 8.436554e-17, 8.437678e-17, 8.437238e-17, 
    8.439529e-17, 8.438542e-17, 8.441154e-17, 8.44053e-17, 8.441305e-17, 
    8.440912e-17, 8.441581e-17, 8.440979e-17, 8.442033e-17, 8.442256e-17, 
    8.442101e-17, 8.442712e-17, 8.440945e-17, 8.441616e-17, 8.436546e-17, 
    8.436575e-17, 8.436715e-17, 8.436096e-17, 8.436062e-17, 8.435512e-17, 
    8.436006e-17, 8.436212e-17, 8.436759e-17, 8.437071e-17, 8.437372e-17, 
    8.438035e-17, 8.438768e-17, 8.43981e-17, 8.440569e-17, 8.441076e-17, 
    8.440769e-17, 8.44104e-17, 8.440736e-17, 8.440595e-17, 8.442168e-17, 
    8.441279e-17, 8.442624e-17, 8.442551e-17, 8.441937e-17, 8.442559e-17, 
    8.436596e-17, 8.436429e-17, 8.435829e-17, 8.436299e-17, 8.435452e-17, 
    8.435919e-17, 8.436183e-17, 8.437235e-17, 8.43748e-17, 8.43769e-17, 
    8.438118e-17, 8.43866e-17, 8.439609e-17, 8.440445e-17, 8.441219e-17, 
    8.441163e-17, 8.441182e-17, 8.441349e-17, 8.440928e-17, 8.441419e-17, 
    8.441495e-17, 8.441286e-17, 8.442541e-17, 8.442183e-17, 8.442549e-17, 
    8.442318e-17, 8.436485e-17, 8.436769e-17, 8.436614e-17, 8.436902e-17, 
    8.436695e-17, 8.4376e-17, 8.437872e-17, 8.439161e-17, 8.438646e-17, 
    8.439482e-17, 8.438735e-17, 8.438864e-17, 8.439485e-17, 8.438779e-17, 
    8.440388e-17, 8.439275e-17, 8.441356e-17, 8.440219e-17, 8.441425e-17, 
    8.441215e-17, 8.441569e-17, 8.44188e-17, 8.442283e-17, 8.443009e-17, 
    8.442843e-17, 8.443461e-17, 8.437199e-17, 8.437563e-17, 8.437541e-17, 
    8.43793e-17, 8.438216e-17, 8.438848e-17, 8.439852e-17, 8.439478e-17, 
    8.440177e-17, 8.440313e-17, 8.439258e-17, 8.439895e-17, 8.437815e-17, 
    8.438139e-17, 8.437954e-17, 8.437221e-17, 8.439549e-17, 8.438346e-17, 
    8.44058e-17, 8.439929e-17, 8.441835e-17, 8.440875e-17, 8.442749e-17, 
    8.443525e-17, 8.444307e-17, 8.445164e-17, 8.437773e-17, 8.437524e-17, 
    8.437979e-17, 8.43859e-17, 8.439188e-17, 8.439967e-17, 8.440053e-17, 
    8.440195e-17, 8.440579e-17, 8.440896e-17, 8.44023e-17, 8.440977e-17, 
    8.438193e-17, 8.439658e-17, 8.43742e-17, 8.438079e-17, 8.438558e-17, 
    8.438359e-17, 8.439438e-17, 8.439688e-17, 8.440704e-17, 8.440185e-17, 
    8.443324e-17, 8.441931e-17, 8.445854e-17, 8.444746e-17, 8.437435e-17, 
    8.437778e-17, 8.438956e-17, 8.438396e-17, 8.440024e-17, 8.440421e-17, 
    8.440753e-17, 8.441161e-17, 8.441213e-17, 8.441456e-17, 8.441057e-17, 
    8.441444e-17, 8.439968e-17, 8.440629e-17, 8.438834e-17, 8.439263e-17, 
    8.439069e-17, 8.438848e-17, 8.439529e-17, 8.440238e-17, 8.44027e-17, 
    8.440495e-17, 8.441097e-17, 8.440032e-17, 8.443472e-17, 8.441313e-17, 
    8.43815e-17, 8.438787e-17, 8.438899e-17, 8.438648e-17, 8.440381e-17, 
    8.43975e-17, 8.441452e-17, 8.440996e-17, 8.441749e-17, 8.441373e-17, 
    8.441317e-17, 8.440838e-17, 8.440536e-17, 8.439775e-17, 8.439163e-17, 
    8.438687e-17, 8.438799e-17, 8.439323e-17, 8.440285e-17, 8.44121e-17, 
    8.441005e-17, 8.441692e-17, 8.439906e-17, 8.440644e-17, 8.440353e-17, 
    8.441117e-17, 8.439464e-17, 8.440818e-17, 8.439112e-17, 8.439265e-17, 
    8.439738e-17, 8.440683e-17, 8.440918e-17, 8.441139e-17, 8.441006e-17, 
    8.440313e-17, 8.440207e-17, 8.43973e-17, 8.43959e-17, 8.439233e-17, 
    8.438929e-17, 8.439202e-17, 8.439486e-17, 8.44032e-17, 8.441064e-17, 
    8.441882e-17, 8.44209e-17, 8.443004e-17, 8.442235e-17, 8.443481e-17, 
    8.442385e-17, 8.444301e-17, 8.440923e-17, 8.442389e-17, 8.439765e-17, 
    8.440051e-17, 8.44055e-17, 8.441735e-17, 8.441113e-17, 8.441849e-17, 
    8.440204e-17, 8.439332e-17, 8.439128e-17, 8.438713e-17, 8.439138e-17, 
    8.439104e-17, 8.43951e-17, 8.43938e-17, 8.440348e-17, 8.439829e-17, 
    8.441311e-17, 8.441848e-17, 8.44339e-17, 8.444328e-17, 8.445312e-17, 
    8.445738e-17, 8.445869e-17, 8.445923e-17 ;

 MEG_carene_3 =
  3.259777e-17, 3.260117e-17, 3.260052e-17, 3.260323e-17, 3.260176e-17, 
    3.260351e-17, 3.259848e-17, 3.260128e-17, 3.259951e-17, 3.259811e-17, 
    3.260842e-17, 3.260336e-17, 3.261397e-17, 3.261069e-17, 3.261903e-17, 
    3.261342e-17, 3.262017e-17, 3.261893e-17, 3.262283e-17, 3.262172e-17, 
    3.262657e-17, 3.262334e-17, 3.26292e-17, 3.262584e-17, 3.262634e-17, 
    3.262323e-17, 3.260444e-17, 3.260777e-17, 3.260423e-17, 3.260471e-17, 
    3.260451e-17, 3.260176e-17, 3.260033e-17, 3.259755e-17, 3.259807e-17, 
    3.260014e-17, 3.260493e-17, 3.260334e-17, 3.260746e-17, 3.260737e-17, 
    3.261192e-17, 3.260987e-17, 3.261758e-17, 3.26154e-17, 3.262177e-17, 
    3.262015e-17, 3.262168e-17, 3.262122e-17, 3.262168e-17, 3.261932e-17, 
    3.262033e-17, 3.261828e-17, 3.261024e-17, 3.261258e-17, 3.260558e-17, 
    3.260128e-17, 3.25986e-17, 3.259664e-17, 3.259691e-17, 3.259743e-17, 
    3.260015e-17, 3.260276e-17, 3.260474e-17, 3.260605e-17, 3.260736e-17, 
    3.261113e-17, 3.261328e-17, 3.261799e-17, 3.26172e-17, 3.261858e-17, 
    3.262e-17, 3.262229e-17, 3.262192e-17, 3.262291e-17, 3.261859e-17, 
    3.262144e-17, 3.261673e-17, 3.261801e-17, 3.260748e-17, 3.260378e-17, 
    3.260201e-17, 3.260064e-17, 3.259712e-17, 3.259954e-17, 3.259858e-17, 
    3.260091e-17, 3.260235e-17, 3.260165e-17, 3.260609e-17, 3.260435e-17, 
    3.261341e-17, 3.26095e-17, 3.261983e-17, 3.261736e-17, 3.262043e-17, 
    3.261887e-17, 3.262152e-17, 3.261914e-17, 3.262331e-17, 3.262419e-17, 
    3.262358e-17, 3.262599e-17, 3.2619e-17, 3.262166e-17, 3.260162e-17, 
    3.260173e-17, 3.260228e-17, 3.259984e-17, 3.25997e-17, 3.259752e-17, 
    3.259948e-17, 3.26003e-17, 3.260245e-17, 3.260369e-17, 3.260488e-17, 
    3.26075e-17, 3.26104e-17, 3.261452e-17, 3.261752e-17, 3.261953e-17, 
    3.261831e-17, 3.261938e-17, 3.261818e-17, 3.261762e-17, 3.262384e-17, 
    3.262033e-17, 3.262564e-17, 3.262536e-17, 3.262293e-17, 3.262539e-17, 
    3.260181e-17, 3.260115e-17, 3.259878e-17, 3.260064e-17, 3.259729e-17, 
    3.259914e-17, 3.260018e-17, 3.260434e-17, 3.260531e-17, 3.260614e-17, 
    3.260783e-17, 3.260997e-17, 3.261372e-17, 3.261703e-17, 3.262009e-17, 
    3.261987e-17, 3.261994e-17, 3.26206e-17, 3.261894e-17, 3.262088e-17, 
    3.262118e-17, 3.262035e-17, 3.262532e-17, 3.26239e-17, 3.262535e-17, 
    3.262443e-17, 3.260137e-17, 3.26025e-17, 3.260188e-17, 3.260302e-17, 
    3.26022e-17, 3.260578e-17, 3.260685e-17, 3.261195e-17, 3.260991e-17, 
    3.261322e-17, 3.261027e-17, 3.261078e-17, 3.261323e-17, 3.261044e-17, 
    3.26168e-17, 3.26124e-17, 3.262063e-17, 3.261614e-17, 3.26209e-17, 
    3.262007e-17, 3.262147e-17, 3.26227e-17, 3.262429e-17, 3.262717e-17, 
    3.262651e-17, 3.262895e-17, 3.260419e-17, 3.260563e-17, 3.260555e-17, 
    3.260709e-17, 3.260821e-17, 3.261072e-17, 3.261468e-17, 3.26132e-17, 
    3.261597e-17, 3.261651e-17, 3.261234e-17, 3.261485e-17, 3.260663e-17, 
    3.260791e-17, 3.260718e-17, 3.260428e-17, 3.261349e-17, 3.260873e-17, 
    3.261756e-17, 3.261499e-17, 3.262252e-17, 3.261873e-17, 3.262614e-17, 
    3.26292e-17, 3.26323e-17, 3.263568e-17, 3.260647e-17, 3.260548e-17, 
    3.260728e-17, 3.26097e-17, 3.261206e-17, 3.261514e-17, 3.261548e-17, 
    3.261604e-17, 3.261756e-17, 3.261881e-17, 3.261618e-17, 3.261913e-17, 
    3.260812e-17, 3.261392e-17, 3.260507e-17, 3.260767e-17, 3.260957e-17, 
    3.260878e-17, 3.261305e-17, 3.261404e-17, 3.261805e-17, 3.2616e-17, 
    3.262841e-17, 3.26229e-17, 3.263841e-17, 3.263403e-17, 3.260513e-17, 
    3.260648e-17, 3.261114e-17, 3.260893e-17, 3.261537e-17, 3.261694e-17, 
    3.261825e-17, 3.261986e-17, 3.262007e-17, 3.262103e-17, 3.261945e-17, 
    3.262098e-17, 3.261514e-17, 3.261776e-17, 3.261066e-17, 3.261236e-17, 
    3.261159e-17, 3.261072e-17, 3.261341e-17, 3.261621e-17, 3.261634e-17, 
    3.261722e-17, 3.261961e-17, 3.261539e-17, 3.262899e-17, 3.262046e-17, 
    3.260796e-17, 3.261047e-17, 3.261092e-17, 3.260993e-17, 3.261677e-17, 
    3.261428e-17, 3.262101e-17, 3.261921e-17, 3.262218e-17, 3.26207e-17, 
    3.262048e-17, 3.261858e-17, 3.261739e-17, 3.261438e-17, 3.261196e-17, 
    3.261008e-17, 3.261052e-17, 3.261259e-17, 3.26164e-17, 3.262005e-17, 
    3.261924e-17, 3.262196e-17, 3.26149e-17, 3.261782e-17, 3.261666e-17, 
    3.261969e-17, 3.261315e-17, 3.26185e-17, 3.261176e-17, 3.261236e-17, 
    3.261423e-17, 3.261797e-17, 3.26189e-17, 3.261977e-17, 3.261925e-17, 
    3.261651e-17, 3.261609e-17, 3.26142e-17, 3.261365e-17, 3.261224e-17, 
    3.261104e-17, 3.261212e-17, 3.261324e-17, 3.261654e-17, 3.261947e-17, 
    3.262271e-17, 3.262353e-17, 3.262715e-17, 3.262411e-17, 3.262903e-17, 
    3.26247e-17, 3.263227e-17, 3.261892e-17, 3.262471e-17, 3.261434e-17, 
    3.261547e-17, 3.261745e-17, 3.262213e-17, 3.261967e-17, 3.262258e-17, 
    3.261608e-17, 3.261263e-17, 3.261182e-17, 3.261018e-17, 3.261186e-17, 
    3.261173e-17, 3.261333e-17, 3.261282e-17, 3.261665e-17, 3.261459e-17, 
    3.262045e-17, 3.262257e-17, 3.262867e-17, 3.263237e-17, 3.263627e-17, 
    3.263795e-17, 3.263847e-17, 3.263868e-17 ;

 MEG_ethanol =
  1.676328e-18, 1.676591e-18, 1.676541e-18, 1.676751e-18, 1.676636e-18, 
    1.676772e-18, 1.676384e-18, 1.676599e-18, 1.676463e-18, 1.676355e-18, 
    1.677151e-18, 1.676761e-18, 1.67758e-18, 1.677327e-18, 1.677971e-18, 
    1.677538e-18, 1.67806e-18, 1.677964e-18, 1.678265e-18, 1.678179e-18, 
    1.678554e-18, 1.678305e-18, 1.678757e-18, 1.678497e-18, 1.678536e-18, 
    1.678296e-18, 1.676844e-18, 1.677101e-18, 1.676828e-18, 1.676865e-18, 
    1.676849e-18, 1.676637e-18, 1.676527e-18, 1.676311e-18, 1.676351e-18, 
    1.676511e-18, 1.676881e-18, 1.676759e-18, 1.677077e-18, 1.67707e-18, 
    1.677422e-18, 1.677263e-18, 1.677859e-18, 1.677691e-18, 1.678183e-18, 
    1.678058e-18, 1.678176e-18, 1.678141e-18, 1.678176e-18, 1.677994e-18, 
    1.678072e-18, 1.677913e-18, 1.677292e-18, 1.677473e-18, 1.676932e-18, 
    1.6766e-18, 1.676392e-18, 1.676241e-18, 1.676262e-18, 1.676302e-18, 
    1.676512e-18, 1.676714e-18, 1.676867e-18, 1.676968e-18, 1.677069e-18, 
    1.677361e-18, 1.677527e-18, 1.677891e-18, 1.67783e-18, 1.677937e-18, 
    1.678046e-18, 1.678223e-18, 1.678194e-18, 1.678271e-18, 1.677937e-18, 
    1.678158e-18, 1.677794e-18, 1.677893e-18, 1.677079e-18, 1.676793e-18, 
    1.676656e-18, 1.67655e-18, 1.676279e-18, 1.676465e-18, 1.676391e-18, 
    1.676571e-18, 1.676682e-18, 1.676628e-18, 1.676971e-18, 1.676837e-18, 
    1.677537e-18, 1.677235e-18, 1.678033e-18, 1.677843e-18, 1.678079e-18, 
    1.677959e-18, 1.678164e-18, 1.67798e-18, 1.678301e-18, 1.67837e-18, 
    1.678323e-18, 1.678509e-18, 1.677969e-18, 1.678174e-18, 1.676626e-18, 
    1.676634e-18, 1.676677e-18, 1.676488e-18, 1.676478e-18, 1.676309e-18, 
    1.676461e-18, 1.676524e-18, 1.67669e-18, 1.676786e-18, 1.676878e-18, 
    1.677081e-18, 1.677304e-18, 1.677623e-18, 1.677855e-18, 1.67801e-18, 
    1.677916e-18, 1.677998e-18, 1.677905e-18, 1.677862e-18, 1.678343e-18, 
    1.678071e-18, 1.678482e-18, 1.67846e-18, 1.678273e-18, 1.678462e-18, 
    1.676641e-18, 1.67659e-18, 1.676407e-18, 1.67655e-18, 1.676291e-18, 
    1.676434e-18, 1.676515e-18, 1.676836e-18, 1.676911e-18, 1.676975e-18, 
    1.677106e-18, 1.677271e-18, 1.677561e-18, 1.677817e-18, 1.678053e-18, 
    1.678036e-18, 1.678042e-18, 1.678093e-18, 1.677964e-18, 1.678114e-18, 
    1.678137e-18, 1.678073e-18, 1.678457e-18, 1.678347e-18, 1.678459e-18, 
    1.678389e-18, 1.676607e-18, 1.676694e-18, 1.676646e-18, 1.676734e-18, 
    1.676671e-18, 1.676948e-18, 1.677031e-18, 1.677424e-18, 1.677267e-18, 
    1.677522e-18, 1.677294e-18, 1.677334e-18, 1.677523e-18, 1.677308e-18, 
    1.677799e-18, 1.677459e-18, 1.678095e-18, 1.677748e-18, 1.678116e-18, 
    1.678052e-18, 1.67816e-18, 1.678255e-18, 1.678378e-18, 1.6786e-18, 
    1.678549e-18, 1.678738e-18, 1.676825e-18, 1.676936e-18, 1.67693e-18, 
    1.677048e-18, 1.677136e-18, 1.677329e-18, 1.677636e-18, 1.677521e-18, 
    1.677735e-18, 1.677777e-18, 1.677454e-18, 1.677649e-18, 1.677013e-18, 
    1.677112e-18, 1.677056e-18, 1.676832e-18, 1.677543e-18, 1.677176e-18, 
    1.677858e-18, 1.677659e-18, 1.678241e-18, 1.677948e-18, 1.67852e-18, 
    1.678757e-18, 1.678996e-18, 1.679258e-18, 1.677e-18, 1.676924e-18, 
    1.677064e-18, 1.67725e-18, 1.677433e-18, 1.677671e-18, 1.677697e-18, 
    1.67774e-18, 1.677858e-18, 1.677954e-18, 1.677751e-18, 1.677979e-18, 
    1.677129e-18, 1.677576e-18, 1.676893e-18, 1.677094e-18, 1.677241e-18, 
    1.67718e-18, 1.677509e-18, 1.677586e-18, 1.677896e-18, 1.677737e-18, 
    1.678696e-18, 1.67827e-18, 1.679468e-18, 1.67913e-18, 1.676897e-18, 
    1.677002e-18, 1.677362e-18, 1.677191e-18, 1.677688e-18, 1.677809e-18, 
    1.677911e-18, 1.678035e-18, 1.678051e-18, 1.678125e-18, 1.678003e-18, 
    1.678122e-18, 1.677671e-18, 1.677873e-18, 1.677324e-18, 1.677456e-18, 
    1.677396e-18, 1.677329e-18, 1.677537e-18, 1.677753e-18, 1.677763e-18, 
    1.677832e-18, 1.678016e-18, 1.67769e-18, 1.678741e-18, 1.678082e-18, 
    1.677116e-18, 1.67731e-18, 1.677344e-18, 1.677268e-18, 1.677797e-18, 
    1.677604e-18, 1.678124e-18, 1.677985e-18, 1.678215e-18, 1.6781e-18, 
    1.678083e-18, 1.677937e-18, 1.677844e-18, 1.677612e-18, 1.677425e-18, 
    1.67728e-18, 1.677314e-18, 1.677474e-18, 1.677768e-18, 1.67805e-18, 
    1.677988e-18, 1.678197e-18, 1.677652e-18, 1.677878e-18, 1.677789e-18, 
    1.678022e-18, 1.677517e-18, 1.677931e-18, 1.677409e-18, 1.677456e-18, 
    1.677601e-18, 1.677889e-18, 1.677961e-18, 1.678029e-18, 1.677988e-18, 
    1.677776e-18, 1.677744e-18, 1.677598e-18, 1.677556e-18, 1.677446e-18, 
    1.677354e-18, 1.677437e-18, 1.677524e-18, 1.677779e-18, 1.678006e-18, 
    1.678256e-18, 1.678319e-18, 1.678598e-18, 1.678364e-18, 1.678744e-18, 
    1.678409e-18, 1.678994e-18, 1.677963e-18, 1.67841e-18, 1.677609e-18, 
    1.677696e-18, 1.677849e-18, 1.678211e-18, 1.678021e-18, 1.678246e-18, 
    1.677743e-18, 1.677477e-18, 1.677414e-18, 1.677287e-18, 1.677417e-18, 
    1.677407e-18, 1.677531e-18, 1.677492e-18, 1.677787e-18, 1.677628e-18, 
    1.678081e-18, 1.678245e-18, 1.678716e-18, 1.679002e-18, 1.679303e-18, 
    1.679433e-18, 1.679473e-18, 1.679489e-18 ;

 MEG_formaldehyde =
  3.352656e-19, 3.353182e-19, 3.353082e-19, 3.353501e-19, 3.353273e-19, 
    3.353544e-19, 3.352767e-19, 3.353199e-19, 3.352926e-19, 3.352709e-19, 
    3.354303e-19, 3.353521e-19, 3.35516e-19, 3.354653e-19, 3.355942e-19, 
    3.355075e-19, 3.356119e-19, 3.355927e-19, 3.35653e-19, 3.356358e-19, 
    3.357108e-19, 3.356609e-19, 3.357514e-19, 3.356994e-19, 3.357071e-19, 
    3.356591e-19, 3.353688e-19, 3.354202e-19, 3.353655e-19, 3.353729e-19, 
    3.353698e-19, 3.353274e-19, 3.353053e-19, 3.352623e-19, 3.352703e-19, 
    3.353023e-19, 3.353763e-19, 3.353518e-19, 3.354155e-19, 3.354141e-19, 
    3.354844e-19, 3.354527e-19, 3.355718e-19, 3.355382e-19, 3.356365e-19, 
    3.356116e-19, 3.356352e-19, 3.356281e-19, 3.356353e-19, 3.355988e-19, 
    3.356143e-19, 3.355826e-19, 3.354584e-19, 3.354945e-19, 3.353864e-19, 
    3.353199e-19, 3.352784e-19, 3.352482e-19, 3.352525e-19, 3.352604e-19, 
    3.353024e-19, 3.353429e-19, 3.353734e-19, 3.353937e-19, 3.354138e-19, 
    3.354722e-19, 3.355054e-19, 3.355782e-19, 3.355659e-19, 3.355874e-19, 
    3.356091e-19, 3.356446e-19, 3.356388e-19, 3.356543e-19, 3.355874e-19, 
    3.356315e-19, 3.355587e-19, 3.355785e-19, 3.354158e-19, 3.353586e-19, 
    3.353312e-19, 3.3531e-19, 3.352557e-19, 3.35293e-19, 3.352782e-19, 
    3.353142e-19, 3.353365e-19, 3.353256e-19, 3.353943e-19, 3.353674e-19, 
    3.355074e-19, 3.35447e-19, 3.356066e-19, 3.355685e-19, 3.356159e-19, 
    3.355919e-19, 3.356327e-19, 3.35596e-19, 3.356603e-19, 3.356739e-19, 
    3.356645e-19, 3.357018e-19, 3.355938e-19, 3.356348e-19, 3.353251e-19, 
    3.353269e-19, 3.353355e-19, 3.352976e-19, 3.352955e-19, 3.352619e-19, 
    3.352921e-19, 3.353047e-19, 3.353381e-19, 3.353572e-19, 3.353756e-19, 
    3.354161e-19, 3.354608e-19, 3.355245e-19, 3.355709e-19, 3.356019e-19, 
    3.355831e-19, 3.355997e-19, 3.35581e-19, 3.355725e-19, 3.356686e-19, 
    3.356143e-19, 3.356964e-19, 3.35692e-19, 3.356545e-19, 3.356925e-19, 
    3.353282e-19, 3.353179e-19, 3.352813e-19, 3.3531e-19, 3.352583e-19, 
    3.352868e-19, 3.353029e-19, 3.353672e-19, 3.353822e-19, 3.35395e-19, 
    3.354211e-19, 3.354543e-19, 3.355122e-19, 3.355633e-19, 3.356106e-19, 
    3.356072e-19, 3.356083e-19, 3.356185e-19, 3.355928e-19, 3.356228e-19, 
    3.356275e-19, 3.356147e-19, 3.356913e-19, 3.356695e-19, 3.356919e-19, 
    3.356777e-19, 3.353213e-19, 3.353387e-19, 3.353293e-19, 3.353469e-19, 
    3.353342e-19, 3.353895e-19, 3.354061e-19, 3.354849e-19, 3.354534e-19, 
    3.355045e-19, 3.354589e-19, 3.354667e-19, 3.355047e-19, 3.354615e-19, 
    3.355599e-19, 3.354918e-19, 3.356189e-19, 3.355495e-19, 3.356232e-19, 
    3.356104e-19, 3.35632e-19, 3.35651e-19, 3.356756e-19, 3.3572e-19, 
    3.357098e-19, 3.357475e-19, 3.35365e-19, 3.353872e-19, 3.353859e-19, 
    3.354097e-19, 3.354271e-19, 3.354658e-19, 3.355271e-19, 3.355042e-19, 
    3.355469e-19, 3.355553e-19, 3.354908e-19, 3.355297e-19, 3.354026e-19, 
    3.354224e-19, 3.354111e-19, 3.353663e-19, 3.355086e-19, 3.354351e-19, 
    3.355716e-19, 3.355318e-19, 3.356482e-19, 3.355896e-19, 3.357041e-19, 
    3.357515e-19, 3.357992e-19, 3.358515e-19, 3.354001e-19, 3.353849e-19, 
    3.354127e-19, 3.3545e-19, 3.354865e-19, 3.355341e-19, 3.355393e-19, 
    3.355481e-19, 3.355715e-19, 3.355909e-19, 3.355502e-19, 3.355958e-19, 
    3.354257e-19, 3.355153e-19, 3.353785e-19, 3.354188e-19, 3.354481e-19, 
    3.354359e-19, 3.355018e-19, 3.355171e-19, 3.355792e-19, 3.355474e-19, 
    3.357392e-19, 3.356541e-19, 3.358936e-19, 3.35826e-19, 3.353794e-19, 
    3.354003e-19, 3.354723e-19, 3.354382e-19, 3.355376e-19, 3.355619e-19, 
    3.355822e-19, 3.356071e-19, 3.356102e-19, 3.356251e-19, 3.356007e-19, 
    3.356244e-19, 3.355342e-19, 3.355746e-19, 3.354649e-19, 3.354911e-19, 
    3.354793e-19, 3.354658e-19, 3.355074e-19, 3.355506e-19, 3.355526e-19, 
    3.355664e-19, 3.356031e-19, 3.355381e-19, 3.357482e-19, 3.356164e-19, 
    3.354231e-19, 3.35462e-19, 3.354689e-19, 3.354536e-19, 3.355594e-19, 
    3.355209e-19, 3.356249e-19, 3.355969e-19, 3.35643e-19, 3.3562e-19, 
    3.356166e-19, 3.355873e-19, 3.355689e-19, 3.355224e-19, 3.35485e-19, 
    3.354559e-19, 3.354628e-19, 3.354948e-19, 3.355535e-19, 3.3561e-19, 
    3.355975e-19, 3.356395e-19, 3.355304e-19, 3.355755e-19, 3.355577e-19, 
    3.356044e-19, 3.355034e-19, 3.355861e-19, 3.354819e-19, 3.354912e-19, 
    3.355201e-19, 3.355779e-19, 3.355922e-19, 3.356057e-19, 3.355976e-19, 
    3.355553e-19, 3.355488e-19, 3.355197e-19, 3.355111e-19, 3.354893e-19, 
    3.354707e-19, 3.354874e-19, 3.355047e-19, 3.355557e-19, 3.356011e-19, 
    3.356511e-19, 3.356638e-19, 3.357197e-19, 3.356727e-19, 3.357488e-19, 
    3.356819e-19, 3.357989e-19, 3.355925e-19, 3.35682e-19, 3.355218e-19, 
    3.355393e-19, 3.355698e-19, 3.356421e-19, 3.356042e-19, 3.356491e-19, 
    3.355486e-19, 3.354953e-19, 3.354829e-19, 3.354575e-19, 3.354835e-19, 
    3.354814e-19, 3.355062e-19, 3.354983e-19, 3.355574e-19, 3.355257e-19, 
    3.356162e-19, 3.35649e-19, 3.357432e-19, 3.358004e-19, 3.358605e-19, 
    3.358866e-19, 3.358946e-19, 3.358979e-19 ;

 MEG_isoprene =
  2.294623e-19, 2.295062e-19, 2.294979e-19, 2.295328e-19, 2.295137e-19, 
    2.295364e-19, 2.294716e-19, 2.295076e-19, 2.294848e-19, 2.294668e-19, 
    2.295996e-19, 2.295345e-19, 2.29671e-19, 2.296288e-19, 2.297361e-19, 
    2.296639e-19, 2.297509e-19, 2.297349e-19, 2.297851e-19, 2.297707e-19, 
    2.298332e-19, 2.297917e-19, 2.29867e-19, 2.298237e-19, 2.298302e-19, 
    2.297902e-19, 2.295484e-19, 2.295912e-19, 2.295456e-19, 2.295518e-19, 
    2.295492e-19, 2.295138e-19, 2.294954e-19, 2.294596e-19, 2.294662e-19, 
    2.294929e-19, 2.295546e-19, 2.295342e-19, 2.295872e-19, 2.295861e-19, 
    2.296447e-19, 2.296182e-19, 2.297175e-19, 2.296894e-19, 2.297713e-19, 
    2.297506e-19, 2.297702e-19, 2.297644e-19, 2.297703e-19, 2.297399e-19, 
    2.297529e-19, 2.297265e-19, 2.29623e-19, 2.296531e-19, 2.29563e-19, 
    2.295076e-19, 2.29473e-19, 2.294479e-19, 2.294514e-19, 2.29458e-19, 
    2.294931e-19, 2.295267e-19, 2.295522e-19, 2.295691e-19, 2.295859e-19, 
    2.296345e-19, 2.296622e-19, 2.297228e-19, 2.297126e-19, 2.297304e-19, 
    2.297486e-19, 2.297781e-19, 2.297733e-19, 2.297861e-19, 2.297305e-19, 
    2.297672e-19, 2.297066e-19, 2.29723e-19, 2.295875e-19, 2.295398e-19, 
    2.295171e-19, 2.294993e-19, 2.294541e-19, 2.294852e-19, 2.294729e-19, 
    2.295028e-19, 2.295214e-19, 2.295124e-19, 2.295696e-19, 2.295472e-19, 
    2.296638e-19, 2.296136e-19, 2.297465e-19, 2.297147e-19, 2.297542e-19, 
    2.297342e-19, 2.297682e-19, 2.297376e-19, 2.297911e-19, 2.298025e-19, 
    2.297947e-19, 2.298257e-19, 2.297358e-19, 2.297699e-19, 2.29512e-19, 
    2.295134e-19, 2.295206e-19, 2.29489e-19, 2.294873e-19, 2.294593e-19, 
    2.294844e-19, 2.294949e-19, 2.295227e-19, 2.295387e-19, 2.29554e-19, 
    2.295878e-19, 2.296251e-19, 2.296781e-19, 2.297167e-19, 2.297425e-19, 
    2.297269e-19, 2.297407e-19, 2.297252e-19, 2.29718e-19, 2.29798e-19, 
    2.297528e-19, 2.298212e-19, 2.298175e-19, 2.297863e-19, 2.298179e-19, 
    2.295145e-19, 2.29506e-19, 2.294755e-19, 2.294993e-19, 2.294562e-19, 
    2.2948e-19, 2.294935e-19, 2.29547e-19, 2.295595e-19, 2.295702e-19, 
    2.295919e-19, 2.296195e-19, 2.296679e-19, 2.297104e-19, 2.297498e-19, 
    2.297469e-19, 2.297479e-19, 2.297564e-19, 2.297349e-19, 2.297599e-19, 
    2.297638e-19, 2.297532e-19, 2.29817e-19, 2.297988e-19, 2.298175e-19, 
    2.298056e-19, 2.295088e-19, 2.295233e-19, 2.295154e-19, 2.295301e-19, 
    2.295195e-19, 2.295656e-19, 2.295795e-19, 2.296451e-19, 2.296188e-19, 
    2.296614e-19, 2.296234e-19, 2.2963e-19, 2.296616e-19, 2.296256e-19, 
    2.297075e-19, 2.296509e-19, 2.297567e-19, 2.296989e-19, 2.297603e-19, 
    2.297496e-19, 2.297676e-19, 2.297834e-19, 2.298039e-19, 2.298408e-19, 
    2.298324e-19, 2.298638e-19, 2.295452e-19, 2.295637e-19, 2.295626e-19, 
    2.295824e-19, 2.29597e-19, 2.296291e-19, 2.296802e-19, 2.296612e-19, 
    2.296968e-19, 2.297037e-19, 2.2965e-19, 2.296824e-19, 2.295765e-19, 
    2.295931e-19, 2.295836e-19, 2.295463e-19, 2.296648e-19, 2.296036e-19, 
    2.297173e-19, 2.296841e-19, 2.297811e-19, 2.297323e-19, 2.298276e-19, 
    2.298671e-19, 2.299068e-19, 2.299503e-19, 2.295744e-19, 2.295617e-19, 
    2.295849e-19, 2.29616e-19, 2.296464e-19, 2.296861e-19, 2.296904e-19, 
    2.296977e-19, 2.297172e-19, 2.297334e-19, 2.296995e-19, 2.297375e-19, 
    2.295958e-19, 2.296704e-19, 2.295565e-19, 2.2959e-19, 2.296144e-19, 
    2.296042e-19, 2.296591e-19, 2.296719e-19, 2.297236e-19, 2.296972e-19, 
    2.298568e-19, 2.29786e-19, 2.299853e-19, 2.299291e-19, 2.295572e-19, 
    2.295746e-19, 2.296346e-19, 2.296061e-19, 2.29689e-19, 2.297092e-19, 
    2.297261e-19, 2.297468e-19, 2.297495e-19, 2.297618e-19, 2.297415e-19, 
    2.297612e-19, 2.296861e-19, 2.297198e-19, 2.296284e-19, 2.296503e-19, 
    2.296404e-19, 2.296292e-19, 2.296638e-19, 2.296999e-19, 2.297015e-19, 
    2.297129e-19, 2.297436e-19, 2.296894e-19, 2.298644e-19, 2.297546e-19, 
    2.295936e-19, 2.29626e-19, 2.296317e-19, 2.29619e-19, 2.297071e-19, 
    2.29675e-19, 2.297616e-19, 2.297384e-19, 2.297767e-19, 2.297576e-19, 
    2.297547e-19, 2.297304e-19, 2.29715e-19, 2.296764e-19, 2.296452e-19, 
    2.296209e-19, 2.296266e-19, 2.296533e-19, 2.297023e-19, 2.297493e-19, 
    2.297389e-19, 2.297738e-19, 2.29683e-19, 2.297206e-19, 2.297057e-19, 
    2.297446e-19, 2.296605e-19, 2.297294e-19, 2.296426e-19, 2.296504e-19, 
    2.296744e-19, 2.297225e-19, 2.297345e-19, 2.297457e-19, 2.297389e-19, 
    2.297037e-19, 2.296983e-19, 2.29674e-19, 2.296669e-19, 2.296487e-19, 
    2.296333e-19, 2.296472e-19, 2.296616e-19, 2.29704e-19, 2.297419e-19, 
    2.297835e-19, 2.29794e-19, 2.298406e-19, 2.298015e-19, 2.298648e-19, 
    2.298091e-19, 2.299065e-19, 2.297347e-19, 2.298093e-19, 2.296758e-19, 
    2.296904e-19, 2.297158e-19, 2.29776e-19, 2.297444e-19, 2.297818e-19, 
    2.296982e-19, 2.296538e-19, 2.296434e-19, 2.296223e-19, 2.296439e-19, 
    2.296422e-19, 2.296628e-19, 2.296563e-19, 2.297055e-19, 2.296791e-19, 
    2.297544e-19, 2.297818e-19, 2.298602e-19, 2.299078e-19, 2.299578e-19, 
    2.299794e-19, 2.299861e-19, 2.299889e-19 ;

 MEG_methanol =
  5.798236e-17, 5.798805e-17, 5.798697e-17, 5.79915e-17, 5.798903e-17, 
    5.799197e-17, 5.798356e-17, 5.798823e-17, 5.798527e-17, 5.798294e-17, 
    5.800016e-17, 5.799171e-17, 5.800943e-17, 5.800395e-17, 5.801787e-17, 
    5.800851e-17, 5.801978e-17, 5.801771e-17, 5.802422e-17, 5.802236e-17, 
    5.803046e-17, 5.802508e-17, 5.803485e-17, 5.802923e-17, 5.803007e-17, 
    5.802488e-17, 5.799352e-17, 5.799907e-17, 5.799316e-17, 5.799396e-17, 
    5.799363e-17, 5.798904e-17, 5.798665e-17, 5.7982e-17, 5.798287e-17, 
    5.798633e-17, 5.799432e-17, 5.799168e-17, 5.799856e-17, 5.799841e-17, 
    5.800601e-17, 5.800258e-17, 5.801546e-17, 5.801182e-17, 5.802244e-17, 
    5.801975e-17, 5.802229e-17, 5.802154e-17, 5.802231e-17, 5.801837e-17, 
    5.802005e-17, 5.801662e-17, 5.80032e-17, 5.800711e-17, 5.799541e-17, 
    5.798823e-17, 5.798375e-17, 5.798048e-17, 5.798094e-17, 5.79818e-17, 
    5.798634e-17, 5.799071e-17, 5.799402e-17, 5.799621e-17, 5.799838e-17, 
    5.80047e-17, 5.800828e-17, 5.801614e-17, 5.801482e-17, 5.801713e-17, 
    5.801949e-17, 5.802331e-17, 5.80227e-17, 5.802436e-17, 5.801714e-17, 
    5.80219e-17, 5.801404e-17, 5.801618e-17, 5.79986e-17, 5.799241e-17, 
    5.798946e-17, 5.798716e-17, 5.798129e-17, 5.798532e-17, 5.798373e-17, 
    5.798761e-17, 5.799003e-17, 5.798885e-17, 5.799627e-17, 5.799337e-17, 
    5.80085e-17, 5.800198e-17, 5.801922e-17, 5.801509e-17, 5.802022e-17, 
    5.801762e-17, 5.802203e-17, 5.801806e-17, 5.802501e-17, 5.802648e-17, 
    5.802546e-17, 5.802949e-17, 5.801783e-17, 5.802226e-17, 5.79888e-17, 
    5.798899e-17, 5.798991e-17, 5.798582e-17, 5.798559e-17, 5.798196e-17, 
    5.798523e-17, 5.798659e-17, 5.79902e-17, 5.799226e-17, 5.799425e-17, 
    5.799863e-17, 5.800347e-17, 5.801035e-17, 5.801536e-17, 5.801871e-17, 
    5.801667e-17, 5.801846e-17, 5.801645e-17, 5.801552e-17, 5.802591e-17, 
    5.802004e-17, 5.802891e-17, 5.802843e-17, 5.802438e-17, 5.802849e-17, 
    5.798913e-17, 5.798802e-17, 5.798406e-17, 5.798716e-17, 5.798157e-17, 
    5.798465e-17, 5.798639e-17, 5.799335e-17, 5.799496e-17, 5.799635e-17, 
    5.799917e-17, 5.800275e-17, 5.800902e-17, 5.801454e-17, 5.801964e-17, 
    5.801928e-17, 5.80194e-17, 5.80205e-17, 5.801772e-17, 5.802096e-17, 
    5.802147e-17, 5.802008e-17, 5.802837e-17, 5.8026e-17, 5.802842e-17, 
    5.802689e-17, 5.798839e-17, 5.799026e-17, 5.798925e-17, 5.799114e-17, 
    5.798977e-17, 5.799576e-17, 5.799755e-17, 5.800606e-17, 5.800266e-17, 
    5.800818e-17, 5.800325e-17, 5.80041e-17, 5.80082e-17, 5.800354e-17, 
    5.801416e-17, 5.800681e-17, 5.802055e-17, 5.801304e-17, 5.8021e-17, 
    5.801962e-17, 5.802196e-17, 5.802401e-17, 5.802666e-17, 5.803145e-17, 
    5.803036e-17, 5.803443e-17, 5.79931e-17, 5.799551e-17, 5.799537e-17, 
    5.799793e-17, 5.799982e-17, 5.8004e-17, 5.801062e-17, 5.800815e-17, 
    5.801276e-17, 5.801367e-17, 5.80067e-17, 5.801091e-17, 5.799717e-17, 
    5.799932e-17, 5.799809e-17, 5.799325e-17, 5.800862e-17, 5.800069e-17, 
    5.801543e-17, 5.801113e-17, 5.80237e-17, 5.801737e-17, 5.802974e-17, 
    5.803485e-17, 5.804001e-17, 5.804565e-17, 5.79969e-17, 5.799525e-17, 
    5.799826e-17, 5.800229e-17, 5.800624e-17, 5.801138e-17, 5.801194e-17, 
    5.801289e-17, 5.801542e-17, 5.801752e-17, 5.801311e-17, 5.801804e-17, 
    5.799967e-17, 5.800935e-17, 5.799457e-17, 5.799892e-17, 5.800209e-17, 
    5.800077e-17, 5.800789e-17, 5.800954e-17, 5.801625e-17, 5.801282e-17, 
    5.803353e-17, 5.802434e-17, 5.80502e-17, 5.80429e-17, 5.799467e-17, 
    5.799693e-17, 5.80047e-17, 5.800101e-17, 5.801176e-17, 5.801438e-17, 
    5.801657e-17, 5.801926e-17, 5.80196e-17, 5.802121e-17, 5.801857e-17, 
    5.802113e-17, 5.801139e-17, 5.801575e-17, 5.80039e-17, 5.800674e-17, 
    5.800546e-17, 5.8004e-17, 5.800849e-17, 5.801317e-17, 5.801339e-17, 
    5.801486e-17, 5.801884e-17, 5.80118e-17, 5.80345e-17, 5.802027e-17, 
    5.799939e-17, 5.800359e-17, 5.800433e-17, 5.800268e-17, 5.801411e-17, 
    5.800995e-17, 5.802118e-17, 5.801817e-17, 5.802314e-17, 5.802066e-17, 
    5.802029e-17, 5.801713e-17, 5.801513e-17, 5.801012e-17, 5.800608e-17, 
    5.800293e-17, 5.800367e-17, 5.800713e-17, 5.801348e-17, 5.801958e-17, 
    5.801823e-17, 5.802276e-17, 5.801098e-17, 5.801585e-17, 5.801393e-17, 
    5.801897e-17, 5.800806e-17, 5.8017e-17, 5.800574e-17, 5.800675e-17, 
    5.800987e-17, 5.801611e-17, 5.801766e-17, 5.801911e-17, 5.801824e-17, 
    5.801366e-17, 5.801297e-17, 5.800982e-17, 5.80089e-17, 5.800654e-17, 
    5.800453e-17, 5.800634e-17, 5.800821e-17, 5.801372e-17, 5.801862e-17, 
    5.802402e-17, 5.802538e-17, 5.803142e-17, 5.802635e-17, 5.803456e-17, 
    5.802734e-17, 5.803997e-17, 5.801769e-17, 5.802736e-17, 5.801005e-17, 
    5.801194e-17, 5.801523e-17, 5.802305e-17, 5.801894e-17, 5.80238e-17, 
    5.801295e-17, 5.800719e-17, 5.800585e-17, 5.80031e-17, 5.800591e-17, 
    5.800568e-17, 5.800837e-17, 5.800751e-17, 5.80139e-17, 5.801047e-17, 
    5.802025e-17, 5.802379e-17, 5.803396e-17, 5.804014e-17, 5.804663e-17, 
    5.804944e-17, 5.80503e-17, 5.805066e-17 ;

 MEG_pinene_a =
  4.796219e-17, 4.796741e-17, 4.796642e-17, 4.797057e-17, 4.796831e-17, 
    4.7971e-17, 4.796329e-17, 4.796758e-17, 4.796487e-17, 4.796272e-17, 
    4.797852e-17, 4.797077e-17, 4.798702e-17, 4.798199e-17, 4.799477e-17, 
    4.798618e-17, 4.799653e-17, 4.799463e-17, 4.80006e-17, 4.799889e-17, 
    4.800633e-17, 4.800139e-17, 4.801036e-17, 4.800521e-17, 4.800597e-17, 
    4.800121e-17, 4.797243e-17, 4.797752e-17, 4.79721e-17, 4.797283e-17, 
    4.797253e-17, 4.796832e-17, 4.796613e-17, 4.796186e-17, 4.796265e-17, 
    4.796583e-17, 4.797316e-17, 4.797074e-17, 4.797705e-17, 4.797691e-17, 
    4.798388e-17, 4.798074e-17, 4.799256e-17, 4.798922e-17, 4.799896e-17, 
    4.79965e-17, 4.799883e-17, 4.799814e-17, 4.799884e-17, 4.799523e-17, 
    4.799677e-17, 4.799362e-17, 4.798131e-17, 4.798489e-17, 4.797416e-17, 
    4.796758e-17, 4.796346e-17, 4.796047e-17, 4.796089e-17, 4.796168e-17, 
    4.796584e-17, 4.796985e-17, 4.797288e-17, 4.797489e-17, 4.797689e-17, 
    4.798268e-17, 4.798597e-17, 4.799318e-17, 4.799197e-17, 4.799409e-17, 
    4.799626e-17, 4.799977e-17, 4.79992e-17, 4.800073e-17, 4.79941e-17, 
    4.799847e-17, 4.799125e-17, 4.799321e-17, 4.797708e-17, 4.797141e-17, 
    4.79687e-17, 4.79666e-17, 4.796121e-17, 4.796491e-17, 4.796344e-17, 
    4.796701e-17, 4.796922e-17, 4.796814e-17, 4.797495e-17, 4.797229e-17, 
    4.798616e-17, 4.798018e-17, 4.7996e-17, 4.799222e-17, 4.799692e-17, 
    4.799454e-17, 4.799859e-17, 4.799495e-17, 4.800132e-17, 4.800267e-17, 
    4.800174e-17, 4.800544e-17, 4.799474e-17, 4.79988e-17, 4.796809e-17, 
    4.796827e-17, 4.796912e-17, 4.796537e-17, 4.796516e-17, 4.796182e-17, 
    4.796482e-17, 4.796607e-17, 4.796938e-17, 4.797127e-17, 4.797309e-17, 
    4.797711e-17, 4.798155e-17, 4.798786e-17, 4.799246e-17, 4.799554e-17, 
    4.799367e-17, 4.799532e-17, 4.799347e-17, 4.799262e-17, 4.800214e-17, 
    4.799676e-17, 4.80049e-17, 4.800447e-17, 4.800075e-17, 4.800452e-17, 
    4.79684e-17, 4.796738e-17, 4.796375e-17, 4.796659e-17, 4.796147e-17, 
    4.796429e-17, 4.796589e-17, 4.797227e-17, 4.797375e-17, 4.797502e-17, 
    4.797761e-17, 4.79809e-17, 4.798664e-17, 4.799171e-17, 4.799639e-17, 
    4.799606e-17, 4.799617e-17, 4.799718e-17, 4.799463e-17, 4.799761e-17, 
    4.799807e-17, 4.79968e-17, 4.80044e-17, 4.800223e-17, 4.800446e-17, 
    4.800305e-17, 4.796772e-17, 4.796944e-17, 4.79685e-17, 4.797025e-17, 
    4.796899e-17, 4.797448e-17, 4.797612e-17, 4.798393e-17, 4.798081e-17, 
    4.798588e-17, 4.798135e-17, 4.798213e-17, 4.79859e-17, 4.798162e-17, 
    4.799136e-17, 4.798462e-17, 4.799722e-17, 4.799034e-17, 4.799765e-17, 
    4.799637e-17, 4.799852e-17, 4.80004e-17, 4.800284e-17, 4.800724e-17, 
    4.800623e-17, 4.800998e-17, 4.797205e-17, 4.797425e-17, 4.797412e-17, 
    4.797648e-17, 4.797821e-17, 4.798204e-17, 4.798812e-17, 4.798585e-17, 
    4.799009e-17, 4.799091e-17, 4.798452e-17, 4.798838e-17, 4.797578e-17, 
    4.797774e-17, 4.797662e-17, 4.797218e-17, 4.798628e-17, 4.7979e-17, 
    4.799253e-17, 4.798859e-17, 4.800013e-17, 4.799431e-17, 4.800567e-17, 
    4.801036e-17, 4.80151e-17, 4.802029e-17, 4.797553e-17, 4.797402e-17, 
    4.797678e-17, 4.798047e-17, 4.79841e-17, 4.798881e-17, 4.798933e-17, 
    4.79902e-17, 4.799252e-17, 4.799445e-17, 4.799041e-17, 4.799493e-17, 
    4.797807e-17, 4.798695e-17, 4.797339e-17, 4.797738e-17, 4.798028e-17, 
    4.797908e-17, 4.798561e-17, 4.798713e-17, 4.799328e-17, 4.799014e-17, 
    4.800915e-17, 4.800071e-17, 4.802446e-17, 4.801776e-17, 4.797348e-17, 
    4.797555e-17, 4.798269e-17, 4.79793e-17, 4.798916e-17, 4.799157e-17, 
    4.799358e-17, 4.799605e-17, 4.799636e-17, 4.799783e-17, 4.799541e-17, 
    4.799776e-17, 4.798882e-17, 4.799282e-17, 4.798195e-17, 4.798455e-17, 
    4.798338e-17, 4.798204e-17, 4.798616e-17, 4.799045e-17, 4.799065e-17, 
    4.799201e-17, 4.799566e-17, 4.79892e-17, 4.801004e-17, 4.799697e-17, 
    4.797781e-17, 4.798167e-17, 4.798235e-17, 4.798083e-17, 4.799132e-17, 
    4.79875e-17, 4.799781e-17, 4.799504e-17, 4.799961e-17, 4.799733e-17, 
    4.799699e-17, 4.799409e-17, 4.799226e-17, 4.798766e-17, 4.798395e-17, 
    4.798106e-17, 4.798174e-17, 4.798491e-17, 4.799074e-17, 4.799634e-17, 
    4.79951e-17, 4.799926e-17, 4.798844e-17, 4.799292e-17, 4.799115e-17, 
    4.799578e-17, 4.798577e-17, 4.799397e-17, 4.798364e-17, 4.798457e-17, 
    4.798743e-17, 4.799315e-17, 4.799458e-17, 4.799591e-17, 4.799511e-17, 
    4.799091e-17, 4.799027e-17, 4.798738e-17, 4.798653e-17, 4.798437e-17, 
    4.798253e-17, 4.798418e-17, 4.79859e-17, 4.799095e-17, 4.799546e-17, 
    4.800041e-17, 4.800167e-17, 4.800721e-17, 4.800255e-17, 4.801009e-17, 
    4.800346e-17, 4.801506e-17, 4.79946e-17, 4.800348e-17, 4.798759e-17, 
    4.798933e-17, 4.799235e-17, 4.799952e-17, 4.799576e-17, 4.800022e-17, 
    4.799025e-17, 4.798497e-17, 4.798373e-17, 4.798122e-17, 4.798379e-17, 
    4.798359e-17, 4.798605e-17, 4.798526e-17, 4.799112e-17, 4.798798e-17, 
    4.799695e-17, 4.800021e-17, 4.800955e-17, 4.801522e-17, 4.802118e-17, 
    4.802376e-17, 4.802455e-17, 4.802488e-17 ;

 MEG_thujene_a =
  1.210192e-18, 1.210318e-18, 1.210294e-18, 1.210395e-18, 1.21034e-18, 
    1.210405e-18, 1.210219e-18, 1.210322e-18, 1.210257e-18, 1.210205e-18, 
    1.210588e-18, 1.2104e-18, 1.210793e-18, 1.210672e-18, 1.210981e-18, 
    1.210773e-18, 1.211024e-18, 1.210978e-18, 1.211123e-18, 1.211081e-18, 
    1.211261e-18, 1.211142e-18, 1.211359e-18, 1.211234e-18, 1.211253e-18, 
    1.211137e-18, 1.21044e-18, 1.210563e-18, 1.210432e-18, 1.21045e-18, 
    1.210442e-18, 1.21034e-18, 1.210287e-18, 1.210184e-18, 1.210203e-18, 
    1.21028e-18, 1.210458e-18, 1.210399e-18, 1.210552e-18, 1.210549e-18, 
    1.210718e-18, 1.210641e-18, 1.210928e-18, 1.210847e-18, 1.211083e-18, 
    1.211023e-18, 1.21108e-18, 1.211063e-18, 1.21108e-18, 1.210992e-18, 
    1.21103e-18, 1.210953e-18, 1.210655e-18, 1.210742e-18, 1.210482e-18, 
    1.210323e-18, 1.210223e-18, 1.21015e-18, 1.21016e-18, 1.21018e-18, 
    1.210281e-18, 1.210378e-18, 1.210451e-18, 1.2105e-18, 1.210548e-18, 
    1.210688e-18, 1.210768e-18, 1.210943e-18, 1.210913e-18, 1.210965e-18, 
    1.211017e-18, 1.211102e-18, 1.211089e-18, 1.211126e-18, 1.210965e-18, 
    1.211071e-18, 1.210896e-18, 1.210944e-18, 1.210553e-18, 1.210415e-18, 
    1.21035e-18, 1.210299e-18, 1.210168e-18, 1.210258e-18, 1.210222e-18, 
    1.210309e-18, 1.210362e-18, 1.210336e-18, 1.210501e-18, 1.210437e-18, 
    1.210773e-18, 1.210628e-18, 1.211011e-18, 1.21092e-18, 1.211033e-18, 
    1.210976e-18, 1.211074e-18, 1.210986e-18, 1.21114e-18, 1.211173e-18, 
    1.21115e-18, 1.21124e-18, 1.210981e-18, 1.211079e-18, 1.210335e-18, 
    1.210339e-18, 1.21036e-18, 1.210269e-18, 1.210264e-18, 1.210183e-18, 
    1.210256e-18, 1.210286e-18, 1.210366e-18, 1.210412e-18, 1.210456e-18, 
    1.210553e-18, 1.210661e-18, 1.210814e-18, 1.210925e-18, 1.211e-18, 
    1.210955e-18, 1.210995e-18, 1.21095e-18, 1.210929e-18, 1.21116e-18, 
    1.21103e-18, 1.211227e-18, 1.211216e-18, 1.211126e-18, 1.211218e-18, 
    1.210342e-18, 1.210318e-18, 1.21023e-18, 1.210299e-18, 1.210174e-18, 
    1.210243e-18, 1.210282e-18, 1.210436e-18, 1.210472e-18, 1.210503e-18, 
    1.210566e-18, 1.210645e-18, 1.210784e-18, 1.210907e-18, 1.211021e-18, 
    1.211013e-18, 1.211015e-18, 1.21104e-18, 1.210978e-18, 1.21105e-18, 
    1.211061e-18, 1.211031e-18, 1.211215e-18, 1.211162e-18, 1.211216e-18, 
    1.211182e-18, 1.210326e-18, 1.210368e-18, 1.210345e-18, 1.210387e-18, 
    1.210357e-18, 1.21049e-18, 1.21053e-18, 1.210719e-18, 1.210643e-18, 
    1.210766e-18, 1.210656e-18, 1.210675e-18, 1.210766e-18, 1.210663e-18, 
    1.210899e-18, 1.210735e-18, 1.211041e-18, 1.210874e-18, 1.211051e-18, 
    1.21102e-18, 1.211072e-18, 1.211118e-18, 1.211177e-18, 1.211283e-18, 
    1.211259e-18, 1.21135e-18, 1.210431e-18, 1.210484e-18, 1.210481e-18, 
    1.210538e-18, 1.21058e-18, 1.210673e-18, 1.21082e-18, 1.210765e-18, 
    1.210868e-18, 1.210888e-18, 1.210733e-18, 1.210827e-18, 1.210521e-18, 
    1.210569e-18, 1.210542e-18, 1.210434e-18, 1.210776e-18, 1.210599e-18, 
    1.210927e-18, 1.210831e-18, 1.211111e-18, 1.21097e-18, 1.211245e-18, 
    1.211359e-18, 1.211474e-18, 1.2116e-18, 1.210515e-18, 1.210479e-18, 
    1.210545e-18, 1.210635e-18, 1.210723e-18, 1.210837e-18, 1.21085e-18, 
    1.210871e-18, 1.210927e-18, 1.210973e-18, 1.210876e-18, 1.210985e-18, 
    1.210577e-18, 1.210792e-18, 1.210463e-18, 1.21056e-18, 1.21063e-18, 
    1.210601e-18, 1.210759e-18, 1.210796e-18, 1.210945e-18, 1.210869e-18, 
    1.21133e-18, 1.211125e-18, 1.211701e-18, 1.211538e-18, 1.210465e-18, 
    1.210516e-18, 1.210689e-18, 1.210607e-18, 1.210845e-18, 1.210904e-18, 
    1.210953e-18, 1.211012e-18, 1.21102e-18, 1.211056e-18, 1.210997e-18, 
    1.211054e-18, 1.210837e-18, 1.210934e-18, 1.210671e-18, 1.210734e-18, 
    1.210705e-18, 1.210673e-18, 1.210773e-18, 1.210877e-18, 1.210882e-18, 
    1.210914e-18, 1.211003e-18, 1.210847e-18, 1.211351e-18, 1.211035e-18, 
    1.21057e-18, 1.210664e-18, 1.21068e-18, 1.210644e-18, 1.210898e-18, 
    1.210805e-18, 1.211055e-18, 1.210988e-18, 1.211099e-18, 1.211043e-18, 
    1.211035e-18, 1.210965e-18, 1.210921e-18, 1.210809e-18, 1.210719e-18, 
    1.210649e-18, 1.210666e-18, 1.210743e-18, 1.210884e-18, 1.211019e-18, 
    1.210989e-18, 1.21109e-18, 1.210828e-18, 1.210936e-18, 1.210894e-18, 
    1.211006e-18, 1.210763e-18, 1.210962e-18, 1.210712e-18, 1.210734e-18, 
    1.210803e-18, 1.210942e-18, 1.210977e-18, 1.211009e-18, 1.21099e-18, 
    1.210888e-18, 1.210872e-18, 1.210802e-18, 1.210782e-18, 1.210729e-18, 
    1.210685e-18, 1.210725e-18, 1.210766e-18, 1.210889e-18, 1.210998e-18, 
    1.211118e-18, 1.211149e-18, 1.211283e-18, 1.21117e-18, 1.211353e-18, 
    1.211192e-18, 1.211473e-18, 1.210977e-18, 1.211192e-18, 1.210807e-18, 
    1.210849e-18, 1.210923e-18, 1.211097e-18, 1.211005e-18, 1.211113e-18, 
    1.210872e-18, 1.210744e-18, 1.210714e-18, 1.210653e-18, 1.210715e-18, 
    1.21071e-18, 1.21077e-18, 1.210751e-18, 1.210893e-18, 1.210817e-18, 
    1.211034e-18, 1.211113e-18, 1.211339e-18, 1.211477e-18, 1.211621e-18, 
    1.211684e-18, 1.211703e-18, 1.211711e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  3.681014e-25, 1.703156e-25, 2.032799e-25, 3.543663e-25, 2.994258e-25, 
    1.071341e-25, 1.538335e-25, -2.142679e-25, -7.966364e-26, -2.142679e-25, 
    3.104139e-25, -3.681012e-25, 1.208692e-25, -6.043446e-26, 6.86757e-26, 
    3.763425e-25, 1.648223e-26, 2.005329e-25, -3.351369e-25, -2.692083e-25, 
    3.296438e-26, -4.50512e-25, 1.373521e-26, 3.845835e-25, 7.416975e-26, 
    -4.093066e-25, -1.977857e-25, -3.296421e-26, 2.472331e-26, -1.922916e-25, 
    4.257889e-25, -9.339876e-26, 1.538335e-25, -8.515768e-26, 4.917175e-25, 
    2.032799e-25, -1.318571e-25, -1.126279e-25, 3.104139e-25, 2.609674e-25, 
    3.021735e-26, -1.703155e-25, -1.922916e-25, -4.972114e-25, 2.14268e-25, 
    -1.098809e-25, -5.136936e-25, -3.571124e-26, 2.637145e-25, -1.703155e-25, 
    -2.33497e-25, -4.120529e-26, -4.752352e-25, -1.483393e-25, -2.582203e-25, 
    3.323901e-25, -9.614578e-26, 2.08774e-25, -3.104137e-25, -4.944636e-26, 
    2.856907e-25, -1.593274e-25, 3.983187e-25, -2.719554e-25, -4.56006e-25, 
    4.148008e-25, 2.856907e-25, -1.922916e-25, -2.719554e-25, -2.33497e-25, 
    -2.801964e-25, 5.76876e-26, 4.120545e-26, 8.241083e-26, -1.593274e-25, 
    -2.115208e-25, 1.098818e-26, -2.692083e-25, -2.774494e-25, 3.790895e-25, 
    8.241083e-26, 2.939317e-25, 1.0164e-25, 2.801966e-25, 1.318573e-25, 
    3.57114e-26, 2.966788e-25, -1.318571e-25, 6.318165e-26, 1.236162e-25, 
    4.669943e-25, 1.538335e-25, 8.241157e-27, -3.104137e-25, -9.339876e-26, 
    2.472331e-26, -1.098809e-25, 1.373521e-26, 5.384169e-25, -2.389911e-25, 
    1.922926e-26, -3.351369e-25, 1.922918e-25, 1.0164e-25, -2.472314e-26, 
    1.263632e-25, -2.417381e-25, -4.669941e-25, -3.241488e-25, 1.785567e-25, 
    -1.648207e-26, -1.538333e-25, -3.818364e-25, 1.236162e-25, -3.571131e-25, 
    1.071341e-25, -4.120529e-26, -1.895446e-25, -5.493967e-27, -2.692083e-25, 
    -3.131607e-25, -1.23616e-25, -1.18122e-25, -1.346041e-25, 1.593275e-25, 
    -4.395231e-26, -2.884375e-25, -7.691661e-26, -2.142679e-25, 3.681014e-25, 
    2.856907e-25, -4.120529e-26, 1.785567e-25, -4.752352e-25, -2.25256e-25, 
    7.691677e-26, -6.592851e-26, 1.483394e-25, -2.746942e-27, -1.098809e-25, 
    -3.708483e-25, -5.219339e-26, 2.719555e-25, -1.428452e-25, -1.758095e-25, 
    -1.071339e-25, -4.944636e-26, -3.268959e-25, 7.96638e-26, 2.747026e-25, 
    1.346043e-25, -1.895446e-25, 6.043463e-26, 1.840507e-25, 9.614595e-26, 
    -4.615001e-25, -3.488721e-25, -2.637143e-25, -2.637143e-25, 3.873306e-25, 
    -3.296429e-25, -9.065174e-26, -3.021719e-26, 7.416975e-26, -1.648214e-25, 
    -8.515768e-26, 2.747107e-27, 2.527264e-25, -1.18122e-25, -2.554732e-25, 
    2.11521e-25, -1.18122e-25, 9.339892e-26, -5.164406e-25, 2.884377e-25, 
    -7.142256e-26, -6.373097e-25, 4.66995e-26, -3.351369e-25, -2.3075e-25, 
    2.225091e-25, -1.291101e-25, -6.867554e-26, 2.005329e-25, -2.747016e-26, 
    3.873306e-25, -3.186548e-25, 1.071341e-25, 2.252561e-25, 2.472323e-25, 
    -5.274287e-25, -6.73021e-25, 2.747107e-27, 1.373513e-25, 3.433782e-25, 
    -5.493967e-27, 1.400983e-25, -8.515768e-26, -1.098809e-25, -7.691661e-26, 
    1.0164e-25, 1.153751e-25, -2.142679e-25, -4.752352e-25, -2.115208e-25, 
    -5.878632e-25, -3.598602e-25, 1.373521e-26, 1.730626e-25, -9.889281e-26, 
    3.296431e-25, -1.785565e-25, -1.071339e-25, 6.86757e-26, -2.472314e-26, 
    -5.439108e-25, -6.043446e-26, 2.719555e-25, 2.582204e-25, 2.389912e-25, 
    -6.812621e-25, -1.922909e-26, 2.747107e-27, 8.257634e-32, -2.115208e-25, 
    -3.076667e-25, -5.521519e-25, 8.790487e-26, -9.889281e-26, -4.120529e-26, 
    -5.384168e-25, 1.126281e-25, -2.142679e-25, -2.966786e-25, -2.197612e-26, 
    2.499793e-25, -2.856905e-25, 7.142273e-26, -4.642471e-25, 1.098811e-25, 
    -3.104137e-25, 2.252561e-25, -3.735953e-25, 3.900776e-25, -2.692083e-25, 
    5.494058e-26, -3.763423e-25, 8.515785e-26, 7.691677e-26, -5.768744e-26, 
    -1.675684e-25, -6.043446e-26, -2.911845e-25, 2.884377e-25, -9.587115e-25, 
    -4.752352e-25, -1.648207e-26, 2.582204e-25, -1.922916e-25, -1.538333e-25, 
    1.648223e-26, 2.197628e-26, -1.785565e-25, 4.477651e-25, -1.043869e-25, 
    5.76876e-26, 2.472323e-25, 3.296431e-25, -1.593274e-25, -1.346041e-25, 
    2.637145e-25, -1.620744e-25, -2.554732e-25, 2.747107e-27, -1.126279e-25, 
    4.148008e-25, 2.829436e-25, -1.428452e-25, 1.565805e-25, -7.691661e-26, 
    3.24149e-25, 3.516192e-25, -1.23616e-25, -3.241488e-25, 2.14268e-25, 
    -4.395239e-25, -6.043446e-26, -2.197612e-26, -1.400982e-25, 
    -1.373512e-25, -5.384168e-25, 2.609674e-25, 1.758097e-25, 9.889298e-26, 
    -3.571131e-25, 7.142273e-26, -3.268959e-25, 1.0164e-25, 3.104139e-25, 
    2.472331e-26, -2.856905e-25, -2.087738e-25, -2.28003e-25, -5.576459e-25, 
    1.236162e-25, -1.648214e-25, 1.098818e-26, 1.373521e-26, 2.08774e-25, 
    -1.675684e-25, 2.14268e-25, 9.889298e-26, 1.428454e-25, -6.043446e-26, 
    7.142273e-26, -4.010655e-25, -4.450179e-25, 1.785567e-25, 3.351371e-25, 
    7.96638e-26, -3.296429e-25, -2.609673e-25, -1.15375e-25, 1.758097e-25, 
    -1.867976e-25, 5.136937e-25, 9.889298e-26, 1.263632e-25, -2.582203e-25, 
    1.648216e-25, -1.455922e-25, -2.747016e-26, 1.098818e-26, 2.609674e-25, 
    -3.37884e-25, 3.406311e-25, -3.845826e-26, -5.494041e-26 ;

 M_LITR2C_TO_LEACHING =
  -2.939316e-25, -2.637143e-25, -1.758095e-25, -8.515771e-26, -1.648209e-26, 
    -1.895447e-25, -3.845829e-26, -8.241069e-26, -1.20869e-25, 1.263632e-25, 
    -8.241069e-26, 1.813037e-25, 1.922923e-26, 6.04346e-26, 2.747078e-27, 
    2.087739e-25, -1.565804e-25, 1.400983e-25, -2.444852e-25, 3.928246e-25, 
    -7.142259e-26, -1.236161e-25, 1.64822e-26, -1.593274e-25, 1.181221e-25, 
    -3.296424e-26, 3.84584e-26, 2.14268e-25, -1.318571e-25, 8.24108e-26, 
    -1.977857e-25, -4.395234e-26, 1.64822e-26, -2.197614e-26, -2.444852e-25, 
    -6.043449e-26, 3.104139e-25, 7.416973e-26, 1.373513e-25, 5.494055e-26, 
    1.04387e-25, -3.845829e-26, -1.20869e-25, -7.966367e-26, -5.494044e-26, 
    2.856906e-25, -1.291101e-25, 2.472323e-25, 6.592865e-26, 2.472328e-26, 
    -9.065177e-26, -1.593274e-25, 3.488722e-25, -1.263631e-25, -1.15375e-25, 
    -6.592854e-26, 2.14268e-25, -3.296424e-26, -1.950387e-25, -1.263631e-25, 
    3.076668e-25, -3.845829e-26, 4.94465e-26, 4.120543e-26, -1.18122e-25, 
    5.768757e-26, 7.416973e-26, -9.339879e-26, -6.043449e-26, -6.592854e-26, 
    -7.416961e-26, -2.966786e-25, -3.571127e-26, 4.94465e-26, -1.291101e-25, 
    -7.142259e-26, -1.20869e-25, 1.236162e-25, -1.648214e-25, -9.339879e-26, 
    2.747025e-25, -7.416961e-26, 3.26896e-25, -5.493996e-27, -1.648209e-26, 
    -3.488721e-25, 5.494055e-26, 7.416973e-26, -1.043869e-25, -1.318571e-25, 
    -3.955715e-25, -6.043449e-26, 1.263632e-25, -9.065177e-26, -5.494044e-26, 
    2.472323e-25, 5.494103e-27, -2.142679e-25, 8.515782e-26, -8.790474e-26, 
    -1.043869e-25, 4.94465e-26, 1.09881e-25, -4.395234e-26, -1.977857e-25, 
    1.565805e-25, -2.197614e-26, 1.64822e-26, -2.966786e-25, -1.730625e-25, 
    -8.241021e-27, 5.494055e-26, -4.010656e-25, 6.867567e-26, -8.241069e-26, 
    -3.296424e-26, 2.417382e-25, 5.768757e-26, 3.818365e-25, 1.648215e-25, 
    3.021733e-26, -3.845829e-26, 1.318572e-25, -9.614581e-26, -1.758095e-25, 
    -3.296424e-26, -1.648209e-26, -1.922912e-26, 2.14268e-25, 8.515782e-26, 
    1.373513e-25, -1.483393e-25, 1.703156e-25, 5.768757e-26, -9.889284e-26, 
    1.565805e-25, -2.637143e-25, 5.494055e-26, 3.84584e-26, 2.252561e-25, 
    -1.648209e-26, 2.17015e-25, -1.867976e-25, -6.043449e-26, -1.730625e-25, 
    1.64822e-26, -1.346042e-25, -2.087738e-25, 1.922923e-26, -5.493996e-27, 
    -3.571132e-25, 9.339889e-26, 8.790485e-26, 1.208691e-25, 1.675686e-25, 
    7.14227e-26, 9.339889e-26, 5.494055e-26, -2.472317e-26, -1.977857e-25, 
    -1.922917e-25, -9.339879e-26, 8.24108e-26, 1.455924e-25, 3.84584e-26, 
    1.867977e-25, -4.065596e-25, 3.3239e-25, 1.758096e-25, -8.790474e-26, 
    -8.790474e-26, 8.241128e-27, 1.04387e-25, 1.840507e-25, -2.74702e-26, 
    1.867977e-25, -2.334971e-25, -1.318571e-25, -4.038126e-25, 5.494103e-27, 
    4.395245e-26, 2.14268e-25, 1.373518e-26, 1.64822e-26, 1.098815e-26, 
    2.362442e-25, -4.395234e-26, 2.499793e-25, -9.065177e-26, -2.362441e-25, 
    -9.889284e-26, 2.032799e-25, -1.043869e-25, -5.494044e-26, 6.592865e-26, 
    -1.016399e-25, 9.339889e-26, -1.20869e-25, -4.120537e-25, -1.675685e-25, 
    -7.142259e-26, -1.538333e-25, 8.515782e-26, 1.703156e-25, -2.499792e-25, 
    -1.675685e-25, -4.944639e-26, 3.021733e-26, -4.944639e-26, -4.395234e-26, 
    7.14227e-26, -5.494044e-26, 7.416973e-26, 1.538334e-25, 1.208691e-25, 
    6.592865e-26, -6.592854e-26, -3.845829e-26, 1.318572e-25, 7.14227e-26, 
    1.400983e-25, -2.060268e-25, 2.307501e-25, 2.527263e-25, 3.84584e-26, 
    6.04346e-26, -1.236161e-25, -9.339879e-26, 1.0164e-25, 3.186549e-25, 
    -3.845834e-25, 2.307501e-25, 3.021728e-25, -4.395234e-26, 1.977858e-25, 
    1.64822e-26, -2.472317e-26, -5.768747e-26, -6.592854e-26, -5.494044e-26, 
    3.29643e-25, -1.043869e-25, -8.241069e-26, 7.14227e-26, 9.065187e-26, 
    -2.25256e-25, -6.318152e-26, -1.016399e-25, -1.373512e-25, 6.592865e-26, 
    -1.813036e-25, 1.400983e-25, 1.098815e-26, -1.758095e-25, -1.098805e-26, 
    -2.3075e-25, -3.021722e-26, -1.400982e-25, 1.126281e-25, 1.922918e-25, 
    1.291102e-25, -1.071339e-25, -1.318571e-25, -3.543661e-25, 2.444853e-25, 
    8.24108e-26, 1.675686e-25, 8.24108e-26, 5.351442e-32, -1.346042e-25, 
    8.790485e-26, 2.747078e-27, 1.126281e-25, 3.26896e-25, 1.64822e-26, 
    2.11521e-25, 6.592865e-26, -1.400982e-25, 5.768757e-26, 1.565805e-25, 
    5.494055e-26, -1.510863e-25, 2.939317e-25, -1.483393e-25, 5.351451e-32, 
    3.516192e-25, -3.845829e-26, 4.120543e-26, -3.571127e-26, 2.19762e-25, 
    -3.268959e-25, 2.74703e-26, -4.862233e-25, -2.197614e-26, 6.867567e-26, 
    -8.515771e-26, -2.087738e-25, -2.170149e-25, -5.494044e-26, 
    -3.900775e-25, -1.648209e-26, 3.131609e-25, 1.263632e-25, 3.21402e-25, 
    -2.362441e-25, 6.04346e-26, 7.966377e-26, -6.043449e-26, 1.373518e-26, 
    1.730626e-25, 1.236162e-25, -2.719554e-25, -1.20869e-25, -1.758095e-25, 
    -1.098805e-26, 1.373513e-25, 4.395245e-26, -1.648209e-26, -9.889284e-26, 
    1.785567e-25, 4.395245e-26, -7.142259e-26, 2.005329e-25, 1.318572e-25, 
    -1.785566e-25, 6.318163e-26, -2.25256e-25, 1.181221e-25, -9.614581e-26, 
    -1.373512e-25, -7.966367e-26, 1.922923e-26, 2.087739e-25, -1.016399e-25, 
    4.120543e-26, -1.648214e-25, 1.291102e-25, 2.19762e-25 ;

 M_LITR3C_TO_LEACHING =
  2.334974e-26, -2.197617e-26, -2.197617e-26, 4.257891e-26, -6.867559e-26, 
    4.395242e-26, -3.159076e-26, -1.332307e-25, -4.120535e-26, -9.614584e-26, 
    -3.021725e-26, 4.12054e-26, -1.085074e-25, -1.648212e-26, -1.387247e-25, 
    -9.339881e-26, 1.208691e-25, -7.416964e-26, -5.768749e-26, -6.043452e-26, 
    -1.071339e-25, -1.922915e-26, -7.00491e-26, -9.61456e-27, -6.180803e-26, 
    -1.607009e-25, -7.966369e-26, -2.197617e-26, 7.691672e-26, 2.197622e-26, 
    6.043457e-26, -2.609671e-26, 1.414718e-25, -3.708481e-26, -5.768749e-26, 
    4.12054e-26, 2.197622e-26, -9.065179e-26, -7.554316e-26, -6.867559e-26, 
    -1.263631e-25, -1.648212e-26, -5.494047e-26, -2.197617e-26, 
    -1.565804e-25, 5.494052e-26, 2.675721e-32, 1.510864e-25, 1.510866e-26, 
    -2.884373e-26, -2.884373e-26, 6.592862e-26, 2.67573e-32, -4.669939e-26, 
    -4.532588e-26, 1.373539e-27, 9.339887e-26, -8.241071e-26, 2.747028e-26, 
    4.12054e-26, -5.356696e-26, 2.334974e-26, 1.359778e-25, 9.614614e-27, 
    -2.115209e-25, 2.675729e-32, -1.785563e-26, 5.906106e-26, 2.472325e-26, 
    -6.043452e-26, -4.807291e-26, 3.296432e-26, -2.060266e-26, 2.67572e-32, 
    -4.120511e-27, 1.373539e-27, 6.867589e-27, -1.414718e-25, -1.194956e-25, 
    2.060271e-26, 7.416969e-26, 3.571135e-26, -2.746998e-27, -2.47232e-26, 
    2.675739e-32, -3.845832e-26, 9.202536e-26, -1.071339e-25, -5.494023e-27, 
    5.494076e-27, -1.373486e-27, -1.167485e-25, 6.867589e-27, 3.708486e-26, 
    2.472325e-26, 1.373539e-27, 1.098813e-26, 5.494052e-26, -4.120535e-26, 
    4.257891e-26, 1.63448e-25, 2.747028e-26, -5.494047e-26, -4.944642e-26, 
    7.142267e-26, 1.648217e-26, -8.241071e-26, 2.005328e-25, -1.593274e-25, 
    1.236164e-26, 1.04387e-25, -4.532588e-26, 2.060271e-26, 5.631404e-26, 
    -4.807291e-26, -1.922915e-26, -2.746998e-27, -9.339881e-26, 1.92292e-26, 
    1.510864e-25, 1.181221e-25, 1.263632e-25, 8.653131e-26, -1.469658e-25, 
    -4.944642e-26, 4.807296e-26, -4.669939e-26, -7.829018e-26, -1.359777e-25, 
    -9.065179e-26, -4.120535e-26, 1.387248e-25, 2.747052e-27, 3.159081e-26, 
    6.043457e-26, -5.081993e-26, -4.120535e-26, 1.277367e-25, 6.043457e-26, 
    1.236164e-26, -1.37351e-26, 3.433784e-26, -1.291101e-25, -1.497128e-25, 
    -3.296427e-26, 3.433784e-26, -5.494047e-26, 3.845837e-26, -1.359777e-25, 
    -4.395237e-26, 1.92292e-26, 1.167486e-25, -5.768749e-26, -4.944642e-26, 
    -1.09881e-25, 2.472325e-26, -9.614584e-26, -8.10372e-26, -1.387247e-25, 
    5.768755e-26, 2.197622e-26, -1.12628e-25, -2.197617e-26, -6.043452e-26, 
    6.867589e-27, -4.120535e-26, 4.532594e-26, -6.730208e-26, 9.339887e-26, 
    -1.071339e-25, 2.747028e-26, 3.159081e-26, -1.098807e-26, -1.922915e-26, 
    4.669945e-26, 1.098813e-26, -2.142679e-25, -7.829018e-26, -6.867559e-26, 
    6.455511e-26, -9.065179e-26, 1.12628e-25, -2.334968e-26, 1.04387e-25, 
    6.31816e-26, 9.339887e-26, -1.222426e-25, 3.845837e-26, -4.669939e-26, 
    2.22509e-25, 2.675725e-32, 5.21935e-26, -1.140015e-25, -2.746998e-27, 
    -3.433778e-26, -9.751935e-26, -2.884373e-26, 7.142267e-26, -3.57113e-26, 
    -2.087739e-25, -1.263631e-25, 3.845837e-26, -5.906101e-26, 9.75194e-26, 
    -1.414718e-25, 6.867589e-27, 4.12054e-26, -1.016399e-25, 5.631404e-26, 
    5.494076e-27, 1.208691e-25, -2.005328e-25, -1.098807e-26, -1.030134e-25, 
    -1.785563e-26, -7.416964e-26, 1.373515e-26, 5.494052e-26, 2.472325e-26, 
    -3.983183e-26, -1.15375e-25, -4.944642e-26, -3.021725e-26, -7.966369e-26, 
    -1.826771e-25, 5.631404e-26, -7.554316e-26, -9.20253e-26, -3.57113e-26, 
    3.845837e-26, 6.592862e-26, -1.359777e-25, -1.964122e-25, 5.21935e-26, 
    -2.609671e-26, -1.538334e-25, -7.00491e-26, -3.296427e-26, -4.669939e-26, 
    1.648215e-25, -1.37351e-26, 7.279618e-26, 3.296432e-26, 2.747052e-27, 
    -2.884373e-26, -7.416964e-26, -2.884373e-26, 3.296432e-26, 1.648217e-26, 
    -2.884373e-26, -2.060266e-26, -6.043452e-26, 7.829024e-26, -4.807291e-26, 
    -1.043869e-25, 3.571135e-26, 4.257891e-26, -1.071339e-25, 1.675685e-25, 
    -2.334971e-25, 8.378428e-26, 9.065185e-26, -1.785566e-25, 5.906106e-26, 
    -3.983183e-26, 3.433784e-26, -2.115209e-25, 9.065185e-26, 7.691672e-26, 
    8.241101e-27, 2.747052e-27, -2.060266e-26, -3.296427e-26, -5.494047e-26, 
    -2.060266e-26, -1.002664e-25, -4.257886e-26, 6.592862e-26, -5.494023e-27, 
    2.884379e-26, 5.906106e-26, -7.966369e-26, -1.15375e-25, -1.922915e-26, 
    5.081998e-26, -7.142262e-26, -1.510863e-25, 3.571135e-26, 1.785569e-26, 
    -7.279613e-26, 1.428453e-25, 7.004916e-26, 5.768755e-26, -1.030134e-25, 
    -1.510863e-25, 2.609676e-26, -4.669939e-26, 2.334974e-26, 7.004916e-26, 
    7.691672e-26, 9.614589e-26, -5.494047e-26, 2.747028e-26, 1.648217e-26, 
    4.12054e-26, 1.263632e-25, -3.983183e-26, -1.840506e-25, -9.065179e-26, 
    -1.373512e-25, 2.675718e-32, -1.277366e-25, 2.472325e-26, 4.532594e-26, 
    1.002664e-25, 2.472325e-26, -1.304836e-25, -4.395237e-26, -5.219344e-26, 
    -3.296427e-26, 1.648217e-26, 3.02173e-26, -5.631398e-26, -2.334971e-25, 
    8.515779e-26, 1.12628e-25, 5.768755e-26, -1.167485e-25, 3.159081e-26, 
    7.554321e-26, -3.708481e-26, -1.66195e-25, 1.016399e-25, -5.219344e-26, 
    1.813037e-25, -3.021725e-26, 3.845837e-26, -1.098807e-26 ;

 M_SOIL1C_TO_LEACHING =
  -4.552245e-21, -1.737775e-20, -1.616201e-20, -2.244318e-21, 2.654419e-20, 
    5.325241e-21, -2.988691e-20, 3.373262e-21, 7.2416e-21, -1.123544e-20, 
    4.592566e-20, -1.225214e-20, 2.33308e-21, 1.85658e-20, 4.193725e-21, 
    2.594166e-20, 1.91577e-21, -1.499096e-20, -3.753677e-20, -3.857044e-20, 
    1.019585e-20, 1.822509e-20, 2.932483e-20, -1.284389e-20, 4.568989e-22, 
    1.895906e-20, -2.475534e-20, 1.294286e-20, 8.670793e-21, 2.877095e-20, 
    -9.759013e-21, 1.707836e-20, -1.944708e-20, 6.757546e-21, 1.23822e-20, 
    -1.457477e-20, 4.127784e-20, 1.939166e-20, -1.53192e-20, -1.190568e-21, 
    2.430776e-20, -1.618435e-20, -3.115981e-21, -4.33625e-21, -9.05614e-21, 
    1.701192e-20, -1.575654e-21, 1.421203e-20, -1.805633e-20, 7.442866e-21, 
    -4.582947e-22, -2.422833e-20, -2.988691e-20, -2.27095e-20, -2.165713e-21, 
    -2.407058e-20, -3.05044e-20, 3.615337e-20, 1.571813e-20, -3.856276e-20, 
    1.03075e-20, 9.166702e-21, 1.651205e-20, 2.599851e-20, -9.90681e-22, 
    2.220283e-21, 1.648237e-20, 6.936515e-21, -1.180627e-20, 9.677044e-21, 
    -7.396517e-21, 2.564735e-20, 1.504135e-21, 2.10462e-20, -1.380179e-20, 
    -6.712593e-21, 3.769792e-20, -1.264174e-20, -3.91537e-20, -1.036663e-20, 
    1.271808e-20, 5.394574e-22, 6.691954e-21, -1.358295e-20, 4.298186e-20, 
    2.691617e-21, 2.10329e-20, 9.12343e-21, -2.596968e-20, -4.224959e-20, 
    -3.176877e-20, 1.52952e-20, -1.439636e-20, 7.387552e-22, -1.123007e-20, 
    4.210398e-20, -4.772298e-20, -4.351821e-20, 3.230476e-21, 9.112417e-21, 
    -2.892621e-21, 2.13832e-20, 9.499749e-22, -1.068636e-20, 6.788081e-21, 
    7.82316e-21, -1.75296e-20, 1.82758e-21, -1.736365e-20, 1.165923e-20, 
    -2.043944e-20, -1.591208e-20, -7.791942e-22, -2.305811e-20, 
    -1.722226e-20, -3.853393e-20, -1.729241e-20, 3.944264e-20, 3.279969e-21, 
    -7.975562e-21, -3.107783e-21, -7.097679e-21, -1.488097e-20, 
    -7.863866e-21, 1.399321e-20, 3.735724e-21, 2.697307e-20, -1.200333e-20, 
    -4.610489e-21, 1.778007e-20, 1.042996e-20, -3.264807e-20, 3.245778e-20, 
    -3.573038e-20, -2.260404e-20, 1.70922e-20, 4.286539e-20, 1.54405e-20, 
    2.75561e-20, 3.103762e-20, -1.012684e-20, 4.2264e-20, 5.540138e-20, 
    -7.766671e-20, 2.024323e-20, -8.018239e-22, 1.443823e-20, -3.253609e-20, 
    2.208159e-20, -2.462757e-20, 4.849285e-20, 1.304972e-20, 2.341266e-20, 
    -2.324924e-20, -1.426688e-20, -1.230925e-20, -2.318817e-20, 
    -1.114807e-20, 3.45666e-21, 2.660921e-20, 7.888111e-22, -1.718014e-20, 
    6.408098e-21, -1.098466e-20, 2.467668e-21, -2.817384e-20, 1.34803e-20, 
    -7.843226e-21, 2.572341e-20, -4.74377e-20, 5.030624e-21, -1.794634e-20, 
    3.14846e-20, 3.76015e-22, 2.72332e-20, -3.851388e-21, 7.267257e-20, 
    -1.435481e-20, 4.351338e-20, -9.521817e-21, 1.354845e-20, 5.159526e-20, 
    2.970227e-20, 8.091888e-22, -1.595224e-20, -1.607266e-20, 1.342407e-20, 
    3.380358e-20, -8.520079e-21, -2.614072e-20, 1.023035e-20, 8.985756e-21, 
    -5.243533e-21, -3.382022e-21, 7.953421e-22, -1.352302e-20, -2.062152e-20, 
    1.881264e-20, -2.324319e-21, -7.456172e-21, -2.307732e-20, 4.762582e-21, 
    -8.700192e-21, 1.451426e-20, -1.917707e-20, -1.465987e-20, -1.599097e-20, 
    -4.249443e-20, 1.179005e-22, -2.224045e-20, 8.224344e-21, 1.24639e-20, 
    -1.61035e-20, 1.943547e-20, -8.980653e-21, 1.129198e-20, 6.306044e-21, 
    -2.812972e-20, 2.462565e-21, -2.588289e-20, 5.869212e-21, 8.871824e-21, 
    -7.215579e-21, 2.226308e-20, -2.904747e-20, -2.277311e-20, 6.372761e-21, 
    2.551956e-20, 1.87637e-20, 1.661525e-20, -1.835768e-21, -4.568618e-20, 
    -6.03743e-21, -5.685719e-21, -1.074207e-20, 1.091765e-20, -1.545096e-20, 
    -6.246933e-21, 1.123204e-20, 1.427865e-22, -1.887652e-20, 2.741443e-20, 
    3.143656e-20, 2.660469e-20, 7.644474e-21, -6.873757e-21, 3.560712e-20, 
    4.181595e-21, -1.456855e-20, 4.119382e-21, 1.11508e-21, 3.633939e-20, 
    -1.782901e-20, -3.803831e-20, -1.903711e-20, 3.058468e-20, 1.785556e-20, 
    4.773032e-20, -6.484981e-21, -3.824699e-20, -2.732029e-21, 2.498914e-20, 
    1.880331e-20, 1.138105e-20, -5.241254e-21, 5.198146e-20, -2.92434e-20, 
    9.142934e-21, 5.205062e-21, 4.826272e-20, -4.400987e-20, -2.634401e-20, 
    3.162316e-20, 4.158601e-20, -2.435442e-20, -1.071918e-20, 5.952343e-21, 
    8.979508e-22, -2.780713e-20, -2.267642e-20, 4.667028e-21, 3.843714e-21, 
    4.39958e-21, 6.544091e-21, 2.015561e-20, -3.144419e-20, -4.851082e-21, 
    1.667551e-21, -1.616232e-20, 5.81661e-21, -5.007999e-21, 3.216639e-21, 
    -2.178863e-20, 2.406548e-20, -6.020187e-21, -1.363835e-20, 2.134278e-20, 
    8.721111e-21, -1.55236e-20, 9.267905e-21, 4.227533e-20, -2.252319e-20, 
    7.837863e-21, 3.548103e-20, 2.301655e-20, 1.743911e-20, 2.656232e-21, 
    -6.93538e-21, -6.83361e-22, -2.927676e-20, 8.008359e-21, 4.943774e-20, 
    1.08221e-20, -1.928157e-22, 3.096638e-20, -2.654789e-22, -4.032309e-21, 
    -3.357174e-20, -7.695998e-22, 1.605541e-20, -1.103638e-20, -2.224526e-20, 
    1.036663e-20, 1.221595e-20, -4.185536e-21, -9.158487e-21, -9.783621e-21, 
    5.90189e-20, 2.007333e-20, 3.172152e-22, 1.457137e-20, -5.258776e-21, 
    2.204792e-20, -1.059703e-20, -1.166094e-20, -1.532599e-20, -5.18582e-20, 
    1.755249e-20 ;

 M_SOIL2C_TO_LEACHING =
  3.744911e-20, 2.087486e-20, -1.060551e-20, 1.278678e-20, -2.114261e-21, 
    -1.111726e-20, 1.174379e-20, 1.931223e-20, -2.832878e-20, 2.39032e-20, 
    2.355656e-20, 7.602062e-21, -2.731745e-20, -1.994439e-20, -8.202881e-21, 
    -1.874136e-20, -1.340963e-20, -2.68368e-21, 8.491251e-21, -1.317101e-20, 
    1.7153e-20, 2.18545e-20, -3.301743e-21, 5.005454e-21, 8.139755e-23, 
    5.158974e-21, 2.444999e-20, 6.058045e-20, 2.873393e-20, 2.525068e-20, 
    1.209836e-20, -3.849803e-20, -1.209267e-20, -1.423408e-20, 4.493498e-20, 
    -2.027151e-20, 4.327751e-21, -1.577949e-20, -2.607851e-20, 2.663098e-20, 
    -1.536529e-20, -1.260119e-21, -2.162864e-20, 3.734166e-20, -1.139603e-20, 
    1.346166e-20, 8.146605e-21, 4.622676e-20, -7.837862e-21, 6.699318e-21, 
    -1.334801e-20, 2.750095e-20, 3.398876e-20, -2.079176e-20, -4.370163e-21, 
    3.03935e-21, -7.200026e-21, 4.100171e-21, -1.420469e-20, 3.381451e-21, 
    -9.766378e-21, 7.881126e-21, 4.600016e-22, -7.998454e-21, 1.622479e-20, 
    2.034259e-21, 2.239906e-20, 9.273581e-21, -4.936847e-20, 1.002706e-20, 
    5.179059e-21, 9.991418e-21, 3.775106e-20, 2.525775e-20, -1.122838e-20, 
    8.496044e-21, 3.044247e-20, 2.989907e-20, -1.357616e-20, -8.855698e-21, 
    -6.581815e-22, 7.511593e-21, -1.508143e-20, 8.468906e-21, 8.224917e-21, 
    -2.054236e-20, 2.201905e-21, -2.723913e-20, 2.714299e-20, 3.874542e-21, 
    -1.776623e-20, -3.054313e-20, 3.980564e-21, -1.046812e-20, -6.237038e-21, 
    1.223998e-20, 1.949597e-20, 1.228436e-20, 4.679875e-20, -1.649904e-20, 
    2.614922e-20, -4.17423e-21, 6.527966e-21, -2.946506e-20, 6.019615e-21, 
    5.257086e-21, 1.536811e-20, -2.460776e-20, 2.451729e-20, 2.674973e-20, 
    -1.970126e-20, 2.301991e-21, -3.560429e-21, 2.765984e-20, 5.389894e-20, 
    -1.243054e-20, -1.203444e-20, 9.35301e-21, -6.46946e-21, 6.675594e-21, 
    2.348759e-20, -6.31535e-21, 3.093584e-20, -3.024368e-21, 2.060457e-20, 
    6.533641e-21, -1.229934e-20, 3.537811e-20, 3.318526e-20, -3.571766e-20, 
    -7.544389e-21, -2.397047e-20, -1.203752e-20, -1.966533e-20, 
    -7.818913e-21, 3.613808e-20, 4.568336e-20, 2.626202e-20, 1.615382e-20, 
    2.627249e-20, 1.157244e-20, 2.561682e-20, 3.53419e-20, 2.846166e-20, 
    -3.109472e-20, 1.567658e-20, -8.749131e-21, -1.786746e-20, -2.995052e-20, 
    2.356589e-20, -1.411362e-20, 4.822822e-20, 8.018254e-21, 1.932147e-21, 
    -2.741639e-20, -1.223291e-20, -3.502891e-20, -8.714056e-21, 2.523062e-20, 
    1.435086e-20, 7.670478e-21, -3.890461e-20, -1.93588e-21, 1.338457e-21, 
    3.616664e-20, 1.286566e-20, -7.295859e-21, 1.666727e-20, -2.314461e-20, 
    -9.270729e-21, 2.266087e-20, -2.440984e-20, -2.492102e-20, 1.835769e-21, 
    -2.412684e-20, 7.409818e-21, -5.939523e-20, 1.583463e-20, 1.611906e-20, 
    9.613125e-21, 7.730723e-21, -1.167826e-22, -4.273873e-20, -7.750203e-21, 
    5.195184e-21, -2.550402e-20, -2.835704e-20, 7.649839e-21, -1.534494e-20, 
    4.279415e-20, -9.64223e-21, 1.391969e-20, 2.948881e-21, -2.72971e-20, 
    -3.133166e-20, -1.294058e-20, 2.099332e-20, 2.343858e-21, -5.89797e-22, 
    -1.347185e-20, 3.210098e-20, -1.228436e-20, 1.07774e-20, -2.716422e-20, 
    -4.341614e-21, 2.029328e-20, 1.046866e-20, -7.229667e-22, -6.79237e-24, 
    -2.621224e-20, -1.776371e-20, 4.078903e-20, 4.326633e-21, 1.772014e-20, 
    -4.198004e-21, -9.20994e-21, 8.703867e-21, 1.198381e-20, -3.153466e-20, 
    -4.117119e-21, -7.153236e-22, -7.611395e-20, -1.964272e-20, 
    -2.382018e-21, -1.898905e-20, -5.2636e-21, -6.282192e-22, 9.343965e-21, 
    2.021487e-22, -3.019282e-21, 1.402683e-20, 6.26078e-21, -3.87556e-20, 
    1.130074e-20, -1.215941e-20, -6.496859e-21, 3.492347e-20, -5.220615e-21, 
    2.203595e-21, 2.180024e-20, 1.407518e-20, -1.575654e-21, 9.184508e-21, 
    -6.194053e-21, -2.139396e-20, 5.042193e-20, 2.926293e-20, -9.728479e-21, 
    2.082795e-20, 8.65187e-21, 1.926237e-21, -8.806786e-21, -1.51032e-20, 
    -1.848324e-20, -3.782258e-20, 1.605918e-22, -1.668224e-20, 6.278235e-20, 
    1.040082e-20, 3.367127e-20, 1.645777e-21, -1.99805e-21, 2.740877e-20, 
    -1.212942e-20, -8.811579e-21, -3.726788e-20, 5.349719e-20, 2.052457e-20, 
    -4.32756e-20, -1.462839e-21, 7.838141e-21, -1.302822e-20, -1.592056e-20, 
    -1.785896e-20, 5.501958e-21, 3.968979e-21, -2.571944e-20, 1.086987e-20, 
    -3.241509e-20, 1.682333e-20, -3.140969e-20, 2.194541e-21, -3.34952e-21, 
    1.878633e-20, 1.072226e-20, -2.514888e-20, -6.282008e-21, -3.277443e-20, 
    -2.247258e-20, -2.386447e-20, -6.810985e-20, 3.228163e-20, -1.1657e-20, 
    3.771915e-20, 1.271158e-21, 2.470189e-20, -2.137332e-20, 1.067083e-20, 
    1.403137e-20, -2.679411e-20, -2.597956e-20, 3.000961e-20, 1.080454e-20, 
    3.223046e-20, -5.051549e-20, -5.618623e-20, -9.208543e-21, 3.6105e-20, 
    -5.212705e-21, 9.257171e-21, 9.222407e-21, 2.360377e-20, -2.126641e-20, 
    -9.911416e-21, -1.68174e-20, -1.879312e-20, 4.296802e-20, -4.249076e-20, 
    -1.529656e-20, -8.881423e-21, 1.701728e-20, -8.281765e-21, -1.132061e-21, 
    -4.539254e-21, -1.729067e-20, 4.156205e-22, 1.187895e-20, 1.762798e-20, 
    3.658706e-20, -3.197373e-20, 7.222088e-21, 5.645862e-21, 5.30572e-21, 
    -1.93942e-20, -2.441209e-20, 1.351623e-20, 3.330341e-20, -3.873186e-20 ;

 M_SOIL3C_TO_LEACHING =
  1.459825e-20, 1.816347e-20, 1.132451e-20, 2.037611e-20, 3.15714e-20, 
    -6.574932e-20, -2.88329e-20, 2.076431e-20, -4.51111e-20, 8.466671e-21, 
    2.439939e-20, 2.807709e-22, 2.746757e-20, -1.681118e-20, 1.047094e-20, 
    1.123544e-20, -1.058093e-20, 2.633693e-20, 1.386767e-20, 4.768802e-21, 
    1.279357e-20, 4.510291e-20, 1.586148e-20, 8.10108e-21, 8.032957e-21, 
    9.486196e-21, -6.994188e-21, 1.539725e-20, 1.522168e-20, -7.734942e-21, 
    -5.411297e-20, 1.654513e-20, 1.355524e-20, 1.028971e-20, 5.44511e-21, 
    2.382292e-20, -2.040131e-20, 2.977044e-20, -1.137032e-20, 1.597233e-20, 
    -7.486161e-21, 2.836723e-20, 8.56505e-21, 6.458153e-21, 1.022636e-20, 
    1.811033e-20, -7.739173e-21, 1.724089e-21, 3.739398e-21, 2.570729e-20, 
    1.509751e-22, -3.533905e-20, -1.233831e-21, -8.824591e-21, 7.314237e-21, 
    7.255992e-21, 1.939451e-20, 3.466026e-20, -8.61988e-21, 8.398783e-21, 
    -1.890819e-20, -1.393296e-20, -4.402414e-21, -2.229644e-20, 1.742493e-21, 
    2.086269e-20, -3.321691e-20, 2.827448e-20, 1.271452e-21, 1.158262e-20, 
    1.306499e-20, -1.252215e-20, -2.262582e-20, -1.571699e-20, 3.639875e-21, 
    -4.500396e-20, 1.161234e-20, 7.069969e-21, -5.372847e-20, 2.144204e-20, 
    1.591501e-21, 1.931164e-20, -1.504135e-21, 2.374654e-21, 1.652166e-20, 
    3.542418e-20, -5.948642e-21, -2.805001e-20, 2.829863e-21, 1.462086e-20, 
    1.771223e-20, 1.66257e-20, 2.947948e-20, 6.25202e-21, 6.467666e-20, 
    -4.112544e-20, 1.847354e-21, -2.916111e-21, 8.847745e-21, 1.453039e-20, 
    1.131124e-20, -7.084378e-21, -2.468608e-20, -3.541034e-20, -1.776171e-20, 
    1.415915e-20, 3.089371e-20, -4.200503e-20, 2.050561e-20, 5.346159e-21, 
    1.545887e-20, 2.070549e-20, 1.028264e-20, 1.869671e-20, -1.504214e-20, 
    -1.542777e-20, -1.628219e-20, 1.105818e-20, -4.565881e-22, -1.016191e-20, 
    -5.697336e-20, -2.15356e-20, -1.565226e-20, -2.979248e-20, 7.946163e-21, 
    1.510235e-20, 1.751431e-20, -9.967676e-21, -8.19212e-21, -6.127327e-21, 
    -1.724347e-20, -1.963791e-20, -1.940949e-20, 1.195216e-20, -2.389945e-21, 
    1.026848e-20, -5.885027e-21, 1.617899e-20, -2.148134e-20, -6.377563e-21, 
    1.381416e-21, -3.149591e-20, -2.408274e-21, -5.870918e-21, 3.453442e-20, 
    -6.930841e-21, 3.322513e-20, -1.694885e-20, -1.654033e-20, 1.120943e-20, 
    3.189655e-20, -2.480455e-20, -2.643647e-20, -1.664493e-20, 5.344191e-21, 
    6.88677e-21, 1.115598e-20, -3.332277e-21, -1.396747e-20, 8.612827e-21, 
    -5.875694e-21, -5.286796e-21, -2.793948e-20, -3.478041e-20, 2.120679e-20, 
    1.570739e-20, 1.713076e-21, 1.965885e-20, 6.361296e-22, -2.054549e-20, 
    -7.357793e-21, -2.501376e-20, 1.595874e-20, -4.950955e-20, -4.551571e-20, 
    -1.10265e-20, -1.777189e-20, -2.567082e-20, -3.221379e-20, 2.694143e-20, 
    -2.451335e-20, 1.016756e-20, -2.939581e-20, 2.448646e-20, -3.329947e-20, 
    1.84171e-20, -2.735815e-20, -1.50653e-20, -2.033687e-21, 2.665529e-20, 
    -1.480294e-20, 1.400337e-20, 4.545378e-20, 4.252072e-20, 1.008503e-21, 
    -1.404917e-20, 2.416211e-21, 3.134296e-20, 6.116003e-20, -1.711284e-20, 
    -2.006539e-20, -2.458684e-20, -5.667064e-21, 1.05976e-20, -1.090153e-20, 
    1.427676e-20, -9.064639e-21, -8.680126e-21, -1.647728e-20, -2.33711e-20, 
    3.365174e-20, -3.922098e-20, 2.795049e-20, 1.746171e-20, 8.902342e-21, 
    1.870234e-20, -5.959951e-22, -4.021859e-21, 3.2028e-20, 2.457723e-20, 
    2.992507e-20, -1.468872e-20, 7.921304e-21, 2.674266e-20, 1.67826e-20, 
    -8.213894e-21, -1.711907e-20, 1.092558e-20, 6.153069e-21, 2.236003e-20, 
    -4.602009e-20, 1.378427e-20, 1.738457e-20, 1.475488e-20, -8.661747e-21, 
    -3.230116e-20, -5.303859e-22, 1.667067e-20, -8.418304e-21, 2.094921e-20, 
    6.557676e-21, -7.130475e-21, 7.444301e-22, -1.231262e-20, -3.947484e-20, 
    1.771112e-20, 5.205634e-21, 9.319079e-21, -5.489555e-20, 1.240848e-20, 
    -1.989378e-20, -9.692286e-21, -3.61081e-20, 3.000254e-20, 2.730925e-20, 
    -1.206121e-21, 4.576507e-20, -6.606849e-21, -2.031392e-20, -2.272899e-20, 
    -1.372799e-20, 1.333273e-20, 1.226188e-21, 3.540637e-20, -1.003468e-20, 
    -3.65769e-21, 2.600283e-21, -3.263222e-20, -2.130093e-20, 2.053444e-21, 
    -2.431502e-21, -2.211972e-20, 1.941258e-20, 4.04898e-21, -1.094364e-20, 
    1.893752e-21, -5.429556e-21, 3.021544e-21, 2.308472e-21, -5.244929e-21, 
    9.386085e-21, -1.516312e-20, 2.85855e-20, 2.169025e-20, -7.835316e-21, 
    9.287999e-21, -1.961615e-20, -2.708758e-20, -5.220615e-21, 1.554058e-20, 
    -3.810067e-21, 6.705801e-21, 2.276971e-20, -6.649262e-21, 3.601698e-21, 
    4.321994e-20, 1.057808e-20, -1.021526e-21, -3.143033e-20, -1.239378e-20, 
    -3.967362e-20, 1.037368e-20, -2.255624e-20, 7.003504e-21, 6.918138e-21, 
    -1.190568e-21, -3.236984e-21, -7.498246e-20, 1.632629e-20, 1.752199e-20, 
    5.66424e-21, 1.015851e-21, -1.534152e-20, -1.276135e-20, -2.068288e-20, 
    4.067622e-20, -2.491705e-20, -2.428712e-20, -2.046772e-20, -5.528263e-20, 
    3.321069e-20, 3.382649e-20, 1.810523e-20, 1.813236e-20, -2.833804e-21, 
    -1.159987e-20, 9.167249e-21, -4.188573e-20, 2.058554e-22, -2.872997e-20, 
    9.09995e-21, 3.147527e-20, -9.574679e-21, 3.15979e-21, 2.644957e-21, 
    -7.046505e-21, 2.689338e-21, -3.624804e-20 ;

 NBP =
  -6.195836e-08, -6.223155e-08, -6.217844e-08, -6.23988e-08, -6.227657e-08, 
    -6.242085e-08, -6.201375e-08, -6.224239e-08, -6.209643e-08, 
    -6.198296e-08, -6.282642e-08, -6.240863e-08, -6.326049e-08, -6.2994e-08, 
    -6.366348e-08, -6.321901e-08, -6.375311e-08, -6.365067e-08, 
    -6.395901e-08, -6.387068e-08, -6.426506e-08, -6.399979e-08, 
    -6.446953e-08, -6.420172e-08, -6.424361e-08, -6.399104e-08, 
    -6.249272e-08, -6.27744e-08, -6.247603e-08, -6.251619e-08, -6.249817e-08, 
    -6.227909e-08, -6.216867e-08, -6.193749e-08, -6.197946e-08, 
    -6.214927e-08, -6.253426e-08, -6.240357e-08, -6.273295e-08, 
    -6.272551e-08, -6.309222e-08, -6.292688e-08, -6.354328e-08, 
    -6.336808e-08, -6.387437e-08, -6.374704e-08, -6.386838e-08, 
    -6.383159e-08, -6.386886e-08, -6.368212e-08, -6.376213e-08, 
    -6.359781e-08, -6.295784e-08, -6.314591e-08, -6.2585e-08, -6.224774e-08, 
    -6.202378e-08, -6.186485e-08, -6.188731e-08, -6.193014e-08, 
    -6.215026e-08, -6.235724e-08, -6.251497e-08, -6.262048e-08, 
    -6.272445e-08, -6.303911e-08, -6.32057e-08, -6.357869e-08, -6.351139e-08, 
    -6.362541e-08, -6.373437e-08, -6.391728e-08, -6.388717e-08, 
    -6.396776e-08, -6.362242e-08, -6.385192e-08, -6.347305e-08, 
    -6.357667e-08, -6.275266e-08, -6.243883e-08, -6.23054e-08, -6.218865e-08, 
    -6.190459e-08, -6.210075e-08, -6.202342e-08, -6.220741e-08, 
    -6.232432e-08, -6.22665e-08, -6.262336e-08, -6.248462e-08, -6.321557e-08, 
    -6.290072e-08, -6.372166e-08, -6.352521e-08, -6.376875e-08, 
    -6.364448e-08, -6.385741e-08, -6.366577e-08, -6.399775e-08, 
    -6.407004e-08, -6.402064e-08, -6.421042e-08, -6.365515e-08, 
    -6.386838e-08, -6.226487e-08, -6.22743e-08, -6.231824e-08, -6.212511e-08, 
    -6.21133e-08, -6.193633e-08, -6.20938e-08, -6.216086e-08, -6.23311e-08, 
    -6.243179e-08, -6.252751e-08, -6.273797e-08, -6.297304e-08, 
    -6.330175e-08, -6.353794e-08, -6.369626e-08, -6.359918e-08, 
    -6.368489e-08, -6.358908e-08, -6.354417e-08, -6.404295e-08, 
    -6.376287e-08, -6.418312e-08, -6.415987e-08, -6.396967e-08, 
    -6.416249e-08, -6.228093e-08, -6.222666e-08, -6.203825e-08, -6.21857e-08, 
    -6.191706e-08, -6.206743e-08, -6.215388e-08, -6.248751e-08, 
    -6.256082e-08, -6.262879e-08, -6.276304e-08, -6.293534e-08, 
    -6.323759e-08, -6.35006e-08, -6.374071e-08, -6.372311e-08, -6.372931e-08, 
    -6.378295e-08, -6.365008e-08, -6.380476e-08, -6.383071e-08, 
    -6.376284e-08, -6.415675e-08, -6.404422e-08, -6.415937e-08, -6.40861e-08, 
    -6.22443e-08, -6.233561e-08, -6.228627e-08, -6.237905e-08, -6.231368e-08, 
    -6.260434e-08, -6.269149e-08, -6.309931e-08, -6.293195e-08, 
    -6.319831e-08, -6.2959e-08, -6.300141e-08, -6.320698e-08, -6.297194e-08, 
    -6.348608e-08, -6.313749e-08, -6.378503e-08, -6.343689e-08, 
    -6.380684e-08, -6.373967e-08, -6.38509e-08, -6.395051e-08, -6.407584e-08, 
    -6.430709e-08, -6.425354e-08, -6.444694e-08, -6.247174e-08, 
    -6.259017e-08, -6.257976e-08, -6.270371e-08, -6.279537e-08, 
    -6.299408e-08, -6.331277e-08, -6.319293e-08, -6.341295e-08, 
    -6.345712e-08, -6.312285e-08, -6.332808e-08, -6.266944e-08, 
    -6.277585e-08, -6.27125e-08, -6.248108e-08, -6.322053e-08, -6.284102e-08, 
    -6.354184e-08, -6.333624e-08, -6.393631e-08, -6.363786e-08, 
    -6.422406e-08, -6.447465e-08, -6.471054e-08, -6.498618e-08, 
    -6.265482e-08, -6.257435e-08, -6.271845e-08, -6.291781e-08, 
    -6.310282e-08, -6.334877e-08, -6.337395e-08, -6.342002e-08, 
    -6.353938e-08, -6.363974e-08, -6.343458e-08, -6.36649e-08, -6.28005e-08, 
    -6.325348e-08, -6.254392e-08, -6.275756e-08, -6.290607e-08, 
    -6.284093e-08, -6.317924e-08, -6.325897e-08, -6.358299e-08, 
    -6.341549e-08, -6.44128e-08, -6.397154e-08, -6.519609e-08, -6.485385e-08, 
    -6.254623e-08, -6.265455e-08, -6.303155e-08, -6.285217e-08, -6.33652e-08, 
    -6.349148e-08, -6.359415e-08, -6.372539e-08, -6.373956e-08, 
    -6.381732e-08, -6.36899e-08, -6.381229e-08, -6.33493e-08, -6.355619e-08, 
    -6.298847e-08, -6.312663e-08, -6.306308e-08, -6.299335e-08, 
    -6.320855e-08, -6.343781e-08, -6.344272e-08, -6.351623e-08, 
    -6.372337e-08, -6.336728e-08, -6.446972e-08, -6.378883e-08, 
    -6.277267e-08, -6.298131e-08, -6.301112e-08, -6.29303e-08, -6.347882e-08, 
    -6.328006e-08, -6.381542e-08, -6.367073e-08, -6.390781e-08, -6.379e-08, 
    -6.377267e-08, -6.362136e-08, -6.352716e-08, -6.328918e-08, 
    -6.309555e-08, -6.294202e-08, -6.297773e-08, -6.314637e-08, 
    -6.345184e-08, -6.374083e-08, -6.367753e-08, -6.388979e-08, -6.3328e-08, 
    -6.356355e-08, -6.347251e-08, -6.370992e-08, -6.318974e-08, 
    -6.363265e-08, -6.307653e-08, -6.312529e-08, -6.327612e-08, 
    -6.357952e-08, -6.364667e-08, -6.371835e-08, -6.367412e-08, 
    -6.345959e-08, -6.342446e-08, -6.327246e-08, -6.323049e-08, 
    -6.311468e-08, -6.301879e-08, -6.310639e-08, -6.319839e-08, 
    -6.345969e-08, -6.369518e-08, -6.395192e-08, -6.401477e-08, 
    -6.431474e-08, -6.407053e-08, -6.447351e-08, -6.413087e-08, 
    -6.472403e-08, -6.365835e-08, -6.412082e-08, -6.328299e-08, 
    -6.337325e-08, -6.353649e-08, -6.391095e-08, -6.37088e-08, -6.394522e-08, 
    -6.342308e-08, -6.315219e-08, -6.308211e-08, -6.295136e-08, -6.30851e-08, 
    -6.307422e-08, -6.320221e-08, -6.316108e-08, -6.346837e-08, -6.33033e-08, 
    -6.377223e-08, -6.394335e-08, -6.442666e-08, -6.472296e-08, 
    -6.502461e-08, -6.515778e-08, -6.519831e-08, -6.521526e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.195836e-08, -6.223155e-08, -6.217844e-08, -6.23988e-08, -6.227657e-08, 
    -6.242085e-08, -6.201375e-08, -6.224239e-08, -6.209643e-08, 
    -6.198296e-08, -6.282642e-08, -6.240863e-08, -6.326049e-08, -6.2994e-08, 
    -6.366348e-08, -6.321901e-08, -6.375311e-08, -6.365067e-08, 
    -6.395901e-08, -6.387068e-08, -6.426506e-08, -6.399979e-08, 
    -6.446953e-08, -6.420172e-08, -6.424361e-08, -6.399104e-08, 
    -6.249272e-08, -6.27744e-08, -6.247603e-08, -6.251619e-08, -6.249817e-08, 
    -6.227909e-08, -6.216867e-08, -6.193749e-08, -6.197946e-08, 
    -6.214927e-08, -6.253426e-08, -6.240357e-08, -6.273295e-08, 
    -6.272551e-08, -6.309222e-08, -6.292688e-08, -6.354328e-08, 
    -6.336808e-08, -6.387437e-08, -6.374704e-08, -6.386838e-08, 
    -6.383159e-08, -6.386886e-08, -6.368212e-08, -6.376213e-08, 
    -6.359781e-08, -6.295784e-08, -6.314591e-08, -6.2585e-08, -6.224774e-08, 
    -6.202378e-08, -6.186485e-08, -6.188731e-08, -6.193014e-08, 
    -6.215026e-08, -6.235724e-08, -6.251497e-08, -6.262048e-08, 
    -6.272445e-08, -6.303911e-08, -6.32057e-08, -6.357869e-08, -6.351139e-08, 
    -6.362541e-08, -6.373437e-08, -6.391728e-08, -6.388717e-08, 
    -6.396776e-08, -6.362242e-08, -6.385192e-08, -6.347305e-08, 
    -6.357667e-08, -6.275266e-08, -6.243883e-08, -6.23054e-08, -6.218865e-08, 
    -6.190459e-08, -6.210075e-08, -6.202342e-08, -6.220741e-08, 
    -6.232432e-08, -6.22665e-08, -6.262336e-08, -6.248462e-08, -6.321557e-08, 
    -6.290072e-08, -6.372166e-08, -6.352521e-08, -6.376875e-08, 
    -6.364448e-08, -6.385741e-08, -6.366577e-08, -6.399775e-08, 
    -6.407004e-08, -6.402064e-08, -6.421042e-08, -6.365515e-08, 
    -6.386838e-08, -6.226487e-08, -6.22743e-08, -6.231824e-08, -6.212511e-08, 
    -6.21133e-08, -6.193633e-08, -6.20938e-08, -6.216086e-08, -6.23311e-08, 
    -6.243179e-08, -6.252751e-08, -6.273797e-08, -6.297304e-08, 
    -6.330175e-08, -6.353794e-08, -6.369626e-08, -6.359918e-08, 
    -6.368489e-08, -6.358908e-08, -6.354417e-08, -6.404295e-08, 
    -6.376287e-08, -6.418312e-08, -6.415987e-08, -6.396967e-08, 
    -6.416249e-08, -6.228093e-08, -6.222666e-08, -6.203825e-08, -6.21857e-08, 
    -6.191706e-08, -6.206743e-08, -6.215388e-08, -6.248751e-08, 
    -6.256082e-08, -6.262879e-08, -6.276304e-08, -6.293534e-08, 
    -6.323759e-08, -6.35006e-08, -6.374071e-08, -6.372311e-08, -6.372931e-08, 
    -6.378295e-08, -6.365008e-08, -6.380476e-08, -6.383071e-08, 
    -6.376284e-08, -6.415675e-08, -6.404422e-08, -6.415937e-08, -6.40861e-08, 
    -6.22443e-08, -6.233561e-08, -6.228627e-08, -6.237905e-08, -6.231368e-08, 
    -6.260434e-08, -6.269149e-08, -6.309931e-08, -6.293195e-08, 
    -6.319831e-08, -6.2959e-08, -6.300141e-08, -6.320698e-08, -6.297194e-08, 
    -6.348608e-08, -6.313749e-08, -6.378503e-08, -6.343689e-08, 
    -6.380684e-08, -6.373967e-08, -6.38509e-08, -6.395051e-08, -6.407584e-08, 
    -6.430709e-08, -6.425354e-08, -6.444694e-08, -6.247174e-08, 
    -6.259017e-08, -6.257976e-08, -6.270371e-08, -6.279537e-08, 
    -6.299408e-08, -6.331277e-08, -6.319293e-08, -6.341295e-08, 
    -6.345712e-08, -6.312285e-08, -6.332808e-08, -6.266944e-08, 
    -6.277585e-08, -6.27125e-08, -6.248108e-08, -6.322053e-08, -6.284102e-08, 
    -6.354184e-08, -6.333624e-08, -6.393631e-08, -6.363786e-08, 
    -6.422406e-08, -6.447465e-08, -6.471054e-08, -6.498618e-08, 
    -6.265482e-08, -6.257435e-08, -6.271845e-08, -6.291781e-08, 
    -6.310282e-08, -6.334877e-08, -6.337395e-08, -6.342002e-08, 
    -6.353938e-08, -6.363974e-08, -6.343458e-08, -6.36649e-08, -6.28005e-08, 
    -6.325348e-08, -6.254392e-08, -6.275756e-08, -6.290607e-08, 
    -6.284093e-08, -6.317924e-08, -6.325897e-08, -6.358299e-08, 
    -6.341549e-08, -6.44128e-08, -6.397154e-08, -6.519609e-08, -6.485385e-08, 
    -6.254623e-08, -6.265455e-08, -6.303155e-08, -6.285217e-08, -6.33652e-08, 
    -6.349148e-08, -6.359415e-08, -6.372539e-08, -6.373956e-08, 
    -6.381732e-08, -6.36899e-08, -6.381229e-08, -6.33493e-08, -6.355619e-08, 
    -6.298847e-08, -6.312663e-08, -6.306308e-08, -6.299335e-08, 
    -6.320855e-08, -6.343781e-08, -6.344272e-08, -6.351623e-08, 
    -6.372337e-08, -6.336728e-08, -6.446972e-08, -6.378883e-08, 
    -6.277267e-08, -6.298131e-08, -6.301112e-08, -6.29303e-08, -6.347882e-08, 
    -6.328006e-08, -6.381542e-08, -6.367073e-08, -6.390781e-08, -6.379e-08, 
    -6.377267e-08, -6.362136e-08, -6.352716e-08, -6.328918e-08, 
    -6.309555e-08, -6.294202e-08, -6.297773e-08, -6.314637e-08, 
    -6.345184e-08, -6.374083e-08, -6.367753e-08, -6.388979e-08, -6.3328e-08, 
    -6.356355e-08, -6.347251e-08, -6.370992e-08, -6.318974e-08, 
    -6.363265e-08, -6.307653e-08, -6.312529e-08, -6.327612e-08, 
    -6.357952e-08, -6.364667e-08, -6.371835e-08, -6.367412e-08, 
    -6.345959e-08, -6.342446e-08, -6.327246e-08, -6.323049e-08, 
    -6.311468e-08, -6.301879e-08, -6.310639e-08, -6.319839e-08, 
    -6.345969e-08, -6.369518e-08, -6.395192e-08, -6.401477e-08, 
    -6.431474e-08, -6.407053e-08, -6.447351e-08, -6.413087e-08, 
    -6.472403e-08, -6.365835e-08, -6.412082e-08, -6.328299e-08, 
    -6.337325e-08, -6.353649e-08, -6.391095e-08, -6.37088e-08, -6.394522e-08, 
    -6.342308e-08, -6.315219e-08, -6.308211e-08, -6.295136e-08, -6.30851e-08, 
    -6.307422e-08, -6.320221e-08, -6.316108e-08, -6.346837e-08, -6.33033e-08, 
    -6.377223e-08, -6.394335e-08, -6.442666e-08, -6.472296e-08, 
    -6.502461e-08, -6.515778e-08, -6.519831e-08, -6.521526e-08 ;

 NET_NMIN =
  8.728431e-09, 8.766915e-09, 8.759435e-09, 8.790474e-09, 8.773257e-09, 
    8.793581e-09, 8.736235e-09, 8.768443e-09, 8.747882e-09, 8.731897e-09, 
    8.850712e-09, 8.79186e-09, 8.911858e-09, 8.874319e-09, 8.968625e-09, 
    8.906015e-09, 8.98125e-09, 8.966821e-09, 9.010256e-09, 8.997812e-09, 
    9.053367e-09, 9.016e-09, 9.08217e-09, 9.044444e-09, 9.050344e-09, 
    9.014766e-09, 8.803704e-09, 8.843384e-09, 8.801353e-09, 8.807011e-09, 
    8.804473e-09, 8.773611e-09, 8.758058e-09, 8.725491e-09, 8.731404e-09, 
    8.755324e-09, 8.809556e-09, 8.791147e-09, 8.837546e-09, 8.836498e-09, 
    8.888154e-09, 8.864864e-09, 8.951692e-09, 8.927014e-09, 8.998332e-09, 
    8.980395e-09, 8.997489e-09, 8.992306e-09, 8.997556e-09, 8.97125e-09, 
    8.982521e-09, 8.959375e-09, 8.869224e-09, 8.895717e-09, 8.816705e-09, 
    8.769196e-09, 8.737647e-09, 8.715258e-09, 8.718423e-09, 8.724457e-09, 
    8.755464e-09, 8.78462e-09, 8.80684e-09, 8.821702e-09, 8.836348e-09, 
    8.880673e-09, 8.90414e-09, 8.956682e-09, 8.947201e-09, 8.963263e-09, 
    8.978611e-09, 9.004377e-09, 9.000136e-09, 9.011488e-09, 8.962841e-09, 
    8.995171e-09, 8.9418e-09, 8.956397e-09, 8.840322e-09, 8.796114e-09, 
    8.777318e-09, 8.760872e-09, 8.720857e-09, 8.74849e-09, 8.737596e-09, 
    8.763514e-09, 8.779983e-09, 8.771838e-09, 8.822108e-09, 8.802564e-09, 
    8.905531e-09, 8.861178e-09, 8.976821e-09, 8.949147e-09, 8.983454e-09, 
    8.965948e-09, 8.995944e-09, 8.968948e-09, 9.015713e-09, 9.025895e-09, 
    9.018937e-09, 9.045669e-09, 8.967452e-09, 8.997488e-09, 8.771609e-09, 
    8.772938e-09, 8.779127e-09, 8.751922e-09, 8.750257e-09, 8.725329e-09, 
    8.747511e-09, 8.756957e-09, 8.780938e-09, 8.795122e-09, 8.808606e-09, 
    8.838254e-09, 8.871366e-09, 8.917671e-09, 8.95094e-09, 8.973243e-09, 
    8.959568e-09, 8.97164e-09, 8.958144e-09, 8.951819e-09, 9.022079e-09, 
    8.982626e-09, 9.041824e-09, 9.038549e-09, 9.011757e-09, 9.038918e-09, 
    8.773871e-09, 8.766227e-09, 8.739685e-09, 8.760456e-09, 8.722615e-09, 
    8.743796e-09, 8.755975e-09, 8.802971e-09, 8.813299e-09, 8.822873e-09, 
    8.841785e-09, 8.866055e-09, 8.908632e-09, 8.945681e-09, 8.979504e-09, 
    8.977026e-09, 8.977898e-09, 8.985453e-09, 8.966738e-09, 8.988526e-09, 
    8.992183e-09, 8.982622e-09, 9.03811e-09, 9.022258e-09, 9.038479e-09, 
    9.028158e-09, 8.768712e-09, 8.781574e-09, 8.774624e-09, 8.787693e-09, 
    8.778485e-09, 8.819429e-09, 8.831705e-09, 8.889153e-09, 8.865577e-09, 
    8.9031e-09, 8.869389e-09, 8.875362e-09, 8.904321e-09, 8.871211e-09, 
    8.943637e-09, 8.894531e-09, 8.985747e-09, 8.936706e-09, 8.98882e-09, 
    8.979358e-09, 8.995026e-09, 9.009058e-09, 9.026713e-09, 9.059287e-09, 
    9.051743e-09, 9.078986e-09, 8.80075e-09, 8.817433e-09, 8.815966e-09, 
    8.833426e-09, 8.846339e-09, 8.874329e-09, 8.919223e-09, 8.902341e-09, 
    8.933335e-09, 8.939557e-09, 8.89247e-09, 8.921379e-09, 8.8286e-09, 
    8.843588e-09, 8.834665e-09, 8.802066e-09, 8.90623e-09, 8.85277e-09, 
    8.95149e-09, 8.922528e-09, 9.007056e-09, 8.965017e-09, 9.047591e-09, 
    9.08289e-09, 9.116119e-09, 9.154946e-09, 8.82654e-09, 8.815204e-09, 
    8.835503e-09, 8.863586e-09, 8.889648e-09, 8.924294e-09, 8.92784e-09, 
    8.934331e-09, 8.951145e-09, 8.965281e-09, 8.936381e-09, 8.968825e-09, 
    8.847062e-09, 8.91087e-09, 8.810917e-09, 8.841012e-09, 8.861932e-09, 
    8.852756e-09, 8.900412e-09, 8.911644e-09, 8.957287e-09, 8.933693e-09, 
    9.074177e-09, 9.01202e-09, 9.184515e-09, 9.136306e-09, 8.811242e-09, 
    8.826501e-09, 8.879608e-09, 8.854339e-09, 8.926608e-09, 8.944397e-09, 
    8.958859e-09, 8.977345e-09, 8.979342e-09, 8.990296e-09, 8.972346e-09, 
    8.989587e-09, 8.924368e-09, 8.953513e-09, 8.873539e-09, 8.893003e-09, 
    8.884049e-09, 8.874227e-09, 8.904541e-09, 8.936836e-09, 8.937528e-09, 
    8.947883e-09, 8.977062e-09, 8.926901e-09, 9.082195e-09, 8.986284e-09, 
    8.84314e-09, 8.87253e-09, 8.87673e-09, 8.865346e-09, 8.942614e-09, 
    8.914616e-09, 8.990028e-09, 8.969647e-09, 9.003043e-09, 8.986447e-09, 
    8.984006e-09, 8.962693e-09, 8.949423e-09, 8.915899e-09, 8.888623e-09, 
    8.866997e-09, 8.872026e-09, 8.895783e-09, 8.938812e-09, 8.979522e-09, 
    8.970604e-09, 9.000504e-09, 8.921368e-09, 8.954549e-09, 8.941724e-09, 
    8.975166e-09, 8.901892e-09, 8.964284e-09, 8.885944e-09, 8.892813e-09, 
    8.91406e-09, 8.956799e-09, 8.966258e-09, 8.976354e-09, 8.970124e-09, 
    8.939905e-09, 8.934955e-09, 8.913544e-09, 8.907631e-09, 8.891318e-09, 
    8.87781e-09, 8.890151e-09, 8.90311e-09, 8.939918e-09, 8.97309e-09, 
    9.009257e-09, 9.018109e-09, 9.060365e-09, 9.025964e-09, 9.08273e-09, 
    9.034465e-09, 9.118018e-09, 8.967902e-09, 9.033048e-09, 8.915027e-09, 
    8.927741e-09, 8.950737e-09, 9.003484e-09, 8.97501e-09, 9.008311e-09, 
    8.934761e-09, 8.896602e-09, 8.88673e-09, 8.868311e-09, 8.887151e-09, 
    8.885619e-09, 8.903648e-09, 8.897855e-09, 8.94114e-09, 8.91789e-09, 
    8.983944e-09, 9.008049e-09, 9.076131e-09, 9.117868e-09, 9.16036e-09, 
    9.179119e-09, 9.184828e-09, 9.187215e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14 ;

 O_SCALAR =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5 ;

 PCH4 =
  0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627 ;

 PCO2 =
  28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  5.044949e-14, 5.058576e-14, 5.055929e-14, 5.066909e-14, 5.060821e-14, 
    5.068008e-14, 5.047715e-14, 5.059115e-14, 5.051839e-14, 5.046179e-14, 
    5.088186e-14, 5.067399e-14, 5.109757e-14, 5.096525e-14, 5.129742e-14, 
    5.107696e-14, 5.134183e-14, 5.129111e-14, 5.144381e-14, 5.140008e-14, 
    5.159509e-14, 5.146398e-14, 5.169611e-14, 5.156382e-14, 5.158451e-14, 
    5.145965e-14, 5.071589e-14, 5.085598e-14, 5.070758e-14, 5.072757e-14, 
    5.07186e-14, 5.060945e-14, 5.055439e-14, 5.04391e-14, 5.046004e-14, 
    5.054473e-14, 5.073656e-14, 5.06715e-14, 5.083547e-14, 5.083177e-14, 
    5.101405e-14, 5.093189e-14, 5.123788e-14, 5.1151e-14, 5.140191e-14, 
    5.133885e-14, 5.139894e-14, 5.138073e-14, 5.139918e-14, 5.130669e-14, 
    5.134632e-14, 5.126492e-14, 5.094728e-14, 5.10407e-14, 5.076183e-14, 
    5.059379e-14, 5.048214e-14, 5.040283e-14, 5.041405e-14, 5.043541e-14, 
    5.054522e-14, 5.064841e-14, 5.072698e-14, 5.07795e-14, 5.083124e-14, 
    5.09876e-14, 5.107037e-14, 5.125542e-14, 5.122208e-14, 5.127858e-14, 
    5.133258e-14, 5.142314e-14, 5.140825e-14, 5.144812e-14, 5.127711e-14, 
    5.139078e-14, 5.120307e-14, 5.125444e-14, 5.084517e-14, 5.068906e-14, 
    5.062253e-14, 5.056437e-14, 5.042267e-14, 5.052053e-14, 5.048196e-14, 
    5.057374e-14, 5.063201e-14, 5.06032e-14, 5.078094e-14, 5.071186e-14, 
    5.107527e-14, 5.091887e-14, 5.132628e-14, 5.122893e-14, 5.134961e-14, 
    5.128805e-14, 5.13935e-14, 5.12986e-14, 5.146297e-14, 5.149871e-14, 
    5.147428e-14, 5.156814e-14, 5.129333e-14, 5.139893e-14, 5.060239e-14, 
    5.060708e-14, 5.062899e-14, 5.053268e-14, 5.05268e-14, 5.043851e-14, 
    5.051708e-14, 5.055051e-14, 5.06354e-14, 5.068555e-14, 5.073322e-14, 
    5.083796e-14, 5.095482e-14, 5.111807e-14, 5.123524e-14, 5.131371e-14, 
    5.126561e-14, 5.130807e-14, 5.126059e-14, 5.123834e-14, 5.148531e-14, 
    5.134668e-14, 5.155464e-14, 5.154315e-14, 5.144906e-14, 5.154445e-14, 
    5.061038e-14, 5.058334e-14, 5.048937e-14, 5.056292e-14, 5.04289e-14, 
    5.050392e-14, 5.054702e-14, 5.071328e-14, 5.074981e-14, 5.078363e-14, 
    5.085044e-14, 5.09361e-14, 5.108622e-14, 5.121671e-14, 5.133573e-14, 
    5.132702e-14, 5.133008e-14, 5.135664e-14, 5.129082e-14, 5.136744e-14, 
    5.138028e-14, 5.134668e-14, 5.154161e-14, 5.148596e-14, 5.154291e-14, 
    5.150668e-14, 5.059214e-14, 5.063764e-14, 5.061305e-14, 5.065928e-14, 
    5.06267e-14, 5.077144e-14, 5.08148e-14, 5.101754e-14, 5.093441e-14, 
    5.106672e-14, 5.094787e-14, 5.096893e-14, 5.107098e-14, 5.09543e-14, 
    5.120949e-14, 5.103649e-14, 5.135767e-14, 5.118507e-14, 5.136848e-14, 
    5.133521e-14, 5.139029e-14, 5.143959e-14, 5.15016e-14, 5.161589e-14, 
    5.158944e-14, 5.168497e-14, 5.070545e-14, 5.07644e-14, 5.075924e-14, 
    5.082092e-14, 5.086651e-14, 5.09653e-14, 5.112355e-14, 5.106407e-14, 
    5.117327e-14, 5.119517e-14, 5.102928e-14, 5.113113e-14, 5.080386e-14, 
    5.085677e-14, 5.082528e-14, 5.071009e-14, 5.107774e-14, 5.088918e-14, 
    5.123717e-14, 5.11352e-14, 5.143256e-14, 5.128474e-14, 5.157487e-14, 
    5.169861e-14, 5.181506e-14, 5.195085e-14, 5.079659e-14, 5.075655e-14, 
    5.082826e-14, 5.092736e-14, 5.101932e-14, 5.114141e-14, 5.115391e-14, 
    5.117676e-14, 5.123596e-14, 5.12857e-14, 5.118396e-14, 5.129817e-14, 
    5.086898e-14, 5.109411e-14, 5.074138e-14, 5.084767e-14, 5.092153e-14, 
    5.088916e-14, 5.105728e-14, 5.109686e-14, 5.125756e-14, 5.117453e-14, 
    5.166806e-14, 5.144996e-14, 5.205423e-14, 5.188567e-14, 5.074255e-14, 
    5.079646e-14, 5.09839e-14, 5.089475e-14, 5.114957e-14, 5.12122e-14, 
    5.126311e-14, 5.132812e-14, 5.133515e-14, 5.137365e-14, 5.131056e-14, 
    5.137117e-14, 5.114167e-14, 5.124429e-14, 5.096252e-14, 5.103114e-14, 
    5.099959e-14, 5.096494e-14, 5.107183e-14, 5.118556e-14, 5.118803e-14, 
    5.122447e-14, 5.132701e-14, 5.115061e-14, 5.16961e-14, 5.135945e-14, 
    5.085523e-14, 5.095891e-14, 5.097376e-14, 5.093361e-14, 5.120592e-14, 
    5.110732e-14, 5.137272e-14, 5.130106e-14, 5.141846e-14, 5.136013e-14, 
    5.135155e-14, 5.12766e-14, 5.122989e-14, 5.111183e-14, 5.10157e-14, 
    5.093944e-14, 5.095718e-14, 5.104094e-14, 5.119252e-14, 5.133577e-14, 
    5.13044e-14, 5.140955e-14, 5.113111e-14, 5.124792e-14, 5.120278e-14, 
    5.132047e-14, 5.106248e-14, 5.128208e-14, 5.100627e-14, 5.103049e-14, 
    5.110536e-14, 5.125581e-14, 5.128914e-14, 5.132463e-14, 5.130274e-14, 
    5.119638e-14, 5.117896e-14, 5.110355e-14, 5.10827e-14, 5.102522e-14, 
    5.097758e-14, 5.102109e-14, 5.106677e-14, 5.119644e-14, 5.131315e-14, 
    5.144028e-14, 5.147139e-14, 5.161961e-14, 5.149891e-14, 5.169796e-14, 
    5.152867e-14, 5.182161e-14, 5.129486e-14, 5.152377e-14, 5.110878e-14, 
    5.115357e-14, 5.123449e-14, 5.141997e-14, 5.131992e-14, 5.143694e-14, 
    5.117828e-14, 5.104381e-14, 5.100904e-14, 5.094406e-14, 5.101053e-14, 
    5.100512e-14, 5.106868e-14, 5.104827e-14, 5.120074e-14, 5.111886e-14, 
    5.135132e-14, 5.143602e-14, 5.167495e-14, 5.182114e-14, 5.196983e-14, 
    5.203539e-14, 5.205534e-14, 5.206367e-14 ;

 POT_F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.904545e-44, 0, 3.640714e-41, 
    2.382207e-44, 1.485699e-40, 2.970192e-41, 3.462017e-39, 9.090784e-40, 
    3.043702e-37, 6.372947e-39, 5.297037e-36, 1.228662e-37, 2.240759e-37, 
    5.592868e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 
    5.327737e-42, 3.012792e-43, 9.616453e-40, 1.350768e-40, 8.778827e-40, 
    4.997395e-40, 8.843286e-40, 4.883105e-41, 1.708729e-40, 1.279946e-41, 0, 
    7.006492e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    1.961818e-44, 9.427936e-42, 3.179546e-42, 1.989283e-41, 1.108483e-40, 
    1.845646e-39, 1.168838e-39, 3.948533e-39, 1.895536e-41, 6.828597e-40, 
    1.702578e-42, 9.121052e-42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.242078e-44, 0, 9.087421e-41, 3.976885e-42, 1.893603e-40, 2.691614e-41, 
    7.425691e-40, 3.771455e-41, 6.183549e-39, 1.806158e-38, 8.695494e-39, 
    1.391768e-37, 3.187954e-41, 8.78027e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9.949219e-44, 4.887729e-42, 6.099011e-41, 1.308112e-41, 
    5.099465e-41, 1.112771e-41, 5.404808e-42, 1.210799e-38, 1.728852e-40, 
    9.393621e-38, 6.709526e-38, 4.063952e-39, 6.969254e-38, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3.363116e-44, 2.668072e-42, 1.22367e-40, 9.295093e-41, 
    1.024097e-40, 2.360095e-40, 2.942166e-41, 3.306658e-40, 4.932346e-40, 
    1.727591e-40, 6.41323e-38, 1.233066e-38, 6.661603e-38, 2.286338e-38, 0, 
    0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 1.681558e-44, 0, 0, 1.961818e-44, 0, 
    2.107553e-42, 5.605194e-45, 2.437545e-40, 9.416726e-43, 3.41488e-40, 
    1.20401e-40, 6.718792e-40, 3.047178e-39, 1.966447e-38, 5.518767e-37, 
    2.580681e-37, 3.881303e-36, 0, 0, 0, 0, 0, 0, 1.191104e-43, 1.541428e-44, 
    6.347882e-43, 1.311615e-42, 4.203895e-45, 1.541428e-43, 0, 0, 0, 0, 
    2.522337e-44, 0, 5.205824e-42, 1.765636e-43, 2.460338e-39, 2.425227e-41, 
    1.693173e-37, 5.68547e-36, 1.346246e-34, 4.604947e-33, 0, 0, 0, 0, 
    2.802597e-45, 2.186026e-43, 3.321077e-43, 7.132609e-43, 5.002636e-42, 
    2.496693e-41, 9.066401e-43, 3.719607e-41, 0, 4.344025e-44, 0, 0, 0, 0, 
    1.261169e-44, 4.764415e-44, 1.009916e-41, 6.614129e-43, 2.424143e-36, 
    4.18154e-39, 6.026268e-32, 8.63849e-34, 0, 0, 1.401298e-45, 0, 
    2.872662e-43, 2.299531e-42, 1.206938e-41, 9.634768e-41, 1.20202e-40, 
    4.013333e-40, 5.518173e-41, 3.713385e-40, 2.200039e-43, 6.562281e-42, 0, 
    5.605194e-45, 1.401298e-45, 0, 2.101948e-44, 9.556856e-43, 1.03556e-42, 
    3.440188e-42, 9.359973e-41, 2.970753e-43, 5.321813e-36, 2.591547e-40, 0, 
    0, 0, 0, 1.870733e-42, 6.866362e-44, 3.897558e-40, 4.0789e-41, 
    1.598796e-39, 2.632255e-40, 2.012363e-40, 1.863867e-41, 4.105805e-42, 
    7.987401e-44, 2.802597e-45, 0, 0, 7.006492e-45, 1.203715e-42, 
    1.226613e-40, 4.54329e-41, 1.216202e-39, 1.541428e-43, 7.390448e-42, 
    1.688565e-42, 7.559725e-41, 1.541428e-44, 2.236612e-41, 1.401298e-45, 
    4.203895e-45, 6.445973e-44, 9.556856e-42, 2.787043e-41, 8.629336e-41, 
    4.303107e-41, 1.366266e-42, 7.665103e-43, 6.025583e-44, 2.942727e-44, 
    4.203895e-45, 1.401298e-45, 4.203895e-45, 1.681558e-44, 1.367667e-42, 
    5.998398e-41, 3.113122e-39, 7.966207e-39, 6.155813e-37, 1.82089e-38, 
    5.606511e-36, 4.415561e-38, 1.609795e-34, 3.358352e-41, 3.807932e-38, 
    7.286752e-44, 3.279038e-43, 4.778428e-42, 1.678356e-39, 7.428563e-41, 
    2.815552e-39, 7.496947e-43, 8.407791e-45, 2.802597e-45, 0, 2.802597e-45, 
    1.401298e-45, 1.821688e-44, 8.407791e-45, 1.576461e-42, 1.022948e-43, 
    1.99912e-40, 2.737107e-39, 2.934797e-36, 1.585659e-34, 7.423095e-33, 
    3.795473e-32, 6.187504e-32, 7.582037e-32 ;

 POT_F_NIT =
  3.837638e-11, 3.870687e-11, 3.864251e-11, 3.890991e-11, 3.876146e-11, 
    3.893671e-11, 3.844325e-11, 3.871999e-11, 3.85432e-11, 3.840604e-11, 
    3.943156e-11, 3.892183e-11, 3.996478e-11, 3.963697e-11, 4.046314e-11, 
    3.991366e-11, 4.057441e-11, 4.044724e-11, 4.083065e-11, 4.072061e-11, 
    4.121304e-11, 4.088148e-11, 4.146955e-11, 4.113373e-11, 4.118616e-11, 
    4.087053e-11, 3.902418e-11, 3.936794e-11, 3.900385e-11, 3.905276e-11, 
    3.903081e-11, 3.87645e-11, 3.863064e-11, 3.835115e-11, 3.84018e-11, 
    3.860712e-11, 3.907473e-11, 3.891567e-11, 3.93172e-11, 3.930811e-11, 
    3.97576e-11, 3.95546e-11, 4.031413e-11, 4.009748e-11, 4.072519e-11, 
    4.056684e-11, 4.071773e-11, 4.067194e-11, 4.071832e-11, 4.048622e-11, 
    4.058556e-11, 4.038165e-11, 3.959263e-11, 3.982369e-11, 3.913661e-11, 
    3.872647e-11, 3.845534e-11, 3.826354e-11, 3.829061e-11, 3.834227e-11, 
    3.860832e-11, 3.885935e-11, 3.905122e-11, 3.917984e-11, 3.930679e-11, 
    3.969234e-11, 3.989723e-11, 4.035799e-11, 4.027464e-11, 4.041589e-11, 
    4.05511e-11, 4.077861e-11, 4.074111e-11, 4.08415e-11, 4.041215e-11, 
    4.069722e-11, 4.022717e-11, 4.035544e-11, 3.934133e-11, 3.895857e-11, 
    3.879643e-11, 3.865483e-11, 3.831144e-11, 3.85484e-11, 3.845489e-11, 
    3.867754e-11, 3.881936e-11, 3.874918e-11, 3.918335e-11, 3.901425e-11, 
    3.990938e-11, 3.952251e-11, 4.053532e-11, 4.029174e-11, 4.059381e-11, 
    4.043952e-11, 4.070406e-11, 4.046593e-11, 4.087889e-11, 4.096911e-11, 
    4.090744e-11, 4.114458e-11, 4.045272e-11, 4.071768e-11, 3.874724e-11, 
    3.875868e-11, 3.8812e-11, 3.857787e-11, 3.856357e-11, 3.834973e-11, 
    3.853997e-11, 3.862113e-11, 3.882758e-11, 3.894995e-11, 3.906647e-11, 
    3.932332e-11, 3.96112e-11, 4.001561e-11, 4.030749e-11, 4.050376e-11, 
    4.038335e-11, 4.048964e-11, 4.037082e-11, 4.031519e-11, 4.093528e-11, 
    4.058647e-11, 4.111041e-11, 4.108133e-11, 4.084385e-11, 4.108459e-11, 
    3.87667e-11, 3.870088e-11, 3.847281e-11, 3.865122e-11, 3.832647e-11, 
    3.850806e-11, 3.861268e-11, 3.901776e-11, 3.910706e-11, 3.918996e-11, 
    3.935395e-11, 3.956494e-11, 3.99365e-11, 4.026126e-11, 4.055896e-11, 
    4.053709e-11, 4.054479e-11, 4.061142e-11, 4.044644e-11, 4.063853e-11, 
    4.06708e-11, 4.058642e-11, 4.107742e-11, 4.093683e-11, 4.108069e-11, 
    4.098911e-11, 3.872226e-11, 3.883307e-11, 3.877316e-11, 3.888584e-11, 
    3.880643e-11, 3.916014e-11, 3.926651e-11, 3.976628e-11, 3.956078e-11, 
    3.988811e-11, 3.959396e-11, 3.964599e-11, 3.989878e-11, 3.960982e-11, 
    4.024329e-11, 3.981321e-11, 4.061401e-11, 4.018243e-11, 4.064112e-11, 
    4.055763e-11, 4.06959e-11, 4.081996e-11, 4.09763e-11, 4.126561e-11, 
    4.119851e-11, 4.144108e-11, 3.899858e-11, 3.914286e-11, 3.913015e-11, 
    3.928143e-11, 3.93935e-11, 3.963701e-11, 4.00292e-11, 3.988147e-11, 
    4.015288e-11, 4.020748e-11, 3.979522e-11, 4.004806e-11, 3.923955e-11, 
    3.936957e-11, 3.929213e-11, 3.900987e-11, 3.991543e-11, 3.944932e-11, 
    4.031227e-11, 4.005809e-11, 4.080224e-11, 4.043125e-11, 4.11616e-11, 
    4.147589e-11, 4.177288e-11, 4.212129e-11, 3.922173e-11, 3.912355e-11, 
    3.929944e-11, 3.954346e-11, 3.97706e-11, 4.007362e-11, 4.010469e-11, 
    4.016161e-11, 4.030926e-11, 4.043362e-11, 4.017959e-11, 4.046481e-11, 
    3.939973e-11, 3.995603e-11, 3.908639e-11, 3.934719e-11, 3.952899e-11, 
    3.944919e-11, 3.986455e-11, 3.996277e-11, 4.036321e-11, 4.015595e-11, 
    4.139818e-11, 4.084614e-11, 4.238762e-11, 4.195382e-11, 3.908927e-11, 
    3.922138e-11, 3.968301e-11, 3.946301e-11, 4.009388e-11, 4.024997e-11, 
    4.03771e-11, 4.05399e-11, 4.05575e-11, 4.065415e-11, 4.049583e-11, 
    4.064788e-11, 4.007421e-11, 4.033004e-11, 3.963006e-11, 3.979982e-11, 
    3.972167e-11, 3.963604e-11, 3.990063e-11, 4.018353e-11, 4.018959e-11, 
    4.028053e-11, 4.053733e-11, 4.009636e-11, 4.146967e-11, 4.061865e-11, 
    3.936571e-11, 3.962132e-11, 3.965791e-11, 3.955874e-11, 4.02343e-11, 
    3.998882e-11, 4.065179e-11, 4.047205e-11, 4.076676e-11, 4.062017e-11, 
    4.059861e-11, 4.04108e-11, 4.029408e-11, 4.000002e-11, 3.976158e-11, 
    3.957306e-11, 3.961685e-11, 3.982409e-11, 4.020086e-11, 4.055902e-11, 
    4.048042e-11, 4.074426e-11, 4.004787e-11, 4.03391e-11, 4.02264e-11, 
    4.05206e-11, 3.987753e-11, 4.042483e-11, 3.973825e-11, 3.97982e-11, 
    3.998394e-11, 4.035896e-11, 4.044219e-11, 4.053113e-11, 4.047623e-11, 
    4.021049e-11, 4.016704e-11, 3.997939e-11, 3.992765e-11, 3.97851e-11, 
    3.966726e-11, 3.97749e-11, 3.98881e-11, 4.021057e-11, 4.050232e-11, 
    4.082166e-11, 4.090002e-11, 4.127515e-11, 4.096961e-11, 4.147441e-11, 
    4.104499e-11, 4.178983e-11, 4.045668e-11, 4.103252e-11, 3.999241e-11, 
    4.010379e-11, 4.030565e-11, 4.077065e-11, 4.051928e-11, 4.081335e-11, 
    4.016533e-11, 3.983125e-11, 3.974506e-11, 3.95845e-11, 3.974873e-11, 
    3.973535e-11, 3.989281e-11, 3.984217e-11, 4.022128e-11, 4.00174e-11, 
    4.0598e-11, 4.081097e-11, 4.141557e-11, 4.178849e-11, 4.216993e-11, 
    4.23389e-11, 4.23904e-11, 4.241194e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.0005857514, 0.0005857557, 0.0005857549, 0.0005857582, 0.0005857564, 
    0.0005857585, 0.0005857524, 0.0005857558, 0.0005857536, 0.0005857519, 
    0.0005857646, 0.0005857584, 0.0005857715, 0.0005857674, 0.0005857777, 
    0.0005857708, 0.0005857791, 0.0005857776, 0.0005857825, 0.0005857811, 
    0.0005857871, 0.0005857831, 0.0005857904, 0.0005857862, 0.0005857868, 
    0.0005857829, 0.0005857597, 0.0005857638, 0.0005857594, 0.00058576, 
    0.0005857598, 0.0005857564, 0.0005857546, 0.0005857512, 0.0005857518, 
    0.0005857544, 0.0005857603, 0.0005857584, 0.0005857634, 0.0005857633, 
    0.0005857689, 0.0005857664, 0.0005857759, 0.0005857732, 0.0005857811, 
    0.0005857791, 0.000585781, 0.0005857804, 0.000585781, 0.0005857781, 
    0.0005857793, 0.0005857768, 0.0005857669, 0.0005857697, 0.0005857611, 
    0.0005857558, 0.0005857525, 0.0005857501, 0.0005857504, 0.000585751, 
    0.0005857544, 0.0005857576, 0.00058576, 0.0005857617, 0.0005857633, 
    0.000585768, 0.0005857706, 0.0005857764, 0.0005857755, 0.0005857772, 
    0.0005857789, 0.0005857818, 0.0005857813, 0.0005857825, 0.0005857772, 
    0.0005857807, 0.0005857749, 0.0005857765, 0.0005857634, 0.0005857589, 
    0.0005857567, 0.000585755, 0.0005857507, 0.0005857536, 0.0005857525, 
    0.0005857553, 0.0005857571, 0.0005857563, 0.0005857617, 0.0005857596, 
    0.0005857708, 0.0005857659, 0.0005857787, 0.0005857756, 0.0005857794, 
    0.0005857775, 0.0005857808, 0.0005857779, 0.000585783, 0.0005857841, 
    0.0005857834, 0.0005857864, 0.0005857777, 0.000585781, 0.0005857562, 
    0.0005857563, 0.000585757, 0.000585754, 0.0005857538, 0.0005857511, 
    0.0005857536, 0.0005857546, 0.0005857573, 0.0005857588, 0.0005857602, 
    0.0005857635, 0.000585767, 0.0005857722, 0.0005857758, 0.0005857783, 
    0.0005857768, 0.0005857782, 0.0005857766, 0.000585776, 0.0005857837, 
    0.0005857793, 0.000585786, 0.0005857855, 0.0005857826, 0.0005857856, 
    0.0005857564, 0.0005857556, 0.0005857527, 0.000585755, 0.0005857509, 
    0.0005857532, 0.0005857545, 0.0005857596, 0.0005857607, 0.0005857618, 
    0.0005857639, 0.0005857665, 0.0005857712, 0.0005857752, 0.000585779, 
    0.0005857787, 0.0005857788, 0.0005857797, 0.0005857776, 0.00058578, 
    0.0005857804, 0.0005857794, 0.0005857855, 0.0005857837, 0.0005857855, 
    0.0005857844, 0.0005857559, 0.0005857573, 0.0005857566, 0.000585758, 
    0.0005857569, 0.0005857613, 0.0005857627, 0.000585769, 0.0005857665, 
    0.0005857705, 0.0005857669, 0.0005857675, 0.0005857705, 0.0005857671, 
    0.0005857749, 0.0005857695, 0.0005857797, 0.0005857741, 0.0005857801, 
    0.000585779, 0.0005857808, 0.0005857823, 0.0005857843, 0.0005857878, 
    0.000585787, 0.00058579, 0.0005857594, 0.0005857612, 0.000585761, 
    0.000585763, 0.0005857644, 0.0005857674, 0.0005857723, 0.0005857705, 
    0.0005857739, 0.0005857746, 0.0005857694, 0.0005857726, 0.0005857624, 
    0.0005857639, 0.0005857631, 0.0005857595, 0.0005857709, 0.000585765, 
    0.0005857759, 0.0005857727, 0.0005857821, 0.0005857773, 0.0005857865, 
    0.0005857904, 0.0005857942, 0.0005857984, 0.0005857622, 0.000585761, 
    0.0005857632, 0.0005857662, 0.0005857691, 0.0005857729, 0.0005857733, 
    0.000585774, 0.0005857759, 0.0005857775, 0.0005857742, 0.0005857779, 
    0.0005857642, 0.0005857714, 0.0005857605, 0.0005857637, 0.000585766, 
    0.0005857651, 0.0005857703, 0.0005857715, 0.0005857765, 0.000585774, 
    0.0005857894, 0.0005857825, 0.0005858018, 0.0005857964, 0.0005857605, 
    0.0005857622, 0.000585768, 0.0005857652, 0.0005857732, 0.0005857751, 
    0.0005857768, 0.0005857787, 0.000585779, 0.0005857802, 0.0005857782, 
    0.0005857801, 0.0005857729, 0.0005857761, 0.0005857674, 0.0005857695, 
    0.0005857685, 0.0005857674, 0.0005857708, 0.0005857743, 0.0005857744, 
    0.0005857755, 0.0005857784, 0.0005857732, 0.0005857901, 0.0005857795, 
    0.000585764, 0.0005857671, 0.0005857677, 0.0005857665, 0.0005857749, 
    0.0005857719, 0.0005857802, 0.0005857779, 0.0005857816, 0.0005857798, 
    0.0005857795, 0.0005857772, 0.0005857757, 0.000585772, 0.000585769, 
    0.0005857666, 0.0005857672, 0.0005857698, 0.0005857745, 0.000585779, 
    0.000585778, 0.0005857814, 0.0005857726, 0.0005857762, 0.0005857748, 
    0.0005857786, 0.0005857705, 0.000585777, 0.0005857687, 0.0005857695, 
    0.0005857718, 0.0005857764, 0.0005857776, 0.0005857786, 0.000585778, 
    0.0005857746, 0.0005857741, 0.0005857717, 0.000585771, 0.0005857693, 
    0.0005857678, 0.0005857692, 0.0005857705, 0.0005857747, 0.0005857783, 
    0.0005857823, 0.0005857833, 0.0005857878, 0.000585784, 0.0005857901, 
    0.0005857847, 0.0005857942, 0.0005857776, 0.0005857848, 0.0005857719, 
    0.0005857733, 0.0005857758, 0.0005857816, 0.0005857785, 0.0005857821, 
    0.0005857741, 0.0005857698, 0.0005857688, 0.0005857667, 0.0005857688, 
    0.0005857687, 0.0005857706, 0.0005857701, 0.0005857748, 0.0005857722, 
    0.0005857795, 0.0005857821, 0.0005857897, 0.0005857943, 0.0005857992, 
    0.0005858013, 0.0005858019, 0.0005858022 ;

 QBOT =
  0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  9.506026e-06, 9.530893e-06, 9.526066e-06, 9.546117e-06, 9.535007e-06, 
    9.548128e-06, 9.511082e-06, 9.531866e-06, 9.518605e-06, 9.508286e-06, 
    9.585023e-06, 9.547017e-06, 9.624719e-06, 9.600413e-06, 9.661561e-06, 
    9.620912e-06, 9.669772e-06, 9.660427e-06, 9.688658e-06, 9.68057e-06, 
    9.716624e-06, 9.692391e-06, 9.735395e-06, 9.710857e-06, 9.714679e-06, 
    9.691586e-06, 9.554697e-06, 9.580276e-06, 9.553174e-06, 9.556822e-06, 
    9.555194e-06, 9.535223e-06, 9.52514e-06, 9.504152e-06, 9.507968e-06, 
    9.523397e-06, 9.558464e-06, 9.54658e-06, 9.576614e-06, 9.575936e-06, 
    9.609384e-06, 9.594297e-06, 9.650604e-06, 9.634598e-06, 9.680908e-06, 
    9.669248e-06, 9.680353e-06, 9.676991e-06, 9.680397e-06, 9.663302e-06, 
    9.670623e-06, 9.655597e-06, 9.597115e-06, 9.614278e-06, 9.563101e-06, 
    9.532318e-06, 9.511986e-06, 9.497542e-06, 9.499583e-06, 9.503467e-06, 
    9.523487e-06, 9.542358e-06, 9.556737e-06, 9.566354e-06, 9.575838e-06, 
    9.604465e-06, 9.619714e-06, 9.653822e-06, 9.647697e-06, 9.658101e-06, 
    9.668091e-06, 9.684825e-06, 9.682076e-06, 9.689443e-06, 9.657851e-06, 
    9.678831e-06, 9.644201e-06, 9.653664e-06, 9.578286e-06, 9.549792e-06, 
    9.537578e-06, 9.526989e-06, 9.50115e-06, 9.518983e-06, 9.511949e-06, 
    9.528716e-06, 9.539358e-06, 9.5341e-06, 9.566617e-06, 9.553965e-06, 
    9.620618e-06, 9.591889e-06, 9.666926e-06, 9.648957e-06, 9.671238e-06, 
    9.659873e-06, 9.679339e-06, 9.66182e-06, 9.692196e-06, 9.6988e-06, 
    9.694284e-06, 9.711677e-06, 9.660846e-06, 9.680341e-06, 9.533946e-06, 
    9.534803e-06, 9.53881e-06, 9.521198e-06, 9.520129e-06, 9.504041e-06, 
    9.518367e-06, 9.52446e-06, 9.539986e-06, 9.549149e-06, 9.557871e-06, 
    9.577059e-06, 9.598484e-06, 9.628508e-06, 9.65012e-06, 9.66461e-06, 
    9.655732e-06, 9.663569e-06, 9.654804e-06, 9.650703e-06, 9.696316e-06, 
    9.670684e-06, 9.709175e-06, 9.707049e-06, 9.689613e-06, 9.707288e-06, 
    9.535407e-06, 9.530473e-06, 9.513307e-06, 9.52674e-06, 9.502292e-06, 
    9.515956e-06, 9.523808e-06, 9.554202e-06, 9.560915e-06, 9.567101e-06, 
    9.579353e-06, 9.595068e-06, 9.622651e-06, 9.646693e-06, 9.668677e-06, 
    9.667068e-06, 9.667634e-06, 9.672533e-06, 9.66038e-06, 9.674531e-06, 
    9.676894e-06, 9.670696e-06, 9.706763e-06, 9.696456e-06, 9.707003e-06, 
    9.700295e-06, 9.53208e-06, 9.540389e-06, 9.535897e-06, 9.544337e-06, 
    9.53838e-06, 9.564844e-06, 9.572783e-06, 9.609998e-06, 9.594752e-06, 
    9.619057e-06, 9.59723e-06, 9.601089e-06, 9.619795e-06, 9.598418e-06, 
    9.645341e-06, 9.613471e-06, 9.672724e-06, 9.640814e-06, 9.674722e-06, 
    9.668583e-06, 9.678762e-06, 9.687867e-06, 9.69935e-06, 9.720511e-06, 
    9.715615e-06, 9.733342e-06, 9.552793e-06, 9.563568e-06, 9.562644e-06, 
    9.573941e-06, 9.582293e-06, 9.600436e-06, 9.629531e-06, 9.618594e-06, 
    9.638702e-06, 9.642732e-06, 9.612199e-06, 9.630919e-06, 9.5708e-06, 
    9.580478e-06, 9.574734e-06, 9.553629e-06, 9.62108e-06, 9.586428e-06, 
    9.650473e-06, 9.631681e-06, 9.686565e-06, 9.659231e-06, 9.712915e-06, 
    9.735828e-06, 9.757526e-06, 9.782765e-06, 9.569477e-06, 9.562151e-06, 
    9.575291e-06, 9.593437e-06, 9.610354e-06, 9.632822e-06, 9.635135e-06, 
    9.63934e-06, 9.650263e-06, 9.659438e-06, 9.640645e-06, 9.661741e-06, 
    9.582674e-06, 9.624101e-06, 9.559359e-06, 9.578805e-06, 9.592378e-06, 
    9.586448e-06, 9.617351e-06, 9.62463e-06, 9.654223e-06, 9.638936e-06, 
    9.730149e-06, 9.689756e-06, 9.802081e-06, 9.770632e-06, 9.559586e-06, 
    9.569463e-06, 9.603832e-06, 9.587478e-06, 9.634336e-06, 9.645871e-06, 
    9.655273e-06, 9.667256e-06, 9.668568e-06, 9.675674e-06, 9.664028e-06, 
    9.675223e-06, 9.632869e-06, 9.651792e-06, 9.59993e-06, 9.61253e-06, 
    9.606742e-06, 9.600375e-06, 9.620025e-06, 9.640935e-06, 9.641421e-06, 
    9.648123e-06, 9.666943e-06, 9.634527e-06, 9.735292e-06, 9.672952e-06, 
    9.580235e-06, 9.599224e-06, 9.601986e-06, 9.594619e-06, 9.644713e-06, 
    9.626547e-06, 9.675507e-06, 9.662274e-06, 9.683969e-06, 9.673183e-06, 
    9.671594e-06, 9.657758e-06, 9.649136e-06, 9.627372e-06, 9.609687e-06, 
    9.595692e-06, 9.598949e-06, 9.614325e-06, 9.642224e-06, 9.668669e-06, 
    9.662868e-06, 9.68232e-06, 9.630934e-06, 9.652449e-06, 9.644118e-06, 
    9.665852e-06, 9.618295e-06, 9.658666e-06, 9.60797e-06, 9.61242e-06, 
    9.626187e-06, 9.653882e-06, 9.660072e-06, 9.666612e-06, 9.662584e-06, 
    9.642939e-06, 9.63974e-06, 9.625861e-06, 9.622011e-06, 9.611455e-06, 
    9.602699e-06, 9.610688e-06, 9.619073e-06, 9.642964e-06, 9.664489e-06, 
    9.68799e-06, 9.69376e-06, 9.721147e-06, 9.698796e-06, 9.735632e-06, 
    9.704228e-06, 9.758653e-06, 9.661067e-06, 9.703386e-06, 9.626826e-06, 
    9.635074e-06, 9.649955e-06, 9.684202e-06, 9.66575e-06, 9.68735e-06, 
    9.639618e-06, 9.614836e-06, 9.608477e-06, 9.596536e-06, 9.608751e-06, 
    9.607758e-06, 9.619449e-06, 9.615694e-06, 9.643758e-06, 9.628681e-06, 
    9.671544e-06, 9.68719e-06, 9.73147e-06, 9.758622e-06, 9.786349e-06, 
    9.798578e-06, 9.802304e-06, 9.803858e-06 ;

 QVEGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  81.68618, 81.68539, 81.68554, 81.6849, 81.68525, 81.68484, 81.68601, 
    81.68536, 81.68578, 81.6861, 81.68369, 81.68487, 81.6824, 81.68316, 
    81.68121, 81.68252, 81.68095, 81.68124, 81.68033, 81.68059, 81.67946, 
    81.68021, 81.67885, 81.67963, 81.67951, 81.68024, 81.68462, 81.68384, 
    81.68467, 81.68456, 81.6846, 81.68524, 81.68558, 81.68623, 81.68611, 
    81.68562, 81.6845, 81.68488, 81.68391, 81.68393, 81.68287, 81.68335, 
    81.68155, 81.68206, 81.68057, 81.68095, 81.6806, 81.6807, 81.6806, 
    81.68114, 81.68091, 81.68139, 81.68327, 81.68272, 81.68435, 81.68536, 
    81.68599, 81.68645, 81.68638, 81.68626, 81.68562, 81.68501, 81.68455, 
    81.68424, 81.68394, 81.68305, 81.68256, 81.68146, 81.68164, 81.68132, 
    81.68098, 81.68046, 81.68054, 81.68031, 81.68131, 81.68065, 81.68175, 
    81.68145, 81.68391, 81.68478, 81.68519, 81.68551, 81.68633, 81.68577, 
    81.68599, 81.68545, 81.6851, 81.68527, 81.68423, 81.68464, 81.68253, 
    81.68343, 81.68103, 81.6816, 81.68089, 81.68125, 81.68063, 81.68119, 
    81.68022, 81.68002, 81.68015, 81.6796, 81.68122, 81.6806, 81.68528, 
    81.68525, 81.68512, 81.6857, 81.68573, 81.68624, 81.68578, 81.68559, 
    81.68508, 81.68479, 81.68452, 81.6839, 81.68323, 81.68227, 81.68156, 
    81.6811, 81.68138, 81.68113, 81.68141, 81.68154, 81.68009, 81.68091, 
    81.67967, 81.67974, 81.68031, 81.67973, 81.68523, 81.68539, 81.68594, 
    81.68551, 81.68629, 81.68586, 81.68562, 81.68464, 81.68442, 81.68422, 
    81.68383, 81.68333, 81.68245, 81.68168, 81.68097, 81.68102, 81.681, 
    81.68085, 81.68124, 81.68079, 81.68071, 81.68091, 81.67975, 81.68008, 
    81.67974, 81.67995, 81.68533, 81.68507, 81.68522, 81.68495, 81.68514, 
    81.6843, 81.68405, 81.68286, 81.68334, 81.68256, 81.68326, 81.68314, 
    81.68256, 81.68321, 81.68173, 81.68275, 81.68084, 81.68188, 81.68078, 
    81.68097, 81.68064, 81.68036, 81.67999, 81.67932, 81.67947, 81.6789, 
    81.68468, 81.68434, 81.68436, 81.684, 81.68374, 81.68315, 81.68223, 
    81.68257, 81.68192, 81.6818, 81.68278, 81.68218, 81.6841, 81.68381, 
    81.68398, 81.68465, 81.6825, 81.68362, 81.68156, 81.68215, 81.6804, 
    81.68128, 81.67956, 81.67885, 81.67813, 81.67735, 81.68414, 81.68437, 
    81.68395, 81.68339, 81.68284, 81.68212, 81.68204, 81.68191, 81.68156, 
    81.68127, 81.68188, 81.68119, 81.68375, 81.6824, 81.68447, 81.68386, 
    81.68342, 81.6836, 81.68261, 81.68237, 81.68144, 81.68192, 81.67903, 
    81.68031, 81.67671, 81.67773, 81.68446, 81.68414, 81.68305, 81.68357, 
    81.68207, 81.6817, 81.6814, 81.68102, 81.68097, 81.68075, 81.68111, 
    81.68076, 81.68212, 81.68151, 81.68317, 81.68277, 81.68295, 81.68315, 
    81.68253, 81.68187, 81.68184, 81.68163, 81.68108, 81.68206, 81.67889, 
    81.68088, 81.6838, 81.6832, 81.68311, 81.68333, 81.68174, 81.68232, 
    81.68075, 81.68118, 81.68048, 81.68082, 81.68088, 81.68132, 81.68159, 
    81.6823, 81.68286, 81.6833, 81.6832, 81.68272, 81.68182, 81.68098, 
    81.68117, 81.68053, 81.68217, 81.6815, 81.68176, 81.68106, 81.68259, 
    81.68134, 81.68291, 81.68277, 81.68233, 81.68146, 81.68124, 81.68104, 
    81.68116, 81.6818, 81.6819, 81.68233, 81.68246, 81.6828, 81.68307, 
    81.68282, 81.68256, 81.68179, 81.68111, 81.68036, 81.68017, 81.67932, 
    81.68003, 81.67889, 81.67989, 81.67813, 81.68124, 81.67989, 81.6823, 
    81.68204, 81.68158, 81.68049, 81.68106, 81.68039, 81.6819, 81.68271, 
    81.68289, 81.68327, 81.68288, 81.68291, 81.68254, 81.68266, 81.68177, 
    81.68224, 81.68089, 81.68039, 81.67897, 81.67811, 81.67721, 81.67682, 
    81.6767, 81.67664 ;

 RH2M_R =
  81.68618, 81.68539, 81.68554, 81.6849, 81.68525, 81.68484, 81.68601, 
    81.68536, 81.68578, 81.6861, 81.68369, 81.68487, 81.6824, 81.68316, 
    81.68121, 81.68252, 81.68095, 81.68124, 81.68033, 81.68059, 81.67946, 
    81.68021, 81.67885, 81.67963, 81.67951, 81.68024, 81.68462, 81.68384, 
    81.68467, 81.68456, 81.6846, 81.68524, 81.68558, 81.68623, 81.68611, 
    81.68562, 81.6845, 81.68488, 81.68391, 81.68393, 81.68287, 81.68335, 
    81.68155, 81.68206, 81.68057, 81.68095, 81.6806, 81.6807, 81.6806, 
    81.68114, 81.68091, 81.68139, 81.68327, 81.68272, 81.68435, 81.68536, 
    81.68599, 81.68645, 81.68638, 81.68626, 81.68562, 81.68501, 81.68455, 
    81.68424, 81.68394, 81.68305, 81.68256, 81.68146, 81.68164, 81.68132, 
    81.68098, 81.68046, 81.68054, 81.68031, 81.68131, 81.68065, 81.68175, 
    81.68145, 81.68391, 81.68478, 81.68519, 81.68551, 81.68633, 81.68577, 
    81.68599, 81.68545, 81.6851, 81.68527, 81.68423, 81.68464, 81.68253, 
    81.68343, 81.68103, 81.6816, 81.68089, 81.68125, 81.68063, 81.68119, 
    81.68022, 81.68002, 81.68015, 81.6796, 81.68122, 81.6806, 81.68528, 
    81.68525, 81.68512, 81.6857, 81.68573, 81.68624, 81.68578, 81.68559, 
    81.68508, 81.68479, 81.68452, 81.6839, 81.68323, 81.68227, 81.68156, 
    81.6811, 81.68138, 81.68113, 81.68141, 81.68154, 81.68009, 81.68091, 
    81.67967, 81.67974, 81.68031, 81.67973, 81.68523, 81.68539, 81.68594, 
    81.68551, 81.68629, 81.68586, 81.68562, 81.68464, 81.68442, 81.68422, 
    81.68383, 81.68333, 81.68245, 81.68168, 81.68097, 81.68102, 81.681, 
    81.68085, 81.68124, 81.68079, 81.68071, 81.68091, 81.67975, 81.68008, 
    81.67974, 81.67995, 81.68533, 81.68507, 81.68522, 81.68495, 81.68514, 
    81.6843, 81.68405, 81.68286, 81.68334, 81.68256, 81.68326, 81.68314, 
    81.68256, 81.68321, 81.68173, 81.68275, 81.68084, 81.68188, 81.68078, 
    81.68097, 81.68064, 81.68036, 81.67999, 81.67932, 81.67947, 81.6789, 
    81.68468, 81.68434, 81.68436, 81.684, 81.68374, 81.68315, 81.68223, 
    81.68257, 81.68192, 81.6818, 81.68278, 81.68218, 81.6841, 81.68381, 
    81.68398, 81.68465, 81.6825, 81.68362, 81.68156, 81.68215, 81.6804, 
    81.68128, 81.67956, 81.67885, 81.67813, 81.67735, 81.68414, 81.68437, 
    81.68395, 81.68339, 81.68284, 81.68212, 81.68204, 81.68191, 81.68156, 
    81.68127, 81.68188, 81.68119, 81.68375, 81.6824, 81.68447, 81.68386, 
    81.68342, 81.6836, 81.68261, 81.68237, 81.68144, 81.68192, 81.67903, 
    81.68031, 81.67671, 81.67773, 81.68446, 81.68414, 81.68305, 81.68357, 
    81.68207, 81.6817, 81.6814, 81.68102, 81.68097, 81.68075, 81.68111, 
    81.68076, 81.68212, 81.68151, 81.68317, 81.68277, 81.68295, 81.68315, 
    81.68253, 81.68187, 81.68184, 81.68163, 81.68108, 81.68206, 81.67889, 
    81.68088, 81.6838, 81.6832, 81.68311, 81.68333, 81.68174, 81.68232, 
    81.68075, 81.68118, 81.68048, 81.68082, 81.68088, 81.68132, 81.68159, 
    81.6823, 81.68286, 81.6833, 81.6832, 81.68272, 81.68182, 81.68098, 
    81.68117, 81.68053, 81.68217, 81.6815, 81.68176, 81.68106, 81.68259, 
    81.68134, 81.68291, 81.68277, 81.68233, 81.68146, 81.68124, 81.68104, 
    81.68116, 81.6818, 81.6819, 81.68233, 81.68246, 81.6828, 81.68307, 
    81.68282, 81.68256, 81.68179, 81.68111, 81.68036, 81.68017, 81.67932, 
    81.68003, 81.67889, 81.67989, 81.67813, 81.68124, 81.67989, 81.6823, 
    81.68204, 81.68158, 81.68049, 81.68106, 81.68039, 81.6819, 81.68271, 
    81.68289, 81.68327, 81.68288, 81.68291, 81.68254, 81.68266, 81.68177, 
    81.68224, 81.68089, 81.68039, 81.67897, 81.67811, 81.67721, 81.67682, 
    81.6767, 81.67664 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004365606, 0.0004384049, 0.0004380463, 0.0004395339, 0.0004387087, 
    0.0004396826, 0.0004369343, 0.0004384778, 0.0004374924, 0.0004367262, 
    0.0004424202, 0.0004395998, 0.0004453503, 0.0004435513, 0.0004480703, 
    0.0004450702, 0.0004486752, 0.0004479837, 0.0004500649, 0.0004494686, 
    0.0004521304, 0.00045034, 0.0004535103, 0.0004517028, 0.0004519854, 
    0.0004502806, 0.0004401679, 0.0004420695, 0.0004400551, 0.0004403263, 
    0.0004402045, 0.0004387254, 0.0004379801, 0.0004364192, 0.0004367025, 
    0.0004378489, 0.0004404478, 0.0004395655, 0.000441789, 0.0004417388, 
    0.0004442141, 0.000443098, 0.0004472587, 0.0004460761, 0.0004494934, 
    0.0004486339, 0.0004494529, 0.0004492045, 0.000449456, 0.0004481956, 
    0.0004487355, 0.0004476264, 0.0004433077, 0.0004445771, 0.0004407907, 
    0.0004385138, 0.0004370017, 0.0004359287, 0.0004360803, 0.0004363695, 
    0.0004378555, 0.0004392526, 0.0004403175, 0.0004410296, 0.0004417314, 
    0.0004438556, 0.00044498, 0.0004474977, 0.0004470434, 0.000447813, 
    0.0004485483, 0.0004497828, 0.0004495796, 0.0004501234, 0.0004477924, 
    0.0004493415, 0.0004467841, 0.0004474835, 0.0004419225, 0.0004398038, 
    0.000438903, 0.0004381147, 0.0004361969, 0.0004375213, 0.0004369991, 
    0.0004382411, 0.0004390304, 0.00043864, 0.0004410491, 0.0004401123, 
    0.0004450466, 0.0004429212, 0.0004484626, 0.0004471365, 0.0004487803, 
    0.0004479415, 0.0004493786, 0.0004480851, 0.0004503258, 0.0004508137, 
    0.0004504801, 0.000451761, 0.0004480131, 0.0004494523, 0.0004386293, 
    0.000438693, 0.0004389895, 0.0004376856, 0.0004376059, 0.000436411, 
    0.0004374741, 0.0004379268, 0.000439076, 0.0004397556, 0.0004404018, 
    0.0004418226, 0.0004434093, 0.0004456282, 0.0004472224, 0.0004482909, 
    0.0004476357, 0.0004482141, 0.0004475673, 0.0004472641, 0.0004506307, 
    0.0004487403, 0.0004515766, 0.0004514197, 0.0004501359, 0.0004514372, 
    0.0004387376, 0.0004383711, 0.0004370991, 0.0004380945, 0.0004362808, 
    0.000437296, 0.0004378796, 0.0004401318, 0.0004406266, 0.0004410855, 
    0.0004419917, 0.0004431547, 0.000445195, 0.0004469702, 0.0004485909, 
    0.0004484721, 0.0004485138, 0.0004488758, 0.000447979, 0.0004490229, 
    0.000449198, 0.0004487399, 0.0004513985, 0.000450639, 0.0004514162, 
    0.0004509215, 0.0004384902, 0.0004391065, 0.0004387734, 0.0004393997, 
    0.0004389583, 0.0004409205, 0.0004415087, 0.0004442616, 0.0004431318, 
    0.0004449299, 0.0004433143, 0.0004436006, 0.0004449883, 0.0004434015, 
    0.0004468721, 0.000444519, 0.0004488898, 0.0004465398, 0.0004490369, 
    0.0004485834, 0.0004493341, 0.0004500065, 0.0004508523, 0.000452413, 
    0.0004520515, 0.0004533568, 0.0004400255, 0.0004408249, 0.0004407545, 
    0.0004415912, 0.0004422099, 0.0004435513, 0.0004457025, 0.0004448934, 
    0.0004463785, 0.0004466767, 0.0004444203, 0.0004458056, 0.0004413595, 
    0.0004420776, 0.00044165, 0.0004400877, 0.0004450793, 0.0004425174, 
    0.0004472481, 0.0004458601, 0.0004499104, 0.0004478961, 0.0004518525, 
    0.0004535438, 0.0004551358, 0.0004569959, 0.0004412612, 0.0004407179, 
    0.0004416906, 0.0004430364, 0.0004442852, 0.0004459455, 0.0004461153, 
    0.0004464262, 0.0004472318, 0.0004479092, 0.0004465244, 0.0004480789, 
    0.0004422441, 0.0004453017, 0.0004405117, 0.000441954, 0.0004429564, 
    0.0004425167, 0.0004448003, 0.0004453384, 0.0004475255, 0.0004463949, 
    0.0004531262, 0.000450148, 0.0004584124, 0.0004561027, 0.000440528, 
    0.0004412592, 0.000443804, 0.0004425932, 0.0004460561, 0.0004469086, 
    0.0004476015, 0.0004484873, 0.0004485828, 0.0004491077, 0.0004482475, 
    0.0004490736, 0.0004459484, 0.0004473449, 0.0004435126, 0.0004444452, 
    0.0004440162, 0.0004435454, 0.000444998, 0.0004465455, 0.0004465786, 
    0.0004470747, 0.0004484729, 0.0004460692, 0.0004535102, 0.0004489145, 
    0.0004420565, 0.0004434648, 0.000443666, 0.0004431204, 0.000446823, 
    0.0004454813, 0.0004490949, 0.0004481182, 0.0004497183, 0.0004489232, 
    0.000448806, 0.0004477848, 0.0004471488, 0.0004455424, 0.0004442353, 
    0.0004431989, 0.0004434398, 0.0004445782, 0.0004466401, 0.0004485908, 
    0.0004481634, 0.000449596, 0.0004458039, 0.0004473939, 0.0004467792, 
    0.0004483818, 0.0004448717, 0.0004478614, 0.0004441074, 0.0004444365, 
    0.0004454546, 0.0004475026, 0.0004479557, 0.0004484394, 0.0004481408, 
    0.0004466928, 0.0004464556, 0.0004454295, 0.0004451461, 0.0004443643, 
    0.000443717, 0.0004443083, 0.0004449292, 0.000446693, 0.0004482825, 
    0.0004500154, 0.0004504395, 0.000452464, 0.0004508157, 0.0004535355, 
    0.000451223, 0.0004552261, 0.0004480347, 0.0004511562, 0.0004455009, 
    0.0004461101, 0.000447212, 0.0004497394, 0.0004483749, 0.0004499706, 
    0.0004464462, 0.0004446176, 0.0004441445, 0.0004432618, 0.0004441646, 
    0.0004440912, 0.000444955, 0.0004446773, 0.0004467515, 0.0004456373, 
    0.0004488023, 0.0004499574, 0.0004532194, 0.000455219, 0.0004572547, 
    0.0004581533, 0.0004584268, 0.0004585411 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.502156e-14, 3.511612e-14, 3.509775e-14, 3.517395e-14, 3.51317e-14, 
    3.518158e-14, 3.504075e-14, 3.511986e-14, 3.506937e-14, 3.503009e-14, 
    3.532161e-14, 3.517735e-14, 3.54713e-14, 3.537948e-14, 3.561e-14, 
    3.545701e-14, 3.564082e-14, 3.560561e-14, 3.571158e-14, 3.568124e-14, 
    3.581657e-14, 3.572558e-14, 3.588667e-14, 3.579486e-14, 3.580922e-14, 
    3.572257e-14, 3.520643e-14, 3.530365e-14, 3.520066e-14, 3.521453e-14, 
    3.520831e-14, 3.513257e-14, 3.509435e-14, 3.501434e-14, 3.502888e-14, 
    3.508765e-14, 3.522077e-14, 3.517562e-14, 3.528942e-14, 3.528685e-14, 
    3.541334e-14, 3.535633e-14, 3.556868e-14, 3.550838e-14, 3.568251e-14, 
    3.563875e-14, 3.568045e-14, 3.566781e-14, 3.568061e-14, 3.561643e-14, 
    3.564393e-14, 3.558744e-14, 3.536701e-14, 3.543184e-14, 3.523831e-14, 
    3.512169e-14, 3.504422e-14, 3.498917e-14, 3.499696e-14, 3.501179e-14, 
    3.508799e-14, 3.51596e-14, 3.521413e-14, 3.525058e-14, 3.528648e-14, 
    3.539499e-14, 3.545243e-14, 3.558085e-14, 3.555771e-14, 3.559692e-14, 
    3.563439e-14, 3.569724e-14, 3.56869e-14, 3.571458e-14, 3.55959e-14, 
    3.567478e-14, 3.554452e-14, 3.558017e-14, 3.529614e-14, 3.518781e-14, 
    3.514164e-14, 3.510128e-14, 3.500294e-14, 3.507086e-14, 3.504409e-14, 
    3.510778e-14, 3.514822e-14, 3.512822e-14, 3.525157e-14, 3.520363e-14, 
    3.545583e-14, 3.534729e-14, 3.563002e-14, 3.556246e-14, 3.564621e-14, 
    3.560349e-14, 3.567667e-14, 3.561081e-14, 3.572488e-14, 3.574968e-14, 
    3.573273e-14, 3.579786e-14, 3.560716e-14, 3.568044e-14, 3.512766e-14, 
    3.513092e-14, 3.514612e-14, 3.507929e-14, 3.50752e-14, 3.501394e-14, 
    3.506846e-14, 3.509166e-14, 3.515057e-14, 3.518537e-14, 3.521845e-14, 
    3.529114e-14, 3.537223e-14, 3.548553e-14, 3.556684e-14, 3.56213e-14, 
    3.558792e-14, 3.561739e-14, 3.558444e-14, 3.556899e-14, 3.574038e-14, 
    3.564418e-14, 3.57885e-14, 3.578052e-14, 3.571523e-14, 3.578142e-14, 
    3.513321e-14, 3.511445e-14, 3.504923e-14, 3.510027e-14, 3.500727e-14, 
    3.505933e-14, 3.508924e-14, 3.520462e-14, 3.522997e-14, 3.525344e-14, 
    3.52998e-14, 3.535925e-14, 3.546343e-14, 3.555398e-14, 3.563658e-14, 
    3.563053e-14, 3.563266e-14, 3.565109e-14, 3.560542e-14, 3.565859e-14, 
    3.56675e-14, 3.564418e-14, 3.577945e-14, 3.574083e-14, 3.578035e-14, 
    3.575521e-14, 3.512055e-14, 3.515212e-14, 3.513506e-14, 3.516714e-14, 
    3.514454e-14, 3.524498e-14, 3.527507e-14, 3.541577e-14, 3.535808e-14, 
    3.544989e-14, 3.536741e-14, 3.538203e-14, 3.545285e-14, 3.537188e-14, 
    3.554898e-14, 3.542891e-14, 3.565181e-14, 3.553202e-14, 3.56593e-14, 
    3.563622e-14, 3.567445e-14, 3.570865e-14, 3.575169e-14, 3.5831e-14, 
    3.581264e-14, 3.587894e-14, 3.519919e-14, 3.524009e-14, 3.523651e-14, 
    3.527932e-14, 3.531095e-14, 3.537951e-14, 3.548933e-14, 3.544806e-14, 
    3.552383e-14, 3.553903e-14, 3.542391e-14, 3.54946e-14, 3.526748e-14, 
    3.530419e-14, 3.528235e-14, 3.52024e-14, 3.545754e-14, 3.532669e-14, 
    3.556818e-14, 3.549742e-14, 3.570377e-14, 3.560119e-14, 3.580253e-14, 
    3.58884e-14, 3.596922e-14, 3.606345e-14, 3.526243e-14, 3.523464e-14, 
    3.528441e-14, 3.535318e-14, 3.5417e-14, 3.550173e-14, 3.55104e-14, 
    3.552626e-14, 3.556734e-14, 3.560186e-14, 3.553126e-14, 3.561052e-14, 
    3.531267e-14, 3.54689e-14, 3.522412e-14, 3.529788e-14, 3.534914e-14, 
    3.532667e-14, 3.544334e-14, 3.547081e-14, 3.558233e-14, 3.552471e-14, 
    3.58672e-14, 3.571585e-14, 3.613519e-14, 3.601822e-14, 3.522493e-14, 
    3.526234e-14, 3.539242e-14, 3.533056e-14, 3.550739e-14, 3.555086e-14, 
    3.558619e-14, 3.56313e-14, 3.563618e-14, 3.56629e-14, 3.561911e-14, 
    3.566117e-14, 3.550191e-14, 3.557312e-14, 3.537758e-14, 3.542521e-14, 
    3.540331e-14, 3.537927e-14, 3.545344e-14, 3.553236e-14, 3.553408e-14, 
    3.555936e-14, 3.563053e-14, 3.550811e-14, 3.588667e-14, 3.565304e-14, 
    3.530313e-14, 3.537508e-14, 3.538539e-14, 3.535752e-14, 3.55465e-14, 
    3.547807e-14, 3.566225e-14, 3.561252e-14, 3.5694e-14, 3.565352e-14, 
    3.564756e-14, 3.559554e-14, 3.556313e-14, 3.54812e-14, 3.541449e-14, 
    3.536157e-14, 3.537387e-14, 3.5432e-14, 3.55372e-14, 3.563661e-14, 
    3.561484e-14, 3.568781e-14, 3.549458e-14, 3.557564e-14, 3.554431e-14, 
    3.562599e-14, 3.544695e-14, 3.559935e-14, 3.540795e-14, 3.542475e-14, 
    3.547671e-14, 3.558112e-14, 3.560425e-14, 3.562888e-14, 3.561369e-14, 
    3.553987e-14, 3.552778e-14, 3.547545e-14, 3.546099e-14, 3.54211e-14, 
    3.538804e-14, 3.541823e-14, 3.544992e-14, 3.553991e-14, 3.562091e-14, 
    3.570914e-14, 3.573072e-14, 3.583358e-14, 3.574982e-14, 3.588796e-14, 
    3.577047e-14, 3.597376e-14, 3.560821e-14, 3.576707e-14, 3.547908e-14, 
    3.551017e-14, 3.556632e-14, 3.569504e-14, 3.562561e-14, 3.570682e-14, 
    3.552731e-14, 3.543399e-14, 3.540987e-14, 3.536478e-14, 3.54109e-14, 
    3.540715e-14, 3.545126e-14, 3.543709e-14, 3.55429e-14, 3.548608e-14, 
    3.56474e-14, 3.570618e-14, 3.587199e-14, 3.597344e-14, 3.607662e-14, 
    3.612212e-14, 3.613596e-14, 3.614175e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.164501e-14, 1.167648e-14, 1.167037e-14, 1.169573e-14, 1.168167e-14, 
    1.169827e-14, 1.16514e-14, 1.167773e-14, 1.166092e-14, 1.164785e-14, 
    1.174488e-14, 1.169687e-14, 1.179471e-14, 1.176414e-14, 1.184087e-14, 
    1.178995e-14, 1.185113e-14, 1.183941e-14, 1.187469e-14, 1.186459e-14, 
    1.190963e-14, 1.187935e-14, 1.193297e-14, 1.190241e-14, 1.190719e-14, 
    1.187835e-14, 1.170654e-14, 1.17389e-14, 1.170462e-14, 1.170924e-14, 
    1.170717e-14, 1.168196e-14, 1.166924e-14, 1.164261e-14, 1.164745e-14, 
    1.166701e-14, 1.171132e-14, 1.169629e-14, 1.173417e-14, 1.173331e-14, 
    1.177541e-14, 1.175644e-14, 1.182712e-14, 1.180705e-14, 1.186501e-14, 
    1.185044e-14, 1.186432e-14, 1.186012e-14, 1.186438e-14, 1.184301e-14, 
    1.185217e-14, 1.183336e-14, 1.175999e-14, 1.178157e-14, 1.171715e-14, 
    1.167834e-14, 1.165255e-14, 1.163423e-14, 1.163682e-14, 1.164176e-14, 
    1.166712e-14, 1.169096e-14, 1.17091e-14, 1.172124e-14, 1.173319e-14, 
    1.176931e-14, 1.178842e-14, 1.183117e-14, 1.182347e-14, 1.183652e-14, 
    1.184899e-14, 1.186991e-14, 1.186647e-14, 1.187568e-14, 1.183618e-14, 
    1.186244e-14, 1.181908e-14, 1.183094e-14, 1.17364e-14, 1.170035e-14, 
    1.168498e-14, 1.167154e-14, 1.163881e-14, 1.166142e-14, 1.165251e-14, 
    1.167371e-14, 1.168717e-14, 1.168051e-14, 1.172157e-14, 1.170561e-14, 
    1.178956e-14, 1.175343e-14, 1.184754e-14, 1.182505e-14, 1.185293e-14, 
    1.183871e-14, 1.186307e-14, 1.184114e-14, 1.187911e-14, 1.188737e-14, 
    1.188173e-14, 1.190341e-14, 1.183993e-14, 1.186432e-14, 1.168033e-14, 
    1.168141e-14, 1.168647e-14, 1.166422e-14, 1.166286e-14, 1.164247e-14, 
    1.166062e-14, 1.166834e-14, 1.168795e-14, 1.169954e-14, 1.171055e-14, 
    1.173474e-14, 1.176173e-14, 1.179944e-14, 1.182651e-14, 1.184463e-14, 
    1.183352e-14, 1.184333e-14, 1.183237e-14, 1.182722e-14, 1.188427e-14, 
    1.185225e-14, 1.190029e-14, 1.189763e-14, 1.18759e-14, 1.189793e-14, 
    1.168217e-14, 1.167593e-14, 1.165422e-14, 1.167121e-14, 1.164025e-14, 
    1.165758e-14, 1.166754e-14, 1.170594e-14, 1.171438e-14, 1.172219e-14, 
    1.173762e-14, 1.175741e-14, 1.179209e-14, 1.182223e-14, 1.184972e-14, 
    1.184771e-14, 1.184842e-14, 1.185455e-14, 1.183935e-14, 1.185705e-14, 
    1.186001e-14, 1.185225e-14, 1.189728e-14, 1.188442e-14, 1.189758e-14, 
    1.188921e-14, 1.167796e-14, 1.168847e-14, 1.168279e-14, 1.169347e-14, 
    1.168594e-14, 1.171937e-14, 1.172939e-14, 1.177622e-14, 1.175702e-14, 
    1.178758e-14, 1.176013e-14, 1.176499e-14, 1.178856e-14, 1.176161e-14, 
    1.182056e-14, 1.17806e-14, 1.185479e-14, 1.181492e-14, 1.185729e-14, 
    1.18496e-14, 1.186233e-14, 1.187371e-14, 1.188804e-14, 1.191444e-14, 
    1.190833e-14, 1.193039e-14, 1.170413e-14, 1.171775e-14, 1.171656e-14, 
    1.17308e-14, 1.174133e-14, 1.176415e-14, 1.180071e-14, 1.178697e-14, 
    1.181219e-14, 1.181725e-14, 1.177893e-14, 1.180246e-14, 1.172686e-14, 
    1.173908e-14, 1.173181e-14, 1.17052e-14, 1.179013e-14, 1.174657e-14, 
    1.182695e-14, 1.18034e-14, 1.187209e-14, 1.183794e-14, 1.190496e-14, 
    1.193354e-14, 1.196044e-14, 1.199181e-14, 1.172518e-14, 1.171593e-14, 
    1.17325e-14, 1.175539e-14, 1.177663e-14, 1.180484e-14, 1.180772e-14, 
    1.1813e-14, 1.182668e-14, 1.183816e-14, 1.181466e-14, 1.184104e-14, 
    1.174191e-14, 1.179391e-14, 1.171243e-14, 1.173698e-14, 1.175404e-14, 
    1.174657e-14, 1.17854e-14, 1.179454e-14, 1.183166e-14, 1.181248e-14, 
    1.192649e-14, 1.187611e-14, 1.201569e-14, 1.197676e-14, 1.17127e-14, 
    1.172515e-14, 1.176845e-14, 1.174786e-14, 1.180672e-14, 1.182119e-14, 
    1.183295e-14, 1.184796e-14, 1.184959e-14, 1.185848e-14, 1.184391e-14, 
    1.185791e-14, 1.180489e-14, 1.18286e-14, 1.176351e-14, 1.177936e-14, 
    1.177207e-14, 1.176407e-14, 1.178876e-14, 1.181503e-14, 1.18156e-14, 
    1.182402e-14, 1.184771e-14, 1.180696e-14, 1.193296e-14, 1.18552e-14, 
    1.173873e-14, 1.176268e-14, 1.176611e-14, 1.175683e-14, 1.181974e-14, 
    1.179696e-14, 1.185827e-14, 1.184171e-14, 1.186883e-14, 1.185536e-14, 
    1.185337e-14, 1.183606e-14, 1.182527e-14, 1.1798e-14, 1.17758e-14, 
    1.175818e-14, 1.176228e-14, 1.178163e-14, 1.181664e-14, 1.184973e-14, 
    1.184248e-14, 1.186677e-14, 1.180246e-14, 1.182944e-14, 1.181901e-14, 
    1.18462e-14, 1.17866e-14, 1.183733e-14, 1.177362e-14, 1.177921e-14, 
    1.179651e-14, 1.183126e-14, 1.183896e-14, 1.184716e-14, 1.18421e-14, 
    1.181753e-14, 1.181351e-14, 1.179609e-14, 1.179127e-14, 1.177799e-14, 
    1.176699e-14, 1.177704e-14, 1.178759e-14, 1.181755e-14, 1.184451e-14, 
    1.187387e-14, 1.188106e-14, 1.19153e-14, 1.188741e-14, 1.193339e-14, 
    1.189429e-14, 1.196196e-14, 1.184028e-14, 1.189316e-14, 1.17973e-14, 
    1.180764e-14, 1.182634e-14, 1.186918e-14, 1.184607e-14, 1.18731e-14, 
    1.181335e-14, 1.178229e-14, 1.177426e-14, 1.175925e-14, 1.17746e-14, 
    1.177335e-14, 1.178804e-14, 1.178332e-14, 1.181854e-14, 1.179963e-14, 
    1.185332e-14, 1.187289e-14, 1.192808e-14, 1.196185e-14, 1.19962e-14, 
    1.201134e-14, 1.201595e-14, 1.201787e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.152213e-11, -8.188185e-11, -8.181192e-11, -8.210205e-11, -8.194111e-11, 
    -8.213109e-11, -8.159506e-11, -8.189612e-11, -8.170394e-11, 
    -8.155453e-11, -8.266511e-11, -8.2115e-11, -8.323666e-11, -8.288577e-11, 
    -8.376728e-11, -8.318205e-11, -8.388529e-11, -8.375042e-11, 
    -8.415642e-11, -8.404011e-11, -8.45594e-11, -8.421011e-11, -8.482864e-11, 
    -8.4476e-11, -8.453115e-11, -8.419859e-11, -8.222572e-11, -8.259662e-11, 
    -8.220374e-11, -8.225663e-11, -8.22329e-11, -8.194444e-11, -8.179905e-11, 
    -8.149465e-11, -8.154992e-11, -8.17735e-11, -8.228041e-11, -8.210835e-11, 
    -8.254204e-11, -8.253224e-11, -8.301509e-11, -8.279739e-11, 
    -8.360901e-11, -8.337833e-11, -8.404497e-11, -8.387731e-11, 
    -8.403709e-11, -8.398864e-11, -8.403772e-11, -8.379183e-11, 
    -8.389717e-11, -8.368082e-11, -8.283815e-11, -8.308579e-11, 
    -8.234723e-11, -8.190316e-11, -8.160827e-11, -8.1399e-11, -8.142858e-11, 
    -8.148498e-11, -8.177481e-11, -8.204733e-11, -8.225502e-11, 
    -8.239395e-11, -8.253084e-11, -8.294516e-11, -8.316452e-11, 
    -8.365564e-11, -8.356703e-11, -8.371717e-11, -8.386063e-11, 
    -8.410147e-11, -8.406183e-11, -8.416794e-11, -8.371322e-11, 
    -8.401541e-11, -8.351654e-11, -8.365298e-11, -8.256799e-11, 
    -8.215477e-11, -8.197908e-11, -8.182536e-11, -8.145132e-11, 
    -8.170962e-11, -8.16078e-11, -8.185005e-11, -8.200399e-11, -8.192786e-11, 
    -8.239775e-11, -8.221506e-11, -8.317751e-11, -8.276294e-11, 
    -8.384389e-11, -8.358522e-11, -8.39059e-11, -8.374226e-11, -8.402264e-11, 
    -8.37703e-11, -8.420743e-11, -8.430261e-11, -8.423757e-11, -8.448745e-11, 
    -8.375631e-11, -8.403708e-11, -8.192572e-11, -8.193814e-11, 
    -8.199599e-11, -8.17417e-11, -8.172614e-11, -8.149313e-11, -8.170047e-11, 
    -8.178876e-11, -8.201292e-11, -8.21455e-11, -8.227154e-11, -8.254866e-11, 
    -8.285816e-11, -8.3291e-11, -8.360198e-11, -8.381044e-11, -8.368262e-11, 
    -8.379547e-11, -8.366931e-11, -8.36102e-11, -8.426694e-11, -8.389816e-11, 
    -8.445151e-11, -8.442089e-11, -8.417046e-11, -8.442434e-11, 
    -8.194686e-11, -8.187541e-11, -8.162732e-11, -8.182147e-11, 
    -8.146776e-11, -8.166574e-11, -8.177958e-11, -8.221886e-11, -8.23154e-11, 
    -8.24049e-11, -8.258166e-11, -8.280852e-11, -8.320651e-11, -8.355282e-11, 
    -8.386897e-11, -8.384581e-11, -8.385397e-11, -8.392459e-11, 
    -8.374965e-11, -8.395331e-11, -8.398748e-11, -8.389812e-11, 
    -8.441679e-11, -8.426861e-11, -8.442024e-11, -8.432376e-11, 
    -8.189863e-11, -8.201886e-11, -8.19539e-11, -8.207606e-11, -8.198999e-11, 
    -8.23727e-11, -8.248745e-11, -8.302442e-11, -8.280406e-11, -8.31548e-11, 
    -8.283969e-11, -8.289552e-11, -8.316621e-11, -8.285672e-11, 
    -8.353371e-11, -8.307471e-11, -8.392733e-11, -8.346892e-11, 
    -8.395606e-11, -8.386761e-11, -8.401406e-11, -8.414523e-11, 
    -8.431025e-11, -8.461474e-11, -8.454423e-11, -8.479888e-11, -8.21981e-11, 
    -8.235405e-11, -8.234033e-11, -8.250353e-11, -8.262423e-11, 
    -8.288587e-11, -8.33055e-11, -8.31477e-11, -8.343741e-11, -8.349556e-11, 
    -8.305544e-11, -8.332566e-11, -8.245842e-11, -8.259852e-11, 
    -8.251511e-11, -8.221041e-11, -8.318405e-11, -8.268435e-11, 
    -8.360712e-11, -8.33364e-11, -8.412652e-11, -8.373355e-11, -8.450542e-11, 
    -8.483537e-11, -8.514598e-11, -8.550892e-11, -8.243917e-11, 
    -8.233321e-11, -8.252295e-11, -8.278545e-11, -8.302906e-11, 
    -8.335291e-11, -8.338605e-11, -8.344672e-11, -8.360389e-11, 
    -8.373603e-11, -8.346589e-11, -8.376915e-11, -8.263099e-11, 
    -8.322742e-11, -8.229314e-11, -8.257444e-11, -8.276999e-11, 
    -8.268421e-11, -8.312967e-11, -8.323466e-11, -8.366131e-11, 
    -8.344075e-11, -8.475393e-11, -8.417292e-11, -8.578532e-11, 
    -8.533468e-11, -8.229618e-11, -8.243881e-11, -8.293521e-11, 
    -8.269902e-11, -8.337454e-11, -8.354081e-11, -8.3676e-11, -8.38488e-11, 
    -8.386746e-11, -8.396984e-11, -8.380207e-11, -8.396322e-11, 
    -8.335359e-11, -8.362602e-11, -8.287848e-11, -8.306041e-11, 
    -8.297672e-11, -8.288491e-11, -8.316827e-11, -8.347014e-11, 
    -8.347661e-11, -8.357341e-11, -8.384615e-11, -8.337727e-11, 
    -8.482888e-11, -8.393234e-11, -8.259434e-11, -8.286905e-11, 
    -8.290831e-11, -8.280189e-11, -8.352415e-11, -8.326244e-11, 
    -8.396735e-11, -8.377683e-11, -8.4089e-11, -8.393387e-11, -8.391105e-11, 
    -8.371183e-11, -8.358779e-11, -8.327443e-11, -8.301948e-11, 
    -8.281733e-11, -8.286434e-11, -8.30864e-11, -8.348861e-11, -8.386914e-11, 
    -8.378578e-11, -8.406528e-11, -8.332555e-11, -8.363572e-11, 
    -8.351583e-11, -8.382843e-11, -8.314351e-11, -8.37267e-11, -8.299444e-11, 
    -8.305864e-11, -8.325724e-11, -8.365674e-11, -8.374516e-11, 
    -8.383953e-11, -8.378129e-11, -8.349883e-11, -8.345256e-11, 
    -8.325242e-11, -8.319715e-11, -8.304466e-11, -8.291841e-11, 
    -8.303376e-11, -8.315489e-11, -8.349895e-11, -8.380902e-11, 
    -8.414709e-11, -8.422983e-11, -8.462481e-11, -8.430326e-11, 
    -8.483387e-11, -8.438272e-11, -8.516374e-11, -8.376053e-11, 
    -8.436948e-11, -8.326628e-11, -8.338513e-11, -8.360008e-11, 
    -8.409313e-11, -8.382697e-11, -8.413825e-11, -8.345075e-11, 
    -8.309405e-11, -8.300179e-11, -8.282962e-11, -8.300573e-11, 
    -8.299141e-11, -8.315992e-11, -8.310577e-11, -8.351038e-11, 
    -8.329304e-11, -8.391048e-11, -8.41358e-11, -8.477219e-11, -8.516234e-11, 
    -8.555952e-11, -8.573487e-11, -8.578824e-11, -8.581056e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -1.964839e-12, -1.973507e-12, -1.971822e-12, -1.978813e-12, -1.974935e-12, 
    -1.979513e-12, -1.966597e-12, -1.973851e-12, -1.96922e-12, -1.96562e-12, 
    -1.992381e-12, -1.979125e-12, -2.006153e-12, -1.997698e-12, -2.01894e-12, 
    -2.004838e-12, -2.021783e-12, -2.018533e-12, -2.028317e-12, 
    -2.025514e-12, -2.038027e-12, -2.02961e-12, -2.044515e-12, -2.036017e-12, 
    -2.037346e-12, -2.029333e-12, -1.981793e-12, -1.99073e-12, -1.981264e-12, 
    -1.982538e-12, -1.981966e-12, -1.975015e-12, -1.971512e-12, 
    -1.964177e-12, -1.965509e-12, -1.970896e-12, -1.983111e-12, 
    -1.978965e-12, -1.989416e-12, -1.98918e-12, -2.000814e-12, -1.995568e-12, 
    -2.015126e-12, -2.009567e-12, -2.025631e-12, -2.021591e-12, 
    -2.025441e-12, -2.024274e-12, -2.025456e-12, -2.019531e-12, -2.02207e-12, 
    -2.016856e-12, -1.996551e-12, -2.002518e-12, -1.984721e-12, 
    -1.974021e-12, -1.966915e-12, -1.961872e-12, -1.962585e-12, 
    -1.963944e-12, -1.970928e-12, -1.977495e-12, -1.982499e-12, 
    -1.985847e-12, -1.989146e-12, -1.99913e-12, -2.004415e-12, -2.01625e-12, 
    -2.014114e-12, -2.017732e-12, -2.021189e-12, -2.026992e-12, 
    -2.026037e-12, -2.028594e-12, -2.017637e-12, -2.024919e-12, 
    -2.012898e-12, -2.016185e-12, -1.990041e-12, -1.980084e-12, -1.97585e-12, 
    -1.972146e-12, -1.963133e-12, -1.969357e-12, -1.966903e-12, 
    -1.972741e-12, -1.97645e-12, -1.974616e-12, -1.985939e-12, -1.981536e-12, 
    -2.004728e-12, -1.994738e-12, -2.020786e-12, -2.014553e-12, -2.02228e-12, 
    -2.018337e-12, -2.025093e-12, -2.019013e-12, -2.029546e-12, 
    -2.031839e-12, -2.030272e-12, -2.036293e-12, -2.018675e-12, 
    -2.025441e-12, -1.974564e-12, -1.974863e-12, -1.976257e-12, -1.97013e-12, 
    -1.969755e-12, -1.96414e-12, -1.969136e-12, -1.971264e-12, -1.976665e-12, 
    -1.97986e-12, -1.982897e-12, -1.989575e-12, -1.997033e-12, -2.007463e-12, 
    -2.014957e-12, -2.01998e-12, -2.0169e-12, -2.019619e-12, -2.016579e-12, 
    -2.015154e-12, -2.03098e-12, -2.022093e-12, -2.035427e-12, -2.034689e-12, 
    -2.028655e-12, -2.034773e-12, -1.975074e-12, -1.973352e-12, 
    -1.967374e-12, -1.972052e-12, -1.963529e-12, -1.9683e-12, -1.971043e-12, 
    -1.981628e-12, -1.983954e-12, -1.986111e-12, -1.99037e-12, -1.995837e-12, 
    -2.005427e-12, -2.013772e-12, -2.02139e-12, -2.020832e-12, -2.021029e-12, 
    -2.02273e-12, -2.018515e-12, -2.023422e-12, -2.024246e-12, -2.022092e-12, 
    -2.034591e-12, -2.03102e-12, -2.034674e-12, -2.032349e-12, -1.973911e-12, 
    -1.976809e-12, -1.975243e-12, -1.978187e-12, -1.976113e-12, 
    -1.985335e-12, -1.9881e-12, -2.001039e-12, -1.995729e-12, -2.004181e-12, 
    -1.996588e-12, -1.997933e-12, -2.004456e-12, -1.996998e-12, 
    -2.013311e-12, -2.002251e-12, -2.022796e-12, -2.01175e-12, -2.023489e-12, 
    -2.021357e-12, -2.024886e-12, -2.028047e-12, -2.032023e-12, -2.03936e-12, 
    -2.037661e-12, -2.043798e-12, -1.981128e-12, -1.984886e-12, 
    -1.984555e-12, -1.988488e-12, -1.991396e-12, -1.997701e-12, 
    -2.007812e-12, -2.00401e-12, -2.010991e-12, -2.012392e-12, -2.001787e-12, 
    -2.008298e-12, -1.987401e-12, -1.990776e-12, -1.988767e-12, 
    -1.981424e-12, -2.004886e-12, -1.992845e-12, -2.01508e-12, -2.008557e-12, 
    -2.027596e-12, -2.018127e-12, -2.036726e-12, -2.044677e-12, 
    -2.052161e-12, -2.060907e-12, -1.986937e-12, -1.984383e-12, 
    -1.988955e-12, -1.995281e-12, -2.001151e-12, -2.008955e-12, 
    -2.009753e-12, -2.011215e-12, -2.015002e-12, -2.018187e-12, 
    -2.011677e-12, -2.018985e-12, -1.991559e-12, -2.005931e-12, 
    -1.983418e-12, -1.990196e-12, -1.994908e-12, -1.992841e-12, 
    -2.003575e-12, -2.006105e-12, -2.016386e-12, -2.011072e-12, 
    -2.042714e-12, -2.028714e-12, -2.067567e-12, -2.056708e-12, 
    -1.983491e-12, -1.986928e-12, -1.99889e-12, -1.993198e-12, -2.009476e-12, 
    -2.013482e-12, -2.01674e-12, -2.020904e-12, -2.021354e-12, -2.023821e-12, 
    -2.019778e-12, -2.023661e-12, -2.008971e-12, -2.015536e-12, 
    -1.997523e-12, -2.001907e-12, -1.99989e-12, -1.997678e-12, -2.004506e-12, 
    -2.01178e-12, -2.011936e-12, -2.014268e-12, -2.02084e-12, -2.009542e-12, 
    -2.04452e-12, -2.022917e-12, -1.990676e-12, -1.997295e-12, -1.998241e-12, 
    -1.995677e-12, -2.013081e-12, -2.006775e-12, -2.023761e-12, -2.01917e-12, 
    -2.026692e-12, -2.022954e-12, -2.022404e-12, -2.017604e-12, 
    -2.014615e-12, -2.007064e-12, -2.00092e-12, -1.996049e-12, -1.997182e-12, 
    -2.002533e-12, -2.012225e-12, -2.021394e-12, -2.019386e-12, -2.02612e-12, 
    -2.008295e-12, -2.015769e-12, -2.012881e-12, -2.020413e-12, 
    -2.003909e-12, -2.017962e-12, -2.000317e-12, -2.001864e-12, 
    -2.006649e-12, -2.016276e-12, -2.018406e-12, -2.02068e-12, -2.019277e-12, 
    -2.012471e-12, -2.011356e-12, -2.006533e-12, -2.005202e-12, 
    -2.001527e-12, -1.998485e-12, -2.001264e-12, -2.004183e-12, 
    -2.012474e-12, -2.019945e-12, -2.028092e-12, -2.030086e-12, 
    -2.039603e-12, -2.031855e-12, -2.044641e-12, -2.033769e-12, 
    -2.052589e-12, -2.018777e-12, -2.03345e-12, -2.006867e-12, -2.009731e-12, 
    -2.014911e-12, -2.026791e-12, -2.020378e-12, -2.027879e-12, 
    -2.011312e-12, -2.002717e-12, -2.000494e-12, -1.996345e-12, 
    -2.000589e-12, -2.000244e-12, -2.004304e-12, -2.003e-12, -2.012749e-12, 
    -2.007512e-12, -2.02239e-12, -2.02782e-12, -2.043154e-12, -2.052555e-12, 
    -2.062126e-12, -2.066351e-12, -2.067638e-12, -2.068175e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.782927e-15, 3.793152e-15, 3.791166e-15, 3.799406e-15, 3.794837e-15, 
    3.80023e-15, 3.785003e-15, 3.793557e-15, 3.788098e-15, 3.78385e-15, 
    3.815371e-15, 3.799773e-15, 3.831558e-15, 3.821628e-15, 3.846554e-15, 
    3.830012e-15, 3.849887e-15, 3.846081e-15, 3.857539e-15, 3.854258e-15, 
    3.868892e-15, 3.859053e-15, 3.876472e-15, 3.866544e-15, 3.868097e-15, 
    3.858728e-15, 3.802917e-15, 3.81343e-15, 3.802294e-15, 3.803793e-15, 
    3.803121e-15, 3.79493e-15, 3.790798e-15, 3.782147e-15, 3.783719e-15, 
    3.790073e-15, 3.804468e-15, 3.799586e-15, 3.811891e-15, 3.811613e-15, 
    3.825291e-15, 3.819126e-15, 3.842086e-15, 3.835567e-15, 3.854395e-15, 
    3.849664e-15, 3.854173e-15, 3.852806e-15, 3.85419e-15, 3.84725e-15, 
    3.850224e-15, 3.844115e-15, 3.82028e-15, 3.827291e-15, 3.806364e-15, 
    3.793755e-15, 3.785378e-15, 3.779426e-15, 3.780267e-15, 3.781871e-15, 
    3.790111e-15, 3.797854e-15, 3.80375e-15, 3.807691e-15, 3.811573e-15, 
    3.823306e-15, 3.829517e-15, 3.843403e-15, 3.840901e-15, 3.845141e-15, 
    3.849193e-15, 3.855988e-15, 3.854871e-15, 3.857863e-15, 3.845031e-15, 
    3.85356e-15, 3.839475e-15, 3.843329e-15, 3.812618e-15, 3.800904e-15, 
    3.795912e-15, 3.791548e-15, 3.780915e-15, 3.788258e-15, 3.785364e-15, 
    3.792251e-15, 3.796623e-15, 3.794461e-15, 3.807798e-15, 3.802615e-15, 
    3.829885e-15, 3.818149e-15, 3.84872e-15, 3.841415e-15, 3.850471e-15, 
    3.845851e-15, 3.853764e-15, 3.846643e-15, 3.858977e-15, 3.861659e-15, 
    3.859826e-15, 3.866869e-15, 3.846248e-15, 3.854171e-15, 3.7944e-15, 
    3.794752e-15, 3.796396e-15, 3.78917e-15, 3.788728e-15, 3.782104e-15, 
    3.787999e-15, 3.790508e-15, 3.796877e-15, 3.800641e-15, 3.804218e-15, 
    3.812077e-15, 3.820846e-15, 3.833096e-15, 3.841888e-15, 3.847777e-15, 
    3.844167e-15, 3.847354e-15, 3.843791e-15, 3.842121e-15, 3.860654e-15, 
    3.850251e-15, 3.865856e-15, 3.864994e-15, 3.857934e-15, 3.865091e-15, 
    3.795e-15, 3.792971e-15, 3.78592e-15, 3.791438e-15, 3.781382e-15, 
    3.787011e-15, 3.790246e-15, 3.802721e-15, 3.805462e-15, 3.808001e-15, 
    3.813013e-15, 3.819441e-15, 3.830707e-15, 3.840498e-15, 3.849429e-15, 
    3.848775e-15, 3.849005e-15, 3.850998e-15, 3.846059e-15, 3.851809e-15, 
    3.852773e-15, 3.850251e-15, 3.864878e-15, 3.860702e-15, 3.864975e-15, 
    3.862257e-15, 3.793631e-15, 3.797045e-15, 3.795201e-15, 3.798669e-15, 
    3.796225e-15, 3.807085e-15, 3.810339e-15, 3.825552e-15, 3.819314e-15, 
    3.829243e-15, 3.820324e-15, 3.821905e-15, 3.829562e-15, 3.820807e-15, 
    3.839957e-15, 3.826974e-15, 3.851076e-15, 3.838124e-15, 3.851887e-15, 
    3.84939e-15, 3.853523e-15, 3.857222e-15, 3.861876e-15, 3.870452e-15, 
    3.868467e-15, 3.875637e-15, 3.802134e-15, 3.806558e-15, 3.80617e-15, 
    3.810798e-15, 3.814219e-15, 3.821632e-15, 3.833507e-15, 3.829044e-15, 
    3.837238e-15, 3.838881e-15, 3.826434e-15, 3.834076e-15, 3.809518e-15, 
    3.813488e-15, 3.811126e-15, 3.802482e-15, 3.83007e-15, 3.815921e-15, 
    3.842033e-15, 3.834381e-15, 3.856695e-15, 3.845603e-15, 3.867374e-15, 
    3.876659e-15, 3.885398e-15, 3.895588e-15, 3.808973e-15, 3.805968e-15, 
    3.811349e-15, 3.818786e-15, 3.825686e-15, 3.834848e-15, 3.835786e-15, 
    3.837501e-15, 3.841943e-15, 3.845675e-15, 3.838041e-15, 3.846611e-15, 
    3.814405e-15, 3.831298e-15, 3.80483e-15, 3.812805e-15, 3.818348e-15, 
    3.815919e-15, 3.828534e-15, 3.831504e-15, 3.843563e-15, 3.837332e-15, 
    3.874367e-15, 3.858001e-15, 3.903345e-15, 3.890697e-15, 3.804917e-15, 
    3.808963e-15, 3.823028e-15, 3.816339e-15, 3.83546e-15, 3.84016e-15, 
    3.84398e-15, 3.848858e-15, 3.849386e-15, 3.852275e-15, 3.84754e-15, 
    3.852089e-15, 3.834867e-15, 3.842568e-15, 3.821424e-15, 3.826573e-15, 
    3.824206e-15, 3.821606e-15, 3.829627e-15, 3.83816e-15, 3.838346e-15, 
    3.84108e-15, 3.848775e-15, 3.835538e-15, 3.876471e-15, 3.851209e-15, 
    3.813373e-15, 3.821153e-15, 3.822268e-15, 3.819254e-15, 3.839688e-15, 
    3.83229e-15, 3.852205e-15, 3.846828e-15, 3.855638e-15, 3.851261e-15, 
    3.850616e-15, 3.844992e-15, 3.841488e-15, 3.832628e-15, 3.825415e-15, 
    3.819692e-15, 3.821023e-15, 3.827308e-15, 3.838683e-15, 3.849432e-15, 
    3.847078e-15, 3.854968e-15, 3.834075e-15, 3.84284e-15, 3.839453e-15, 
    3.848284e-15, 3.828925e-15, 3.845403e-15, 3.824707e-15, 3.826524e-15, 
    3.832143e-15, 3.843432e-15, 3.845933e-15, 3.848596e-15, 3.846953e-15, 
    3.838972e-15, 3.837665e-15, 3.832007e-15, 3.830442e-15, 3.826129e-15, 
    3.822554e-15, 3.82582e-15, 3.829246e-15, 3.838977e-15, 3.847735e-15, 
    3.857275e-15, 3.859609e-15, 3.870731e-15, 3.861674e-15, 3.876611e-15, 
    3.863907e-15, 3.88589e-15, 3.846362e-15, 3.86354e-15, 3.832399e-15, 
    3.83576e-15, 3.841832e-15, 3.85575e-15, 3.848243e-15, 3.857024e-15, 
    3.837614e-15, 3.827524e-15, 3.824915e-15, 3.820039e-15, 3.825026e-15, 
    3.824621e-15, 3.82939e-15, 3.827858e-15, 3.8393e-15, 3.833156e-15, 
    3.850599e-15, 3.856955e-15, 3.874884e-15, 3.885855e-15, 3.897012e-15, 
    3.901931e-15, 3.903429e-15, 3.904054e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.535308e-09, -8.572939e-09, -8.565624e-09, -8.595976e-09, -8.579139e-09, 
    -8.599014e-09, -8.542937e-09, -8.574432e-09, -8.554327e-09, 
    -8.538696e-09, -8.65488e-09, -8.597331e-09, -8.714673e-09, -8.677964e-09, 
    -8.770182e-09, -8.708959e-09, -8.782528e-09, -8.768418e-09, 
    -8.810892e-09, -8.798724e-09, -8.853048e-09, -8.816508e-09, 
    -8.881213e-09, -8.844323e-09, -8.850092e-09, -8.815302e-09, 
    -8.608914e-09, -8.647715e-09, -8.606614e-09, -8.612147e-09, 
    -8.609665e-09, -8.579486e-09, -8.564277e-09, -8.532433e-09, 
    -8.538214e-09, -8.561604e-09, -8.614635e-09, -8.596635e-09, 
    -8.642005e-09, -8.64098e-09, -8.691494e-09, -8.668718e-09, -8.753624e-09, 
    -8.729493e-09, -8.799232e-09, -8.781692e-09, -8.798407e-09, 
    -8.793339e-09, -8.798473e-09, -8.772751e-09, -8.783771e-09, 
    -8.761137e-09, -8.672983e-09, -8.698889e-09, -8.621626e-09, 
    -8.575169e-09, -8.544318e-09, -8.522425e-09, -8.525521e-09, -8.53142e-09, 
    -8.561742e-09, -8.590251e-09, -8.611979e-09, -8.626513e-09, 
    -8.640834e-09, -8.684178e-09, -8.707125e-09, -8.758503e-09, 
    -8.749232e-09, -8.76494e-09, -8.779947e-09, -8.805142e-09, -8.800995e-09, 
    -8.812096e-09, -8.764526e-09, -8.79614e-09, -8.743951e-09, -8.758225e-09, 
    -8.64472e-09, -8.601491e-09, -8.583112e-09, -8.56703e-09, -8.5279e-09, 
    -8.554921e-09, -8.544269e-09, -8.569613e-09, -8.585717e-09, 
    -8.577753e-09, -8.62691e-09, -8.607798e-09, -8.708485e-09, -8.665114e-09, 
    -8.778197e-09, -8.751136e-09, -8.784683e-09, -8.767565e-09, 
    -8.796896e-09, -8.770498e-09, -8.816228e-09, -8.826184e-09, -8.81938e-09, 
    -8.845521e-09, -8.769035e-09, -8.798406e-09, -8.577529e-09, 
    -8.578828e-09, -8.584879e-09, -8.558277e-09, -8.55665e-09, -8.532274e-09, 
    -8.553965e-09, -8.563201e-09, -8.586651e-09, -8.600521e-09, 
    -8.613706e-09, -8.642698e-09, -8.675077e-09, -8.720356e-09, -8.75289e-09, 
    -8.774697e-09, -8.761326e-09, -8.773132e-09, -8.759934e-09, 
    -8.753749e-09, -8.822453e-09, -8.783873e-09, -8.841761e-09, 
    -8.838558e-09, -8.81236e-09, -8.838919e-09, -8.57974e-09, -8.572266e-09, 
    -8.546312e-09, -8.566623e-09, -8.529619e-09, -8.550331e-09, -8.56224e-09, 
    -8.608196e-09, -8.618295e-09, -8.627658e-09, -8.64615e-09, -8.669883e-09, 
    -8.711518e-09, -8.747747e-09, -8.780821e-09, -8.778398e-09, -8.77925e-09, 
    -8.786638e-09, -8.768337e-09, -8.789643e-09, -8.793219e-09, -8.78387e-09, 
    -8.838128e-09, -8.822627e-09, -8.83849e-09, -8.828397e-09, -8.574696e-09, 
    -8.587273e-09, -8.580477e-09, -8.593257e-09, -8.584252e-09, -8.62429e-09, 
    -8.636294e-09, -8.692469e-09, -8.669416e-09, -8.706108e-09, 
    -8.673144e-09, -8.678985e-09, -8.707302e-09, -8.674926e-09, 
    -8.745747e-09, -8.69773e-09, -8.786926e-09, -8.73897e-09, -8.789931e-09, 
    -8.780678e-09, -8.795999e-09, -8.80972e-09, -8.826984e-09, -8.858836e-09, 
    -8.851461e-09, -8.878101e-09, -8.606024e-09, -8.622338e-09, 
    -8.620903e-09, -8.637977e-09, -8.650604e-09, -8.677975e-09, 
    -8.721874e-09, -8.705366e-09, -8.735674e-09, -8.741758e-09, 
    -8.695713e-09, -8.723982e-09, -8.633258e-09, -8.647913e-09, 
    -8.639188e-09, -8.607311e-09, -8.709168e-09, -8.656892e-09, 
    -8.753427e-09, -8.725106e-09, -8.807763e-09, -8.766654e-09, -8.8474e-09, 
    -8.881917e-09, -8.914411e-09, -8.952378e-09, -8.631243e-09, 
    -8.620158e-09, -8.640008e-09, -8.667469e-09, -8.692954e-09, 
    -8.726833e-09, -8.7303e-09, -8.736647e-09, -8.753089e-09, -8.766913e-09, 
    -8.738653e-09, -8.770378e-09, -8.651311e-09, -8.713706e-09, 
    -8.615967e-09, -8.645395e-09, -8.665851e-09, -8.656879e-09, -8.70348e-09, 
    -8.714463e-09, -8.759096e-09, -8.736023e-09, -8.873397e-09, 
    -8.812616e-09, -8.981292e-09, -8.93415e-09, -8.616285e-09, -8.631206e-09, 
    -8.683136e-09, -8.658428e-09, -8.729096e-09, -8.746491e-09, 
    -8.760633e-09, -8.778709e-09, -8.780662e-09, -8.791373e-09, 
    -8.773822e-09, -8.79068e-09, -8.726905e-09, -8.755404e-09, -8.677202e-09, 
    -8.696235e-09, -8.687479e-09, -8.677874e-09, -8.707517e-09, 
    -8.739097e-09, -8.739774e-09, -8.7499e-09, -8.778432e-09, -8.729383e-09, 
    -8.881239e-09, -8.78745e-09, -8.647477e-09, -8.676215e-09, -8.680323e-09, 
    -8.66919e-09, -8.744746e-09, -8.717369e-09, -8.791112e-09, -8.771182e-09, 
    -8.803838e-09, -8.787611e-09, -8.785222e-09, -8.764381e-09, 
    -8.751405e-09, -8.718624e-09, -8.691952e-09, -8.670805e-09, 
    -8.675722e-09, -8.698953e-09, -8.74103e-09, -8.780838e-09, -8.772117e-09, 
    -8.801356e-09, -8.723972e-09, -8.756419e-09, -8.743877e-09, 
    -8.776579e-09, -8.704927e-09, -8.765936e-09, -8.689332e-09, 
    -8.696049e-09, -8.716825e-09, -8.758618e-09, -8.767867e-09, -8.77774e-09, 
    -8.771648e-09, -8.742099e-09, -8.737258e-09, -8.716321e-09, 
    -8.710539e-09, -8.694586e-09, -8.681379e-09, -8.693446e-09, 
    -8.706118e-09, -8.742111e-09, -8.774548e-09, -8.809915e-09, 
    -8.818571e-09, -8.859891e-09, -8.826252e-09, -8.881761e-09, 
    -8.834564e-09, -8.916268e-09, -8.769476e-09, -8.83318e-09, -8.717771e-09, 
    -8.730204e-09, -8.75269e-09, -8.80427e-09, -8.776426e-09, -8.808991e-09, 
    -8.737068e-09, -8.699754e-09, -8.690101e-09, -8.67209e-09, -8.690513e-09, 
    -8.689015e-09, -8.706644e-09, -8.700979e-09, -8.743307e-09, -8.72057e-09, 
    -8.785162e-09, -8.808734e-09, -8.875308e-09, -8.916121e-09, 
    -8.957672e-09, -8.976015e-09, -8.981599e-09, -8.983933e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.012876e-10, -1.017343e-10, -1.016474e-10, -1.020078e-10, -1.018079e-10, 
    -1.020438e-10, -1.013781e-10, -1.01752e-10, -1.015133e-10, -1.013278e-10, 
    -1.02707e-10, -1.020238e-10, -1.034169e-10, -1.029811e-10, -1.040759e-10, 
    -1.033491e-10, -1.042225e-10, -1.040549e-10, -1.045592e-10, 
    -1.044147e-10, -1.050597e-10, -1.046259e-10, -1.053941e-10, 
    -1.049561e-10, -1.050246e-10, -1.046115e-10, -1.021614e-10, -1.02622e-10, 
    -1.021341e-10, -1.021997e-10, -1.021703e-10, -1.01812e-10, -1.016315e-10, 
    -1.012534e-10, -1.013221e-10, -1.015997e-10, -1.022293e-10, 
    -1.020156e-10, -1.025542e-10, -1.02542e-10, -1.031417e-10, -1.028713e-10, 
    -1.038793e-10, -1.035928e-10, -1.044207e-10, -1.042125e-10, -1.04411e-10, 
    -1.043508e-10, -1.044118e-10, -1.041064e-10, -1.042372e-10, 
    -1.039685e-10, -1.02922e-10, -1.032295e-10, -1.023123e-10, -1.017608e-10, 
    -1.013945e-10, -1.011346e-10, -1.011714e-10, -1.012414e-10, 
    -1.016014e-10, -1.019398e-10, -1.021977e-10, -1.023703e-10, 
    -1.025403e-10, -1.030549e-10, -1.033273e-10, -1.039372e-10, 
    -1.038272e-10, -1.040136e-10, -1.041918e-10, -1.044909e-10, 
    -1.044417e-10, -1.045735e-10, -1.040087e-10, -1.043841e-10, 
    -1.037645e-10, -1.039339e-10, -1.025864e-10, -1.020732e-10, 
    -1.018551e-10, -1.016641e-10, -1.011996e-10, -1.015204e-10, 
    -1.013939e-10, -1.016948e-10, -1.01886e-10, -1.017914e-10, -1.02375e-10, 
    -1.021481e-10, -1.033434e-10, -1.028285e-10, -1.04171e-10, -1.038498e-10, 
    -1.04248e-10, -1.040448e-10, -1.04393e-10, -1.040796e-10, -1.046225e-10, 
    -1.047407e-10, -1.0466e-10, -1.049703e-10, -1.040623e-10, -1.04411e-10, 
    -1.017888e-10, -1.018042e-10, -1.01876e-10, -1.015602e-10, -1.015409e-10, 
    -1.012515e-10, -1.01509e-10, -1.016187e-10, -1.018971e-10, -1.020617e-10, 
    -1.022182e-10, -1.025624e-10, -1.029468e-10, -1.034844e-10, 
    -1.038706e-10, -1.041295e-10, -1.039707e-10, -1.041109e-10, 
    -1.039542e-10, -1.038808e-10, -1.046964e-10, -1.042384e-10, 
    -1.049257e-10, -1.048876e-10, -1.045766e-10, -1.048919e-10, -1.01815e-10, 
    -1.017263e-10, -1.014182e-10, -1.016593e-10, -1.0122e-10, -1.014659e-10, 
    -1.016073e-10, -1.021528e-10, -1.022727e-10, -1.023839e-10, 
    -1.026034e-10, -1.028852e-10, -1.033794e-10, -1.038095e-10, 
    -1.042022e-10, -1.041734e-10, -1.041835e-10, -1.042712e-10, -1.04054e-10, 
    -1.043069e-10, -1.043494e-10, -1.042384e-10, -1.048825e-10, 
    -1.046985e-10, -1.048868e-10, -1.04767e-10, -1.017551e-10, -1.019045e-10, 
    -1.018238e-10, -1.019755e-10, -1.018686e-10, -1.023439e-10, 
    -1.024864e-10, -1.031533e-10, -1.028796e-10, -1.033152e-10, 
    -1.029239e-10, -1.029932e-10, -1.033294e-10, -1.02945e-10, -1.037858e-10, 
    -1.032157e-10, -1.042747e-10, -1.037053e-10, -1.043103e-10, 
    -1.042005e-10, -1.043824e-10, -1.045453e-10, -1.047502e-10, 
    -1.051284e-10, -1.050408e-10, -1.053571e-10, -1.021271e-10, 
    -1.023207e-10, -1.023037e-10, -1.025064e-10, -1.026563e-10, 
    -1.029812e-10, -1.035024e-10, -1.033064e-10, -1.036662e-10, 
    -1.037384e-10, -1.031918e-10, -1.035274e-10, -1.024504e-10, 
    -1.026243e-10, -1.025208e-10, -1.021423e-10, -1.033515e-10, 
    -1.027309e-10, -1.03877e-10, -1.035407e-10, -1.04522e-10, -1.04034e-10, 
    -1.049926e-10, -1.054024e-10, -1.057882e-10, -1.06239e-10, -1.024264e-10, 
    -1.022948e-10, -1.025305e-10, -1.028565e-10, -1.03159e-10, -1.035612e-10, 
    -1.036024e-10, -1.036778e-10, -1.038729e-10, -1.040371e-10, 
    -1.037016e-10, -1.040782e-10, -1.026647e-10, -1.034054e-10, 
    -1.022451e-10, -1.025944e-10, -1.028373e-10, -1.027308e-10, -1.03284e-10, 
    -1.034144e-10, -1.039443e-10, -1.036704e-10, -1.053013e-10, 
    -1.045797e-10, -1.065822e-10, -1.060226e-10, -1.022489e-10, -1.02426e-10, 
    -1.030425e-10, -1.027492e-10, -1.035881e-10, -1.037946e-10, 
    -1.039625e-10, -1.041771e-10, -1.042003e-10, -1.043275e-10, 
    -1.041191e-10, -1.043192e-10, -1.035621e-10, -1.039004e-10, -1.02972e-10, 
    -1.03198e-10, -1.03094e-10, -1.0298e-10, -1.033319e-10, -1.037068e-10, 
    -1.037149e-10, -1.038351e-10, -1.041738e-10, -1.035915e-10, 
    -1.053944e-10, -1.042809e-10, -1.026191e-10, -1.029603e-10, 
    -1.030091e-10, -1.028769e-10, -1.037739e-10, -1.034489e-10, 
    -1.043244e-10, -1.040877e-10, -1.044754e-10, -1.042828e-10, 
    -1.042544e-10, -1.04007e-10, -1.03853e-10, -1.034638e-10, -1.031472e-10, 
    -1.028961e-10, -1.029545e-10, -1.032303e-10, -1.037298e-10, 
    -1.042024e-10, -1.040989e-10, -1.04446e-10, -1.035273e-10, -1.039125e-10, 
    -1.037636e-10, -1.041518e-10, -1.033012e-10, -1.040255e-10, -1.03116e-10, 
    -1.031958e-10, -1.034424e-10, -1.039386e-10, -1.040484e-10, 
    -1.041656e-10, -1.040933e-10, -1.037425e-10, -1.03685e-10, -1.034364e-10, 
    -1.033678e-10, -1.031784e-10, -1.030216e-10, -1.031649e-10, 
    -1.033153e-10, -1.037426e-10, -1.041277e-10, -1.045476e-10, 
    -1.046504e-10, -1.051409e-10, -1.047415e-10, -1.054006e-10, 
    -1.048402e-10, -1.058102e-10, -1.040675e-10, -1.048238e-10, 
    -1.034537e-10, -1.036013e-10, -1.038682e-10, -1.044806e-10, -1.0415e-10, 
    -1.045366e-10, -1.036828e-10, -1.032398e-10, -1.031252e-10, 
    -1.029114e-10, -1.031301e-10, -1.031123e-10, -1.033216e-10, 
    -1.032543e-10, -1.037568e-10, -1.034869e-10, -1.042537e-10, 
    -1.045336e-10, -1.053239e-10, -1.058085e-10, -1.063018e-10, 
    -1.065196e-10, -1.065859e-10, -1.066136e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.400407e-12, -8.437474e-12, -8.430269e-12, -8.460165e-12, -8.443581e-12, 
    -8.463157e-12, -8.407923e-12, -8.438944e-12, -8.419141e-12, 
    -8.403745e-12, -8.518184e-12, -8.461499e-12, -8.57708e-12, -8.540922e-12, 
    -8.631758e-12, -8.571453e-12, -8.643918e-12, -8.630019e-12, 
    -8.671857e-12, -8.659871e-12, -8.713382e-12, -8.677389e-12, 
    -8.741124e-12, -8.704787e-12, -8.71047e-12, -8.676201e-12, -8.472908e-12, 
    -8.511127e-12, -8.470643e-12, -8.476093e-12, -8.473648e-12, 
    -8.443923e-12, -8.428942e-12, -8.397575e-12, -8.40327e-12, -8.426309e-12, 
    -8.478544e-12, -8.460814e-12, -8.505503e-12, -8.504494e-12, 
    -8.554248e-12, -8.531815e-12, -8.615448e-12, -8.591678e-12, 
    -8.660371e-12, -8.643095e-12, -8.659559e-12, -8.654567e-12, 
    -8.659624e-12, -8.634287e-12, -8.645142e-12, -8.622847e-12, 
    -8.536016e-12, -8.561533e-12, -8.485429e-12, -8.43967e-12, -8.409283e-12, 
    -8.387718e-12, -8.390767e-12, -8.396579e-12, -8.426444e-12, 
    -8.454526e-12, -8.475927e-12, -8.490243e-12, -8.504349e-12, 
    -8.547043e-12, -8.569646e-12, -8.620254e-12, -8.611122e-12, 
    -8.626593e-12, -8.641376e-12, -8.666194e-12, -8.662109e-12, 
    -8.673042e-12, -8.626187e-12, -8.657326e-12, -8.60592e-12, -8.61998e-12, 
    -8.508178e-12, -8.465597e-12, -8.447494e-12, -8.431653e-12, 
    -8.393111e-12, -8.419727e-12, -8.409234e-12, -8.434198e-12, -8.45006e-12, 
    -8.442215e-12, -8.490634e-12, -8.471809e-12, -8.570985e-12, 
    -8.528266e-12, -8.639651e-12, -8.612997e-12, -8.646041e-12, 
    -8.629179e-12, -8.658071e-12, -8.632069e-12, -8.677112e-12, -8.68692e-12, 
    -8.680218e-12, -8.705967e-12, -8.630627e-12, -8.659558e-12, 
    -8.441994e-12, -8.443274e-12, -8.449235e-12, -8.423032e-12, 
    -8.421429e-12, -8.397419e-12, -8.418784e-12, -8.427882e-12, 
    -8.450979e-12, -8.464641e-12, -8.477629e-12, -8.506185e-12, 
    -8.538078e-12, -8.582679e-12, -8.614724e-12, -8.636205e-12, 
    -8.623034e-12, -8.634662e-12, -8.621662e-12, -8.61557e-12, -8.683245e-12, 
    -8.645243e-12, -8.702263e-12, -8.699108e-12, -8.673303e-12, 
    -8.699464e-12, -8.444172e-12, -8.43681e-12, -8.411247e-12, -8.431252e-12, 
    -8.394804e-12, -8.415205e-12, -8.426935e-12, -8.472201e-12, 
    -8.482149e-12, -8.491371e-12, -8.509586e-12, -8.532963e-12, 
    -8.573973e-12, -8.609657e-12, -8.642236e-12, -8.639849e-12, -8.64069e-12, 
    -8.647967e-12, -8.62994e-12, -8.650926e-12, -8.654449e-12, -8.64524e-12, 
    -8.698686e-12, -8.683416e-12, -8.699041e-12, -8.689099e-12, 
    -8.439203e-12, -8.451593e-12, -8.444898e-12, -8.457486e-12, 
    -8.448617e-12, -8.488053e-12, -8.499878e-12, -8.55521e-12, -8.532503e-12, 
    -8.568644e-12, -8.536174e-12, -8.541927e-12, -8.56982e-12, -8.537929e-12, 
    -8.607689e-12, -8.560391e-12, -8.64825e-12, -8.601013e-12, -8.65121e-12, 
    -8.642096e-12, -8.657187e-12, -8.670702e-12, -8.687708e-12, 
    -8.719083e-12, -8.711818e-12, -8.738059e-12, -8.470062e-12, 
    -8.486131e-12, -8.484718e-12, -8.501535e-12, -8.513973e-12, 
    -8.540933e-12, -8.584173e-12, -8.567913e-12, -8.597766e-12, 
    -8.603758e-12, -8.558406e-12, -8.586251e-12, -8.496887e-12, 
    -8.511323e-12, -8.502728e-12, -8.47133e-12, -8.571658e-12, -8.520167e-12, 
    -8.615253e-12, -8.587357e-12, -8.668775e-12, -8.628282e-12, 
    -8.707818e-12, -8.741818e-12, -8.773825e-12, -8.811223e-12, 
    -8.494903e-12, -8.483984e-12, -8.503536e-12, -8.530585e-12, 
    -8.555687e-12, -8.589058e-12, -8.592474e-12, -8.598725e-12, -8.61492e-12, 
    -8.628536e-12, -8.600701e-12, -8.63195e-12, -8.514669e-12, -8.576129e-12, 
    -8.479855e-12, -8.508842e-12, -8.528991e-12, -8.520153e-12, 
    -8.566055e-12, -8.576874e-12, -8.620837e-12, -8.598111e-12, 
    -8.733425e-12, -8.673556e-12, -8.839705e-12, -8.793269e-12, 
    -8.480169e-12, -8.494865e-12, -8.546017e-12, -8.521679e-12, 
    -8.591287e-12, -8.608421e-12, -8.622351e-12, -8.640157e-12, -8.64208e-12, 
    -8.652631e-12, -8.635342e-12, -8.651948e-12, -8.589129e-12, 
    -8.617202e-12, -8.540171e-12, -8.558918e-12, -8.550294e-12, 
    -8.540834e-12, -8.570033e-12, -8.601139e-12, -8.601805e-12, -8.61178e-12, 
    -8.639884e-12, -8.591569e-12, -8.741149e-12, -8.648766e-12, 
    -8.510893e-12, -8.5392e-12, -8.543246e-12, -8.532279e-12, -8.606703e-12, 
    -8.579736e-12, -8.652373e-12, -8.632742e-12, -8.664908e-12, 
    -8.648924e-12, -8.646572e-12, -8.626043e-12, -8.613262e-12, 
    -8.580972e-12, -8.5547e-12, -8.53387e-12, -8.538714e-12, -8.561596e-12, 
    -8.603042e-12, -8.642254e-12, -8.633664e-12, -8.662464e-12, 
    -8.586239e-12, -8.6182e-12, -8.605847e-12, -8.638058e-12, -8.567481e-12, 
    -8.627575e-12, -8.55212e-12, -8.558735e-12, -8.579201e-12, -8.620367e-12, 
    -8.629477e-12, -8.639201e-12, -8.633202e-12, -8.604095e-12, 
    -8.599327e-12, -8.578704e-12, -8.573009e-12, -8.557295e-12, 
    -8.544286e-12, -8.556171e-12, -8.568654e-12, -8.604107e-12, 
    -8.636058e-12, -8.670894e-12, -8.679421e-12, -8.720121e-12, 
    -8.686987e-12, -8.741664e-12, -8.695174e-12, -8.775655e-12, 
    -8.631061e-12, -8.69381e-12, -8.580132e-12, -8.592379e-12, -8.614527e-12, 
    -8.665334e-12, -8.637907e-12, -8.669984e-12, -8.59914e-12, -8.562385e-12, 
    -8.552877e-12, -8.535136e-12, -8.553283e-12, -8.551808e-12, 
    -8.569172e-12, -8.563592e-12, -8.605285e-12, -8.582889e-12, 
    -8.646512e-12, -8.669732e-12, -8.735308e-12, -8.77551e-12, -8.816438e-12, 
    -8.834507e-12, -8.840007e-12, -8.842306e-12 ;

 SMIN_NH4 =
  0.0004353462, 0.00043718, 0.0004368234, 0.0004383026, 0.000437482, 
    0.0004384504, 0.0004357177, 0.0004372525, 0.0004362726, 0.0004355108, 
    0.0004411724, 0.0004383681, 0.0004440855, 0.0004422969, 0.0004467897, 
    0.000443807, 0.0004473911, 0.0004467036, 0.0004487727, 0.0004481798, 
    0.000450826, 0.0004490461, 0.0004521978, 0.0004504009, 0.0004506819, 
    0.0004489871, 0.0004389329, 0.0004408236, 0.0004388208, 0.0004390904, 
    0.0004389693, 0.0004374987, 0.0004367575, 0.0004352055, 0.0004354872, 
    0.0004366271, 0.0004392112, 0.000438334, 0.0004405447, 0.0004404948, 
    0.0004429559, 0.0004418462, 0.0004459828, 0.0004448071, 0.0004482045, 
    0.00044735, 0.0004481643, 0.0004479173, 0.0004481673, 0.0004469142, 
    0.000447451, 0.0004463484, 0.0004420547, 0.0004433168, 0.0004395522, 
    0.0004372883, 0.0004357848, 0.0004347179, 0.0004348686, 0.0004351561, 
    0.0004366337, 0.0004380229, 0.0004390816, 0.0004397898, 0.0004404875, 
    0.0004425995, 0.0004437174, 0.0004462204, 0.0004457688, 0.0004465339, 
    0.000447265, 0.0004484922, 0.0004482902, 0.0004488309, 0.0004465134, 
    0.0004480535, 0.000445511, 0.0004462064, 0.0004406775, 0.0004385709, 
    0.0004376753, 0.0004368915, 0.0004349845, 0.0004363014, 0.0004357822, 
    0.0004370172, 0.0004378019, 0.0004374137, 0.0004398091, 0.0004388777, 
    0.0004437836, 0.0004416704, 0.0004471797, 0.0004458613, 0.0004474956, 
    0.0004466617, 0.0004480904, 0.0004468044, 0.000449032, 0.000449517, 
    0.0004491855, 0.0004504588, 0.0004467328, 0.0004481637, 0.0004374031, 
    0.0004374664, 0.0004377613, 0.0004364648, 0.0004363855, 0.0004351975, 
    0.0004362545, 0.0004367046, 0.0004378473, 0.000438523, 0.0004391655, 
    0.0004405782, 0.0004421557, 0.0004443618, 0.0004459467, 0.000447009, 
    0.0004463576, 0.0004469326, 0.0004462897, 0.0004459883, 0.0004493351, 
    0.0004474558, 0.0004502755, 0.0004501195, 0.0004488433, 0.000450137, 
    0.0004375108, 0.0004371464, 0.0004358817, 0.0004368714, 0.000435068, 
    0.0004360774, 0.0004366577, 0.000438897, 0.0004393891, 0.0004398453, 
    0.0004407463, 0.0004419026, 0.0004439311, 0.000445696, 0.0004473073, 
    0.0004471891, 0.0004472307, 0.0004475905, 0.0004466989, 0.0004477368, 
    0.0004479109, 0.0004474554, 0.0004500985, 0.0004493434, 0.000450116, 
    0.0004496243, 0.0004372648, 0.0004378776, 0.0004375463, 0.0004381691, 
    0.0004377303, 0.0004396812, 0.0004402661, 0.0004430031, 0.0004418798, 
    0.0004436676, 0.0004420613, 0.0004423459, 0.0004437256, 0.000442148, 
    0.0004455985, 0.000443259, 0.0004476044, 0.0004452681, 0.0004477507, 
    0.0004472999, 0.0004480461, 0.0004487146, 0.0004495554, 0.000451107, 
    0.0004507476, 0.0004520452, 0.0004387913, 0.0004395862, 0.0004395162, 
    0.0004403481, 0.0004409633, 0.0004422969, 0.0004444357, 0.0004436313, 
    0.0004451078, 0.0004454042, 0.0004431609, 0.0004445381, 0.0004401177, 
    0.0004408317, 0.0004404065, 0.0004388531, 0.0004438161, 0.000441269, 
    0.0004459723, 0.0004445924, 0.0004486191, 0.0004466165, 0.0004505498, 
    0.0004522311, 0.0004538137, 0.0004556628, 0.00044002, 0.0004394798, 
    0.0004404469, 0.000441785, 0.0004430266, 0.0004446772, 0.0004448461, 
    0.0004451552, 0.0004459561, 0.0004466296, 0.0004452528, 0.0004467983, 
    0.0004409972, 0.0004440372, 0.0004392748, 0.0004407088, 0.0004417054, 
    0.0004412682, 0.0004435387, 0.0004440737, 0.0004462481, 0.0004451241, 
    0.000451816, 0.0004488553, 0.0004570708, 0.0004547749, 0.000439291, 
    0.000440018, 0.0004425482, 0.0004413443, 0.0004447873, 0.0004456348, 
    0.0004463236, 0.0004472042, 0.0004472992, 0.000447821, 0.0004469659, 
    0.0004477872, 0.0004446801, 0.0004460686, 0.0004422584, 0.0004431857, 
    0.0004427591, 0.000442291, 0.0004437352, 0.0004452738, 0.0004453067, 
    0.0004458, 0.00044719, 0.0004448002, 0.0004521977, 0.000447629, 
    0.0004408107, 0.0004422109, 0.000442411, 0.0004418685, 0.0004455496, 
    0.0004442158, 0.0004478083, 0.0004468373, 0.0004484281, 0.0004476376, 
    0.0004475212, 0.0004465058, 0.0004458736, 0.0004442765, 0.0004429769, 
    0.0004419466, 0.000442186, 0.0004433179, 0.0004453678, 0.0004473072, 
    0.0004468822, 0.0004483065, 0.0004445365, 0.0004461173, 0.0004455062, 
    0.0004470994, 0.0004436097, 0.0004465821, 0.0004428498, 0.000443177, 
    0.0004441892, 0.0004462253, 0.0004466758, 0.0004471567, 0.0004468598, 
    0.0004454202, 0.0004451844, 0.0004441642, 0.0004438825, 0.0004431053, 
    0.0004424616, 0.0004430496, 0.0004436669, 0.0004454204, 0.0004470006, 
    0.0004487234, 0.000449145, 0.0004511577, 0.0004495191, 0.0004522229, 
    0.0004499239, 0.0004539035, 0.0004467543, 0.0004498576, 0.0004442353, 
    0.0004448409, 0.0004459364, 0.000448449, 0.0004470925, 0.0004486789, 
    0.0004451751, 0.000443357, 0.0004428867, 0.0004420091, 0.0004429066, 
    0.0004428336, 0.0004436925, 0.0004434164, 0.0004454785, 0.0004443708, 
    0.0004475175, 0.0004486658, 0.0004519086, 0.0004538964, 0.00045592, 
    0.0004568133, 0.0004570851, 0.0004571987 ;

 SMIN_NH4_vr =
  0.002856641, 0.002861575, 0.002860609, 0.002864585, 0.002862377, 
    0.002864974, 0.002857627, 0.002861748, 0.002859114, 0.00285706, 
    0.00287226, 0.002864738, 0.002880068, 0.002875273, 0.002887296, 
    0.002879313, 0.0028889, 0.002887059, 0.002892588, 0.002891, 0.002898056, 
    0.00289331, 0.002901709, 0.002896918, 0.002897663, 0.002893138, 
    0.002866277, 0.002871347, 0.002865969, 0.002866693, 0.002866365, 
    0.002862409, 0.002860413, 0.002856236, 0.00285699, 0.002860056, 
    0.002866996, 0.002864637, 0.002870569, 0.002870436, 0.002877027, 
    0.002874054, 0.002885129, 0.002881978, 0.002891062, 0.002888774, 
    0.002890948, 0.002890284, 0.002890948, 0.002887599, 0.002889028, 
    0.002886081, 0.002874648, 0.002878025, 0.002867928, 0.002861838, 
    0.002857794, 0.002854924, 0.002855323, 0.002856097, 0.002860068, 
    0.002863799, 0.002866642, 0.002868538, 0.002870407, 0.002876067, 
    0.002879061, 0.002885756, 0.002884548, 0.002886589, 0.002888543, 
    0.002891818, 0.002891277, 0.002892716, 0.00288652, 0.002890636, 
    0.002883833, 0.002885693, 0.00287094, 0.002865287, 0.002862876, 
    0.002860766, 0.002855633, 0.002859176, 0.002857776, 0.002861093, 
    0.002863201, 0.002862154, 0.002868587, 0.002866081, 0.002879233, 
    0.002873572, 0.002888319, 0.002884789, 0.002889155, 0.002886927, 
    0.002890738, 0.002887303, 0.002893247, 0.002894542, 0.002893651, 
    0.00289705, 0.002887093, 0.002890917, 0.002862143, 0.002862313, 
    0.002863102, 0.002859611, 0.002859396, 0.002856196, 0.002859036, 
    0.002860247, 0.002863316, 0.002865126, 0.002866848, 0.00287064, 
    0.002874867, 0.002880773, 0.002885014, 0.002887851, 0.002886108, 
    0.002887641, 0.00288592, 0.00288511, 0.002894048, 0.002889029, 
    0.002896553, 0.002896137, 0.002892726, 0.002896175, 0.002862427, 
    0.002861443, 0.002858039, 0.002860697, 0.002855842, 0.002858558, 
    0.002860114, 0.002866128, 0.002867447, 0.002868671, 0.002871086, 
    0.002874183, 0.002879616, 0.002884336, 0.002888645, 0.002888324, 
    0.002888434, 0.002889391, 0.002887006, 0.002889776, 0.002890236, 
    0.002889021, 0.002896072, 0.002894058, 0.002896116, 0.002894799, 
    0.002861758, 0.0028634, 0.002862506, 0.00286418, 0.002862994, 
    0.002868233, 0.002869799, 0.002877134, 0.002874121, 0.002878912, 
    0.002874602, 0.002875365, 0.002879055, 0.002874827, 0.002884065, 
    0.002877795, 0.002889425, 0.002883168, 0.00288981, 0.002888601, 
    0.002890591, 0.002892376, 0.002894615, 0.002898754, 0.00289779, 
    0.00290125, 0.002865851, 0.00286798, 0.002867793, 0.00287002, 
    0.002871667, 0.002875244, 0.00288097, 0.002878811, 0.002882761, 
    0.002883554, 0.002877542, 0.00288123, 0.002869376, 0.002871287, 
    0.002870146, 0.002865971, 0.00287928, 0.002872448, 0.002885047, 
    0.00288135, 0.002892113, 0.002886761, 0.00289726, 0.002901741, 
    0.002905955, 0.002910867, 0.002869142, 0.002867688, 0.00287028, 
    0.002873868, 0.002877191, 0.002881612, 0.002882061, 0.002882883, 
    0.002885023, 0.002886825, 0.002883136, 0.002887267, 0.002871724, 
    0.002879872, 0.002867098, 0.002870945, 0.002873613, 0.002872442, 
    0.002878525, 0.002879953, 0.002885767, 0.002882762, 0.002900625, 
    0.002892728, 0.002914606, 0.002908501, 0.002867178, 0.002869125, 
    0.002875906, 0.00287268, 0.002881899, 0.002884167, 0.002886004, 
    0.002888358, 0.002888606, 0.002890001, 0.002887709, 0.002889905, 
    0.002881588, 0.002885304, 0.002875098, 0.002877578, 0.002876434, 
    0.002875175, 0.002879041, 0.002883159, 0.002883245, 0.002884559, 
    0.002888268, 0.002881879, 0.002901627, 0.002889432, 0.002871249, 
    0.002874997, 0.002875531, 0.002874078, 0.002883931, 0.002880361, 
    0.002889967, 0.002887368, 0.002891615, 0.002889503, 0.002889185, 
    0.002886472, 0.002884774, 0.0028805, 0.002877012, 0.002874252, 
    0.002874888, 0.002877921, 0.002883402, 0.00288859, 0.00288745, 
    0.002891253, 0.002881167, 0.002885396, 0.002883755, 0.002888017, 
    0.002878741, 0.002886691, 0.002876703, 0.002877575, 0.002880281, 
    0.002885729, 0.002886929, 0.002888215, 0.002887416, 0.002883565, 
    0.00288293, 0.002880195, 0.002879436, 0.002877356, 0.002875624, 
    0.0028772, 0.002878847, 0.002883543, 0.002887764, 0.002892363, 
    0.002893489, 0.002898849, 0.002894477, 0.002901679, 0.002895547, 
    0.002906152, 0.002887145, 0.002895435, 0.002880406, 0.002882023, 
    0.00288495, 0.002891662, 0.002888035, 0.002892273, 0.002882903, 
    0.002878029, 0.002876767, 0.002874415, 0.002876815, 0.00287662, 
    0.002878917, 0.002878173, 0.002883689, 0.002880726, 0.002889135, 
    0.002892203, 0.002900851, 0.00290614, 0.002911525, 0.002913895, 
    0.002914616, 0.002914914,
  0.001594047, 0.001600114, 0.001598935, 0.001603825, 0.001601113, 
    0.001604314, 0.001595278, 0.001600354, 0.001597114, 0.001594594, 
    0.001613302, 0.001604043, 0.001622913, 0.001617017, 0.00163182, 
    0.001621995, 0.0016338, 0.001631538, 0.001638346, 0.001636396, 
    0.001645092, 0.001639245, 0.001649598, 0.001643697, 0.00164462, 
    0.001639052, 0.001605909, 0.00161215, 0.001605538, 0.001606429, 
    0.00160603, 0.001601169, 0.001598717, 0.001593584, 0.001594516, 
    0.001598287, 0.001606829, 0.001603932, 0.001611235, 0.00161107, 
    0.001619191, 0.00161553, 0.001629166, 0.001625293, 0.001636478, 
    0.001633667, 0.001636345, 0.001635533, 0.001636356, 0.001632233, 
    0.001634, 0.001630371, 0.001616216, 0.001620379, 0.001607955, 
    0.001600472, 0.0015955, 0.001591969, 0.001592468, 0.00159342, 
    0.001598309, 0.001602904, 0.001606403, 0.001608742, 0.001611046, 
    0.001618013, 0.001621701, 0.001629948, 0.001628461, 0.00163098, 
    0.001633387, 0.001637424, 0.00163676, 0.001638538, 0.001630914, 
    0.001635982, 0.001627614, 0.001629904, 0.001611668, 0.001604714, 
    0.001601752, 0.001599161, 0.001592852, 0.00159721, 0.001595492, 
    0.001599578, 0.001602173, 0.00160089, 0.001608806, 0.001605729, 
    0.001621919, 0.00161495, 0.001633106, 0.001628766, 0.001634146, 
    0.001631402, 0.001636103, 0.001631872, 0.0016392, 0.001640794, 
    0.001639705, 0.00164389, 0.001631637, 0.001636345, 0.001600854, 
    0.001601063, 0.001602038, 0.00159775, 0.001597488, 0.001593558, 
    0.001597056, 0.001598544, 0.001602324, 0.001604557, 0.00160668, 
    0.001611346, 0.001616552, 0.001623826, 0.001629048, 0.001632545, 
    0.001630401, 0.001632294, 0.001630178, 0.001629186, 0.001640196, 
    0.001634016, 0.001643288, 0.001642775, 0.00163858, 0.001642833, 
    0.00160121, 0.001600006, 0.001595822, 0.001599096, 0.00159313, 
    0.00159647, 0.001598389, 0.001605793, 0.001607419, 0.001608926, 
    0.001611902, 0.001615718, 0.001622407, 0.001628222, 0.001633527, 
    0.001633139, 0.001633275, 0.001634459, 0.001631525, 0.001634941, 
    0.001635514, 0.001634016, 0.001642707, 0.001640225, 0.001642764, 
    0.001641149, 0.001600398, 0.001602424, 0.001601329, 0.001603387, 
    0.001601937, 0.001608383, 0.001610314, 0.001619347, 0.001615642, 
    0.001621538, 0.001616242, 0.00161718, 0.001621728, 0.001616528, 
    0.001627901, 0.001620191, 0.001634505, 0.001626812, 0.001634987, 
    0.001633504, 0.00163596, 0.001638158, 0.001640922, 0.001646019, 
    0.00164484, 0.001649101, 0.001605444, 0.001608069, 0.001607839, 
    0.001610587, 0.001612618, 0.001617019, 0.00162407, 0.00162142, 
    0.001626286, 0.001627262, 0.001619869, 0.001624408, 0.001609827, 
    0.001612184, 0.001610781, 0.00160565, 0.001622029, 0.001613628, 
    0.001629134, 0.001624589, 0.001637844, 0.001631255, 0.00164419, 
    0.001649709, 0.001654903, 0.001660963, 0.001609503, 0.001607719, 
    0.001610914, 0.001615329, 0.001619425, 0.001624866, 0.001625423, 
    0.001626442, 0.00162908, 0.001631297, 0.001626763, 0.001631853, 
    0.001612729, 0.001622758, 0.001607044, 0.001611779, 0.001615069, 
    0.001613627, 0.001621117, 0.001622881, 0.001630043, 0.001626342, 
    0.001648347, 0.00163862, 0.001665575, 0.001658054, 0.001607096, 
    0.001609497, 0.001617847, 0.001613876, 0.00162523, 0.001628021, 
    0.00163029, 0.001633188, 0.001633502, 0.001635218, 0.001632405, 
    0.001635107, 0.001624878, 0.001629451, 0.001616895, 0.001619952, 
    0.001618546, 0.001617003, 0.001621765, 0.001626834, 0.001626944, 
    0.001628568, 0.00163314, 0.001625276, 0.001649598, 0.001634586, 
    0.001612115, 0.001616734, 0.001617396, 0.001615607, 0.001627741, 
    0.001623347, 0.001635176, 0.001631982, 0.001637216, 0.001634615, 
    0.001634232, 0.001630891, 0.00162881, 0.001623548, 0.001619264, 
    0.001615866, 0.001616657, 0.001620389, 0.001627144, 0.001633529, 
    0.001632131, 0.001636818, 0.001624407, 0.001629613, 0.001627601, 
    0.001632847, 0.001621349, 0.001631137, 0.001618844, 0.001619923, 
    0.00162326, 0.001629965, 0.00163145, 0.001633033, 0.001632057, 
    0.001627316, 0.00162654, 0.001623179, 0.00162225, 0.001619688, 
    0.001617566, 0.001619505, 0.00162154, 0.001627318, 0.001632521, 
    0.001638189, 0.001639575, 0.001646186, 0.001640803, 0.001649681, 
    0.001642131, 0.001655197, 0.001631706, 0.001641912, 0.001623412, 
    0.001625408, 0.001629015, 0.001637283, 0.001632822, 0.00163804, 
    0.001626509, 0.001620517, 0.001618968, 0.001616073, 0.001619034, 
    0.001618793, 0.001621625, 0.001620715, 0.00162751, 0.001623861, 
    0.001634222, 0.001637999, 0.001648654, 0.001655175, 0.001661809, 
    0.001664735, 0.001665625, 0.001665997,
  0.001500661, 0.001507298, 0.001506009, 0.00151136, 0.001508392, 
    0.001511895, 0.001502007, 0.001507562, 0.001504016, 0.001501259, 
    0.001521736, 0.001511598, 0.001532258, 0.0015258, 0.001542016, 
    0.001531253, 0.001544185, 0.001541706, 0.001549166, 0.001547029, 
    0.001556563, 0.001550152, 0.001561502, 0.001555033, 0.001556045, 
    0.00154994, 0.00151364, 0.001520474, 0.001513235, 0.00151421, 
    0.001513772, 0.001508453, 0.001505771, 0.001500154, 0.001501174, 
    0.0015053, 0.001514648, 0.001511476, 0.00151947, 0.001519289, 
    0.001528181, 0.001524173, 0.001539107, 0.001534865, 0.001547119, 
    0.001544038, 0.001546974, 0.001546084, 0.001546985, 0.001542467, 
    0.001544403, 0.001540427, 0.001524923, 0.001529482, 0.00151588, 
    0.001507691, 0.001502251, 0.001498388, 0.001498934, 0.001499975, 
    0.001505324, 0.001510351, 0.00151418, 0.001516741, 0.001519263, 
    0.001526893, 0.001530931, 0.001539964, 0.001538335, 0.001541095, 
    0.001543732, 0.001548156, 0.001547428, 0.001549377, 0.001541023, 
    0.001546576, 0.001537407, 0.001539915, 0.001519946, 0.001512332, 
    0.001509092, 0.001506256, 0.001499354, 0.001504121, 0.001502242, 
    0.001506712, 0.001509552, 0.001508147, 0.001516811, 0.001513444, 
    0.00153117, 0.001523538, 0.001543424, 0.001538669, 0.001544564, 
    0.001541557, 0.001546708, 0.001542072, 0.001550102, 0.00155185, 
    0.001550656, 0.001555243, 0.001541815, 0.001546974, 0.001508108, 
    0.001508337, 0.001509404, 0.001504713, 0.001504426, 0.001500126, 
    0.001503952, 0.001505581, 0.001509716, 0.001512161, 0.001514485, 
    0.001519592, 0.001525292, 0.001533258, 0.001538978, 0.00154281, 
    0.00154046, 0.001542534, 0.001540216, 0.001539129, 0.001551195, 
    0.001544421, 0.001554583, 0.001554021, 0.001549423, 0.001554085, 
    0.001508498, 0.00150718, 0.001502602, 0.001506185, 0.001499657, 
    0.001503311, 0.001505412, 0.001513513, 0.001515293, 0.001516943, 
    0.0015202, 0.001524378, 0.001531704, 0.001538074, 0.001543885, 
    0.00154346, 0.001543609, 0.001544907, 0.001541692, 0.001545435, 
    0.001546063, 0.001544421, 0.001553946, 0.001551226, 0.00155401, 
    0.001552238, 0.001507608, 0.001509826, 0.001508628, 0.001510881, 
    0.001509293, 0.001516349, 0.001518463, 0.001528352, 0.001524296, 
    0.001530752, 0.001524952, 0.00152598, 0.001530961, 0.001525266, 
    0.001537722, 0.001529278, 0.001544958, 0.00153653, 0.001545485, 
    0.00154386, 0.001546551, 0.00154896, 0.00155199, 0.001557578, 
    0.001556285, 0.001560957, 0.001513131, 0.001516005, 0.001515753, 
    0.00151876, 0.001520984, 0.001525802, 0.001533525, 0.001530622, 
    0.001535952, 0.001537021, 0.001528924, 0.001533896, 0.001517929, 
    0.00152051, 0.001518973, 0.001513358, 0.00153129, 0.001522091, 
    0.001539072, 0.001534093, 0.001548616, 0.001541396, 0.001555573, 
    0.001561625, 0.00156732, 0.001573969, 0.001517574, 0.001515621, 
    0.001519118, 0.001523953, 0.001528438, 0.001534397, 0.001535007, 
    0.001536123, 0.001539013, 0.001541442, 0.001536475, 0.001542051, 
    0.001521107, 0.001532088, 0.001514883, 0.001520066, 0.001523668, 
    0.001522089, 0.00153029, 0.001532222, 0.001540068, 0.001536013, 
    0.001560131, 0.001549468, 0.001579029, 0.001570778, 0.001514939, 
    0.001517568, 0.00152671, 0.001522361, 0.001534795, 0.001537853, 
    0.001540339, 0.001543514, 0.001543857, 0.001545739, 0.001542656, 
    0.001545617, 0.00153441, 0.00153942, 0.001525666, 0.001529015, 
    0.001527475, 0.001525785, 0.001531, 0.001536553, 0.001536672, 
    0.001538452, 0.001543464, 0.001534845, 0.001561505, 0.001545048, 
    0.001520433, 0.001525492, 0.001526215, 0.001524256, 0.001537546, 
    0.001532733, 0.001545693, 0.001542192, 0.001547928, 0.001545078, 
    0.001544658, 0.001540997, 0.001538717, 0.001532953, 0.001528262, 
    0.00152454, 0.001525406, 0.001529493, 0.001536893, 0.001543888, 
    0.001542356, 0.001547492, 0.001533894, 0.001539598, 0.001537393, 
    0.00154314, 0.001530544, 0.001541269, 0.001527801, 0.001528983, 
    0.001532637, 0.001539984, 0.00154161, 0.001543344, 0.001542274, 
    0.001537081, 0.00153623, 0.001532549, 0.001531531, 0.001528725, 
    0.001526401, 0.001528525, 0.001530754, 0.001537083, 0.001542783, 
    0.001548994, 0.001550514, 0.001557763, 0.001551861, 0.001561597, 
    0.001553319, 0.001567645, 0.001541891, 0.001553077, 0.001532804, 
    0.00153499, 0.001538942, 0.001548003, 0.001543113, 0.001548832, 
    0.001536197, 0.001529634, 0.001527936, 0.001524766, 0.001528009, 
    0.001527745, 0.001530847, 0.00152985, 0.001537293, 0.001533296, 
    0.001544648, 0.001548787, 0.001560467, 0.00156762, 0.001574896, 
    0.001578106, 0.001579083, 0.001579492,
  0.00142892, 0.001435685, 0.00143437, 0.001439825, 0.001436799, 0.001440371, 
    0.001430292, 0.001435953, 0.001432339, 0.001429529, 0.00145041, 
    0.001440069, 0.001461149, 0.001454556, 0.001471115, 0.001460123, 
    0.001473331, 0.001470799, 0.001478422, 0.001476238, 0.001485987, 
    0.00147943, 0.001491039, 0.001484421, 0.001485456, 0.001479213, 
    0.00144215, 0.001449122, 0.001441737, 0.001442731, 0.001442285, 
    0.001436862, 0.001434128, 0.001428403, 0.001429443, 0.001433647, 
    0.001443178, 0.001439943, 0.001448096, 0.001447912, 0.001456986, 
    0.001452895, 0.001468143, 0.00146381, 0.001476329, 0.001473181, 
    0.001476181, 0.001475272, 0.001476193, 0.001471576, 0.001473554, 
    0.001469491, 0.001453661, 0.001458314, 0.001444434, 0.001436086, 
    0.00143054, 0.001426604, 0.00142716, 0.001428221, 0.001433672, 
    0.001438796, 0.001442701, 0.001445312, 0.001447885, 0.001455672, 
    0.001459793, 0.001469019, 0.001467354, 0.001470174, 0.001472868, 
    0.00147739, 0.001476646, 0.001478638, 0.0014701, 0.001475775, 
    0.001466406, 0.001468969, 0.001448584, 0.001440816, 0.001437513, 
    0.001434623, 0.001427588, 0.001432446, 0.001430531, 0.001435087, 
    0.001437981, 0.00143655, 0.001445384, 0.00144195, 0.001460038, 
    0.001452248, 0.001472554, 0.001467696, 0.001473718, 0.001470645, 
    0.00147591, 0.001471172, 0.00147938, 0.001481166, 0.001479945, 
    0.001484636, 0.001470909, 0.001476181, 0.00143651, 0.001436743, 
    0.001437831, 0.001433049, 0.001432757, 0.001428375, 0.001432274, 
    0.001433934, 0.001438149, 0.001440642, 0.001443011, 0.00144822, 
    0.001454037, 0.001462169, 0.001468011, 0.001471926, 0.001469525, 
    0.001471645, 0.001469275, 0.001468165, 0.001480497, 0.001473573, 
    0.001483961, 0.001483387, 0.001478686, 0.001483451, 0.001436907, 
    0.001435564, 0.001430898, 0.001434549, 0.001427897, 0.001431621, 
    0.001433762, 0.001442021, 0.001443836, 0.001445518, 0.001448841, 
    0.001453104, 0.001460582, 0.001467087, 0.001473025, 0.00147259, 
    0.001472743, 0.001474069, 0.001470784, 0.001474608, 0.00147525, 
    0.001473572, 0.00148331, 0.001480528, 0.001483374, 0.001481563, 0.001436, 
    0.001438261, 0.001437039, 0.001439336, 0.001437718, 0.001444913, 
    0.00144707, 0.001457161, 0.00145302, 0.001459611, 0.00145369, 
    0.001454739, 0.001459825, 0.00145401, 0.001466729, 0.001458106, 
    0.001474121, 0.001465512, 0.00147466, 0.001472999, 0.001475749, 
    0.001478212, 0.00148131, 0.001487025, 0.001485702, 0.001490481, 
    0.001441631, 0.001444562, 0.001444304, 0.001447372, 0.001449641, 
    0.001454558, 0.001462442, 0.001459477, 0.00146492, 0.001466012, 
    0.001457744, 0.001462821, 0.001446524, 0.001449158, 0.00144759, 
    0.001441862, 0.00146016, 0.001450771, 0.001468107, 0.001463022, 
    0.001477861, 0.001470482, 0.001484973, 0.001491166, 0.001496993, 
    0.001503802, 0.001446162, 0.001444171, 0.001447737, 0.001452671, 
    0.001457248, 0.001463332, 0.001463955, 0.001465095, 0.001468046, 
    0.001470528, 0.001465455, 0.00147115, 0.001449768, 0.001460975, 
    0.001443417, 0.001448705, 0.00145238, 0.001450768, 0.001459138, 
    0.001461111, 0.001469125, 0.001464983, 0.001489638, 0.001478732, 
    0.001508985, 0.001500533, 0.001443475, 0.001446156, 0.001455485, 
    0.001451046, 0.001463739, 0.001466862, 0.001469401, 0.001472646, 
    0.001472996, 0.001474919, 0.001471768, 0.001474794, 0.001463345, 
    0.001468462, 0.001454419, 0.001457837, 0.001456265, 0.00145454, 
    0.001459864, 0.001465535, 0.001465656, 0.001467474, 0.001472597, 
    0.00146379, 0.001491045, 0.001474215, 0.001449079, 0.001454242, 
    0.001454979, 0.00145298, 0.001466549, 0.001461633, 0.001474872, 
    0.001471295, 0.001477156, 0.001474243, 0.001473815, 0.001470074, 
    0.001467744, 0.001461858, 0.001457068, 0.00145327, 0.001454153, 
    0.001458326, 0.001465882, 0.001473028, 0.001471463, 0.001476711, 
    0.001462818, 0.001468644, 0.001466393, 0.001472263, 0.001459399, 
    0.001470354, 0.001456598, 0.001457804, 0.001461535, 0.001469039, 
    0.0014707, 0.001472472, 0.001471378, 0.001466073, 0.001465204, 
    0.001461445, 0.001460406, 0.001457541, 0.001455169, 0.001457336, 
    0.001459613, 0.001466076, 0.001471899, 0.001478247, 0.0014798, 
    0.001487215, 0.001481179, 0.001491138, 0.001482671, 0.001497327, 
    0.001470989, 0.001482422, 0.001461705, 0.001463938, 0.001467975, 
    0.001477234, 0.001472236, 0.001478081, 0.00146517, 0.00145847, 
    0.001456736, 0.001453501, 0.00145681, 0.001456541, 0.001459707, 
    0.001458689, 0.00146629, 0.001462208, 0.001473804, 0.001478035, 
    0.00148998, 0.0014973, 0.00150475, 0.001508039, 0.00150904, 0.001509458,
  0.001343027, 0.001349267, 0.001348053, 0.001353088, 0.001350295, 
    0.001353592, 0.001344292, 0.001349515, 0.00134618, 0.001343588, 
    0.001362868, 0.001353313, 0.001372802, 0.001366701, 0.001382034, 
    0.001371852, 0.001384088, 0.00138174, 0.001388809, 0.001386783, 
    0.001395833, 0.001389744, 0.001400527, 0.001394378, 0.00139534, 
    0.001389544, 0.001355235, 0.001361678, 0.001354853, 0.001355772, 
    0.001355359, 0.001350353, 0.001347831, 0.00134255, 0.001343508, 
    0.001347387, 0.001356185, 0.001353197, 0.001360728, 0.001360558, 
    0.001368948, 0.001365164, 0.001379278, 0.001375265, 0.001386868, 
    0.001383948, 0.001386731, 0.001385887, 0.001386742, 0.001382461, 
    0.001384295, 0.001380528, 0.001365873, 0.001370178, 0.001357345, 
    0.001349637, 0.001344521, 0.001340892, 0.001341405, 0.001342383, 
    0.00134741, 0.001352138, 0.001355743, 0.001358156, 0.001360533, 
    0.001367734, 0.001371547, 0.00138009, 0.001378548, 0.001381161, 
    0.001383658, 0.001387852, 0.001387162, 0.00138901, 0.001381092, 
    0.001386354, 0.001377669, 0.001380044, 0.001361181, 0.001354003, 
    0.001350955, 0.001348287, 0.001341799, 0.001346279, 0.001344513, 
    0.001348715, 0.001351386, 0.001350065, 0.001358222, 0.00135505, 
    0.001371773, 0.001364566, 0.001383367, 0.001378864, 0.001384446, 
    0.001381597, 0.001386479, 0.001382086, 0.001389698, 0.001391357, 
    0.001390223, 0.001394577, 0.001381842, 0.001386731, 0.001350028, 
    0.001350243, 0.001351247, 0.001346835, 0.001346565, 0.001342524, 
    0.00134612, 0.001347651, 0.001351541, 0.001353842, 0.00135603, 
    0.001360843, 0.001366221, 0.001373746, 0.001379156, 0.001382784, 
    0.001380559, 0.001382524, 0.001380328, 0.001379299, 0.001390735, 
    0.001384312, 0.001393951, 0.001393417, 0.001389054, 0.001393477, 
    0.001350394, 0.001349155, 0.001344851, 0.001348219, 0.001342084, 
    0.001345517, 0.001347492, 0.001355116, 0.001356792, 0.001358346, 
    0.001361416, 0.001365358, 0.001372277, 0.001378301, 0.001383803, 
    0.0013834, 0.001383542, 0.001384772, 0.001381726, 0.001385272, 
    0.001385867, 0.001384311, 0.001393346, 0.001390764, 0.001393406, 
    0.001391725, 0.001349557, 0.001351644, 0.001350516, 0.001352637, 
    0.001351143, 0.001357787, 0.00135978, 0.001369111, 0.00136528, 
    0.001371378, 0.001365899, 0.00136687, 0.001371577, 0.001366195, 
    0.001377969, 0.001369986, 0.00138482, 0.001376842, 0.00138532, 
    0.00138378, 0.00138633, 0.001388614, 0.001391489, 0.001396797, 
    0.001395567, 0.001400007, 0.001354755, 0.001357463, 0.001357224, 
    0.001360059, 0.001362156, 0.001366702, 0.001373998, 0.001371254, 
    0.001376293, 0.001377304, 0.001369649, 0.001374349, 0.001359276, 
    0.00136171, 0.00136026, 0.001354969, 0.001371886, 0.001363201, 
    0.001379246, 0.001374535, 0.001388289, 0.001381447, 0.001394891, 
    0.001400645, 0.001406063, 0.001412399, 0.001358941, 0.001357101, 
    0.001360396, 0.001364957, 0.001369191, 0.001374823, 0.001375399, 
    0.001376455, 0.001379189, 0.001381489, 0.001376789, 0.001382066, 
    0.001362275, 0.001372641, 0.001356405, 0.001361291, 0.001364688, 
    0.001363198, 0.00137094, 0.001372766, 0.001380189, 0.001376351, 
    0.001399225, 0.001389097, 0.001417227, 0.001409357, 0.001356458, 
    0.001358935, 0.00136756, 0.001363455, 0.001375199, 0.001378092, 
    0.001380444, 0.001383452, 0.001383777, 0.00138556, 0.001382639, 
    0.001385444, 0.001374835, 0.001379574, 0.001366573, 0.001369736, 
    0.001368281, 0.001366685, 0.001371611, 0.001376863, 0.001376975, 
    0.001378659, 0.001383408, 0.001375246, 0.001400533, 0.001384909, 
    0.001361636, 0.001366411, 0.001367092, 0.001365242, 0.001377802, 
    0.001373249, 0.001385516, 0.001382199, 0.001387635, 0.001384933, 
    0.001384536, 0.001381068, 0.001378909, 0.001373458, 0.001369025, 
    0.001365511, 0.001366328, 0.001370188, 0.001377184, 0.001383807, 
    0.001382356, 0.001387222, 0.001374347, 0.001379743, 0.001377657, 
    0.001383098, 0.001371181, 0.001381329, 0.001368589, 0.001369705, 
    0.001373159, 0.00138011, 0.001381648, 0.001383291, 0.001382277, 
    0.001377361, 0.001376556, 0.001373075, 0.001372114, 0.001369462, 
    0.001367267, 0.001369273, 0.001371379, 0.001377363, 0.00138276, 
    0.001388647, 0.001390088, 0.001396974, 0.001391369, 0.00140062, 
    0.001392755, 0.001406374, 0.001381917, 0.001392523, 0.001373316, 
    0.001375383, 0.001379124, 0.001387708, 0.001383072, 0.001388494, 
    0.001376525, 0.001370321, 0.001368717, 0.001365724, 0.001368785, 
    0.001368536, 0.001371466, 0.001370525, 0.001377562, 0.001373781, 
    0.001384526, 0.001388451, 0.001399542, 0.001406349, 0.001413282, 
    0.001416345, 0.001417278, 0.001417667,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.21443e-06, 1.224907e-06, 1.222866e-06, 1.231344e-06, 1.226637e-06, 
    1.232193e-06, 1.21655e-06, 1.225323e-06, 1.219718e-06, 1.21537e-06, 
    1.24788e-06, 1.231722e-06, 1.264784e-06, 1.254392e-06, 1.280581e-06, 
    1.263163e-06, 1.284108e-06, 1.280077e-06, 1.292231e-06, 1.288743e-06, 
    1.304352e-06, 1.293842e-06, 1.312482e-06, 1.301838e-06, 1.3035e-06, 
    1.293495e-06, 1.234966e-06, 1.245863e-06, 1.234322e-06, 1.235872e-06, 
    1.235176e-06, 1.226734e-06, 1.22249e-06, 1.21363e-06, 1.215236e-06, 
    1.221745e-06, 1.236569e-06, 1.231526e-06, 1.244255e-06, 1.243967e-06, 
    1.258216e-06, 1.251781e-06, 1.275858e-06, 1.26899e-06, 1.288888e-06, 
    1.283868e-06, 1.288651e-06, 1.2872e-06, 1.28867e-06, 1.281313e-06, 
    1.284462e-06, 1.277998e-06, 1.252986e-06, 1.260311e-06, 1.23853e-06, 
    1.225528e-06, 1.216933e-06, 1.210853e-06, 1.211711e-06, 1.213349e-06, 
    1.221783e-06, 1.229741e-06, 1.235823e-06, 1.239901e-06, 1.243925e-06, 
    1.256147e-06, 1.262642e-06, 1.277248e-06, 1.274606e-06, 1.279084e-06, 
    1.283369e-06, 1.290581e-06, 1.289393e-06, 1.292575e-06, 1.278965e-06, 
    1.288001e-06, 1.273101e-06, 1.277167e-06, 1.24502e-06, 1.232886e-06, 
    1.227746e-06, 1.223257e-06, 1.212371e-06, 1.219883e-06, 1.216919e-06, 
    1.223977e-06, 1.228473e-06, 1.226248e-06, 1.240012e-06, 1.234651e-06, 
    1.263028e-06, 1.250764e-06, 1.282869e-06, 1.275148e-06, 1.284723e-06, 
    1.279833e-06, 1.288218e-06, 1.28067e-06, 1.29376e-06, 1.29662e-06, 
    1.294665e-06, 1.302182e-06, 1.280251e-06, 1.28865e-06, 1.226187e-06, 
    1.226549e-06, 1.22824e-06, 1.220817e-06, 1.220364e-06, 1.213585e-06, 
    1.219616e-06, 1.222189e-06, 1.228734e-06, 1.232613e-06, 1.236307e-06, 
    1.244449e-06, 1.253575e-06, 1.266395e-06, 1.275647e-06, 1.281869e-06, 
    1.278052e-06, 1.281421e-06, 1.277655e-06, 1.275891e-06, 1.295547e-06, 
    1.284491e-06, 1.301099e-06, 1.300177e-06, 1.292649e-06, 1.30028e-06, 
    1.226804e-06, 1.224717e-06, 1.217487e-06, 1.223143e-06, 1.212848e-06, 
    1.218605e-06, 1.221921e-06, 1.234763e-06, 1.237594e-06, 1.240222e-06, 
    1.24542e-06, 1.252109e-06, 1.263887e-06, 1.274182e-06, 1.283618e-06, 
    1.282926e-06, 1.283169e-06, 1.285282e-06, 1.280052e-06, 1.286141e-06, 
    1.287164e-06, 1.284489e-06, 1.300053e-06, 1.295597e-06, 1.300157e-06, 
    1.297254e-06, 1.225395e-06, 1.228908e-06, 1.227009e-06, 1.230581e-06, 
    1.228063e-06, 1.239276e-06, 1.242648e-06, 1.258491e-06, 1.251977e-06, 
    1.262353e-06, 1.253029e-06, 1.254678e-06, 1.262691e-06, 1.253531e-06, 
    1.273612e-06, 1.259979e-06, 1.285364e-06, 1.271683e-06, 1.286223e-06, 
    1.283576e-06, 1.28796e-06, 1.291892e-06, 1.296848e-06, 1.306018e-06, 
    1.303891e-06, 1.31158e-06, 1.234155e-06, 1.238728e-06, 1.238326e-06, 
    1.243121e-06, 1.246674e-06, 1.254393e-06, 1.266826e-06, 1.262143e-06, 
    1.270746e-06, 1.272477e-06, 1.259409e-06, 1.267424e-06, 1.241793e-06, 
    1.245915e-06, 1.24346e-06, 1.234513e-06, 1.263219e-06, 1.248444e-06, 
    1.275799e-06, 1.267741e-06, 1.29133e-06, 1.27957e-06, 1.302721e-06, 
    1.312684e-06, 1.322097e-06, 1.33314e-06, 1.241229e-06, 1.238116e-06, 
    1.243692e-06, 1.251428e-06, 1.258628e-06, 1.268234e-06, 1.269219e-06, 
    1.271023e-06, 1.275703e-06, 1.279646e-06, 1.271593e-06, 1.280634e-06, 
    1.246872e-06, 1.264506e-06, 1.236938e-06, 1.245206e-06, 1.250969e-06, 
    1.24844e-06, 1.261606e-06, 1.26472e-06, 1.277414e-06, 1.270844e-06, 
    1.31022e-06, 1.292722e-06, 1.341582e-06, 1.327832e-06, 1.23703e-06, 
    1.241218e-06, 1.255851e-06, 1.248878e-06, 1.268876e-06, 1.273824e-06, 
    1.277854e-06, 1.283015e-06, 1.283572e-06, 1.286636e-06, 1.281617e-06, 
    1.286437e-06, 1.268253e-06, 1.276362e-06, 1.254173e-06, 1.259555e-06, 
    1.257077e-06, 1.254363e-06, 1.26275e-06, 1.271718e-06, 1.27191e-06, 
    1.274793e-06, 1.282933e-06, 1.268955e-06, 1.312486e-06, 1.285511e-06, 
    1.245793e-06, 1.253896e-06, 1.255056e-06, 1.251912e-06, 1.273327e-06, 
    1.265546e-06, 1.286561e-06, 1.280864e-06, 1.290206e-06, 1.285559e-06, 
    1.284876e-06, 1.278922e-06, 1.275222e-06, 1.265901e-06, 1.258342e-06, 
    1.252366e-06, 1.253754e-06, 1.260324e-06, 1.272267e-06, 1.283621e-06, 
    1.281129e-06, 1.289493e-06, 1.267418e-06, 1.27665e-06, 1.273077e-06, 
    1.282403e-06, 1.262018e-06, 1.279367e-06, 1.257603e-06, 1.259503e-06, 
    1.265391e-06, 1.277279e-06, 1.279917e-06, 1.282737e-06, 1.280996e-06, 
    1.272572e-06, 1.271195e-06, 1.265247e-06, 1.263607e-06, 1.259088e-06, 
    1.255352e-06, 1.258765e-06, 1.262353e-06, 1.272575e-06, 1.281823e-06, 
    1.291946e-06, 1.29443e-06, 1.306321e-06, 1.296636e-06, 1.312637e-06, 
    1.299025e-06, 1.322634e-06, 1.280377e-06, 1.29863e-06, 1.26566e-06, 
    1.26919e-06, 1.275589e-06, 1.290329e-06, 1.282361e-06, 1.291682e-06, 
    1.271141e-06, 1.260551e-06, 1.257819e-06, 1.252729e-06, 1.257935e-06, 
    1.257511e-06, 1.262502e-06, 1.260897e-06, 1.272915e-06, 1.266452e-06, 
    1.284856e-06, 1.291607e-06, 1.310771e-06, 1.322592e-06, 1.334682e-06, 
    1.340038e-06, 1.34167e-06, 1.342352e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  7.62962e-06, 7.663833e-06, 7.657164e-06, 7.684774e-06, 7.66945e-06, 
    7.687516e-06, 7.636518e-06, 7.66513e-06, 7.646854e-06, 7.632637e-06, 
    7.738333e-06, 7.685942e-06, 7.792898e-06, 7.759395e-06, 7.843597e-06, 
    7.787654e-06, 7.854883e-06, 7.841975e-06, 7.880833e-06, 7.869683e-06, 
    7.919392e-06, 7.885952e-06, 7.945202e-06, 7.911397e-06, 7.916667e-06, 
    7.884806e-06, 7.696551e-06, 7.731862e-06, 7.69444e-06, 7.699475e-06, 
    7.697209e-06, 7.669728e-06, 7.655881e-06, 7.626941e-06, 7.632183e-06, 
    7.653437e-06, 7.70168e-06, 7.685288e-06, 7.7266e-06, 7.725669e-06, 
    7.771707e-06, 7.750935e-06, 7.828442e-06, 7.806382e-06, 7.870139e-06, 
    7.854078e-06, 7.869366e-06, 7.864717e-06, 7.869403e-06, 7.845872e-06, 
    7.855933e-06, 7.83524e-06, 7.754918e-06, 7.778539e-06, 7.708093e-06, 
    7.665777e-06, 7.637736e-06, 7.617852e-06, 7.620644e-06, 7.626002e-06, 
    7.653545e-06, 7.679474e-06, 7.69925e-06, 7.712473e-06, 7.725511e-06, 
    7.765004e-06, 7.785947e-06, 7.832876e-06, 7.824408e-06, 7.838745e-06, 
    7.852473e-06, 7.875509e-06, 7.871713e-06, 7.881856e-06, 7.838332e-06, 
    7.867242e-06, 7.819513e-06, 7.832556e-06, 7.729092e-06, 7.689746e-06, 
    7.672996e-06, 7.65837e-06, 7.622798e-06, 7.647351e-06, 7.637659e-06, 
    7.660695e-06, 7.675338e-06, 7.668083e-06, 7.712826e-06, 7.695407e-06, 
    7.787176e-06, 7.747614e-06, 7.850882e-06, 7.826128e-06, 7.856793e-06, 
    7.84114e-06, 7.867944e-06, 7.843806e-06, 7.885624e-06, 7.894736e-06, 
    7.88849e-06, 7.912437e-06, 7.842415e-06, 7.869278e-06, 7.667925e-06, 
    7.669108e-06, 7.674605e-06, 7.650387e-06, 7.648907e-06, 7.626746e-06, 
    7.646447e-06, 7.654842e-06, 7.676169e-06, 7.688775e-06, 7.700769e-06, 
    7.72718e-06, 7.75668e-06, 7.797995e-06, 7.827722e-06, 7.84765e-06, 
    7.835421e-06, 7.846201e-06, 7.83413e-06, 7.828466e-06, 7.891294e-06, 
    7.855992e-06, 7.908968e-06, 7.906036e-06, 7.882031e-06, 7.906344e-06, 
    7.669922e-06, 7.663112e-06, 7.639507e-06, 7.657964e-06, 7.624319e-06, 
    7.643137e-06, 7.653946e-06, 7.695749e-06, 7.704944e-06, 7.71347e-06, 
    7.730312e-06, 7.751934e-06, 7.789917e-06, 7.822998e-06, 7.85324e-06, 
    7.851011e-06, 7.851788e-06, 7.85853e-06, 7.84179e-06, 7.861262e-06, 
    7.864518e-06, 7.855972e-06, 7.905619e-06, 7.891425e-06, 7.905941e-06, 
    7.896686e-06, 7.665313e-06, 7.676741e-06, 7.670547e-06, 7.682174e-06, 
    7.673962e-06, 7.710403e-06, 7.721325e-06, 7.772536e-06, 7.751506e-06, 
    7.784981e-06, 7.754892e-06, 7.760217e-06, 7.786025e-06, 7.756498e-06, 
    7.821137e-06, 7.777266e-06, 7.858783e-06, 7.814904e-06, 7.861517e-06, 
    7.853042e-06, 7.867047e-06, 7.879601e-06, 7.89539e-06, 7.924562e-06, 
    7.917789e-06, 7.942207e-06, 7.693799e-06, 7.708634e-06, 7.707333e-06, 
    7.722871e-06, 7.734366e-06, 7.759329e-06, 7.799381e-06, 7.784301e-06, 
    7.811968e-06, 7.817525e-06, 7.775465e-06, 7.801265e-06, 7.718498e-06, 
    7.731832e-06, 7.723888e-06, 7.694839e-06, 7.78769e-06, 7.739985e-06, 
    7.828112e-06, 7.802225e-06, 7.877786e-06, 7.840174e-06, 7.914063e-06, 
    7.945681e-06, 7.975496e-06, 8.010316e-06, 7.716741e-06, 7.706636e-06, 
    7.724708e-06, 7.749729e-06, 7.772967e-06, 7.8039e-06, 7.807061e-06, 
    7.812843e-06, 7.82786e-06, 7.840498e-06, 7.814647e-06, 7.843643e-06, 
    7.7349e-06, 7.791836e-06, 7.702704e-06, 7.729504e-06, 7.748142e-06, 
    7.739968e-06, 7.782474e-06, 7.792487e-06, 7.833243e-06, 7.81217e-06, 
    7.937842e-06, 7.882179e-06, 8.036875e-06, 7.99357e-06, 7.703098e-06, 
    7.716677e-06, 7.763999e-06, 7.741472e-06, 7.805947e-06, 7.821838e-06, 
    7.834751e-06, 7.851274e-06, 7.853047e-06, 7.862844e-06, 7.846776e-06, 
    7.862197e-06, 7.803877e-06, 7.829922e-06, 7.758506e-06, 7.775853e-06, 
    7.767866e-06, 7.759091e-06, 7.78613e-06, 7.814959e-06, 7.815579e-06, 
    7.824812e-06, 7.85085e-06, 7.806057e-06, 7.944974e-06, 7.859075e-06, 
    7.731493e-06, 7.757667e-06, 7.761417e-06, 7.751268e-06, 7.82022e-06, 
    7.795214e-06, 7.862606e-06, 7.844366e-06, 7.874229e-06, 7.859382e-06, 
    7.857178e-06, 7.838124e-06, 7.826242e-06, 7.796291e-06, 7.771928e-06, 
    7.752645e-06, 7.757111e-06, 7.778301e-06, 7.816702e-06, 7.853101e-06, 
    7.845111e-06, 7.871855e-06, 7.801097e-06, 7.830738e-06, 7.819257e-06, 
    7.849161e-06, 7.783862e-06, 7.839561e-06, 7.769627e-06, 7.775742e-06, 
    7.794693e-06, 7.832864e-06, 7.84132e-06, 7.850343e-06, 7.844761e-06, 
    7.817742e-06, 7.813313e-06, 7.794182e-06, 7.788886e-06, 7.774335e-06, 
    7.762265e-06, 7.773275e-06, 7.784816e-06, 7.817694e-06, 7.84733e-06, 
    7.879676e-06, 7.887601e-06, 7.925402e-06, 7.894592e-06, 7.945408e-06, 
    7.902154e-06, 7.977059e-06, 7.84279e-06, 7.901083e-06, 7.795563e-06, 
    7.806905e-06, 7.827432e-06, 7.874589e-06, 7.849121e-06, 7.878903e-06, 
    7.813136e-06, 7.779038e-06, 7.770233e-06, 7.753802e-06, 7.770593e-06, 
    7.769228e-06, 7.785307e-06, 7.780124e-06, 7.818763e-06, 7.797999e-06, 
    7.85701e-06, 7.878574e-06, 7.939547e-06, 7.976959e-06, 8.015115e-06, 
    8.031952e-06, 8.037081e-06, 8.039216e-06,
  3.976129e-06, 4.006499e-06, 4.00059e-06, 4.025133e-06, 4.011514e-06, 
    4.027592e-06, 3.982283e-06, 4.007704e-06, 3.99147e-06, 3.978864e-06, 
    4.072916e-06, 4.026229e-06, 4.121659e-06, 4.091719e-06, 4.167096e-06, 
    4.116991e-06, 4.177228e-06, 4.165655e-06, 4.200542e-06, 4.190537e-06, 
    4.235262e-06, 4.205163e-06, 4.258528e-06, 4.228071e-06, 4.232827e-06, 
    4.20417e-06, 4.035615e-06, 4.06709e-06, 4.033751e-06, 4.038234e-06, 
    4.036224e-06, 4.011792e-06, 3.999497e-06, 3.973817e-06, 3.978475e-06, 
    3.997342e-06, 4.04025e-06, 4.02567e-06, 4.062469e-06, 4.061636e-06, 
    4.102747e-06, 4.084191e-06, 4.153529e-06, 4.133779e-06, 4.190954e-06, 
    4.176547e-06, 4.190276e-06, 4.186112e-06, 4.19033e-06, 4.169207e-06, 
    4.178252e-06, 4.159686e-06, 4.087663e-06, 4.108778e-06, 4.045921e-06, 
    4.008294e-06, 3.983395e-06, 3.965757e-06, 3.968249e-06, 3.972999e-06, 
    3.997452e-06, 4.020503e-06, 4.038101e-06, 4.049889e-06, 4.061516e-06, 
    4.096772e-06, 4.115496e-06, 4.157524e-06, 4.149933e-06, 4.1628e-06, 
    4.175115e-06, 4.195812e-06, 4.192404e-06, 4.20153e-06, 4.162465e-06, 
    4.18841e-06, 4.145611e-06, 4.157299e-06, 4.064656e-06, 4.029602e-06, 
    4.014717e-06, 4.001725e-06, 3.970164e-06, 3.991948e-06, 3.983354e-06, 
    4.003815e-06, 4.016833e-06, 4.010394e-06, 4.050211e-06, 4.034712e-06, 
    4.116606e-06, 4.081255e-06, 4.173678e-06, 4.151491e-06, 4.179003e-06, 
    4.164957e-06, 4.189033e-06, 4.167362e-06, 4.204931e-06, 4.213125e-06, 
    4.207524e-06, 4.229063e-06, 4.166162e-06, 4.190274e-06, 4.010212e-06, 
    4.011262e-06, 4.016157e-06, 3.994656e-06, 3.993343e-06, 3.973688e-06, 
    3.991177e-06, 3.998633e-06, 4.017591e-06, 4.028816e-06, 4.0395e-06, 
    4.063029e-06, 4.089365e-06, 4.126307e-06, 4.152928e-06, 4.170808e-06, 
    4.159842e-06, 4.169523e-06, 4.158701e-06, 4.153633e-06, 4.210052e-06, 
    4.178335e-06, 4.225963e-06, 4.223323e-06, 4.201746e-06, 4.22362e-06, 
    4.012e-06, 4.005959e-06, 3.985003e-06, 4.001399e-06, 3.97155e-06, 
    3.988244e-06, 3.997854e-06, 4.035031e-06, 4.043222e-06, 4.050816e-06, 
    4.065836e-06, 4.08514e-06, 4.119086e-06, 4.148713e-06, 4.175833e-06, 
    4.173844e-06, 4.174544e-06, 4.180607e-06, 4.165589e-06, 4.183075e-06, 
    4.18601e-06, 4.178334e-06, 4.222969e-06, 4.2102e-06, 4.223266e-06, 
    4.214951e-06, 4.007923e-06, 4.018093e-06, 4.012596e-06, 4.022934e-06, 
    4.015647e-06, 4.048079e-06, 4.057822e-06, 4.103538e-06, 4.084759e-06, 
    4.114668e-06, 4.087795e-06, 4.09255e-06, 4.115635e-06, 4.089247e-06, 
    4.147073e-06, 4.107826e-06, 4.180843e-06, 4.141521e-06, 4.183312e-06, 
    4.175715e-06, 4.188298e-06, 4.199576e-06, 4.213786e-06, 4.240045e-06, 
    4.23396e-06, 4.255959e-06, 4.033275e-06, 4.046498e-06, 4.045338e-06, 
    4.059195e-06, 4.069454e-06, 4.09173e-06, 4.127549e-06, 4.114067e-06, 
    4.138835e-06, 4.143812e-06, 4.106192e-06, 4.129271e-06, 4.05536e-06, 
    4.067263e-06, 4.060178e-06, 4.034315e-06, 4.117166e-06, 4.074563e-06, 
    4.153368e-06, 4.130191e-06, 4.197967e-06, 4.164205e-06, 4.230611e-06, 
    4.259105e-06, 4.28601e-06, 4.317503e-06, 4.053727e-06, 4.044733e-06, 
    4.060846e-06, 4.08317e-06, 4.103938e-06, 4.131603e-06, 4.13444e-06, 
    4.139631e-06, 4.153093e-06, 4.164422e-06, 4.141268e-06, 4.167264e-06, 
    4.070016e-06, 4.120874e-06, 4.041331e-06, 4.065215e-06, 4.081855e-06, 
    4.074557e-06, 4.112529e-06, 4.121496e-06, 4.15801e-06, 4.139122e-06, 
    4.252062e-06, 4.201954e-06, 4.341555e-06, 4.302371e-06, 4.041592e-06, 
    4.053698e-06, 4.095932e-06, 4.075817e-06, 4.133455e-06, 4.147687e-06, 
    4.159275e-06, 4.174097e-06, 4.175702e-06, 4.184495e-06, 4.170089e-06, 
    4.183928e-06, 4.131662e-06, 4.154988e-06, 4.091102e-06, 4.106614e-06, 
    4.099476e-06, 4.09165e-06, 4.115824e-06, 4.141631e-06, 4.14219e-06, 
    4.150477e-06, 4.173849e-06, 4.133689e-06, 4.258531e-06, 4.181255e-06, 
    4.066914e-06, 4.09029e-06, 4.093642e-06, 4.084577e-06, 4.146259e-06, 
    4.123868e-06, 4.184282e-06, 4.167923e-06, 4.194741e-06, 4.181406e-06, 
    4.179445e-06, 4.162346e-06, 4.151712e-06, 4.124892e-06, 4.103121e-06, 
    4.085892e-06, 4.089896e-06, 4.108831e-06, 4.143213e-06, 4.175844e-06, 
    4.168687e-06, 4.192701e-06, 4.129265e-06, 4.155817e-06, 4.145544e-06, 
    4.172351e-06, 4.113707e-06, 4.163603e-06, 4.100988e-06, 4.106465e-06, 
    4.123424e-06, 4.157615e-06, 4.165205e-06, 4.173301e-06, 4.168306e-06, 
    4.144089e-06, 4.140129e-06, 4.123013e-06, 4.118288e-06, 4.105273e-06, 
    4.094505e-06, 4.10434e-06, 4.114678e-06, 4.144102e-06, 4.170682e-06, 
    4.199736e-06, 4.20686e-06, 4.240905e-06, 4.213173e-06, 4.258961e-06, 
    4.220005e-06, 4.287532e-06, 4.166512e-06, 4.218877e-06, 4.124199e-06, 
    4.134362e-06, 4.15276e-06, 4.195088e-06, 4.172224e-06, 4.198972e-06, 
    4.139975e-06, 4.109481e-06, 4.101614e-06, 4.086937e-06, 4.10195e-06, 
    4.100728e-06, 4.115112e-06, 4.110488e-06, 4.14508e-06, 4.126486e-06, 
    4.179394e-06, 4.198762e-06, 4.253649e-06, 4.28742e-06, 4.321911e-06, 
    4.337166e-06, 4.341813e-06, 4.343756e-06,
  3.78041e-06, 3.813993e-06, 3.807456e-06, 3.834614e-06, 3.81954e-06, 
    3.837337e-06, 3.78721e-06, 3.815328e-06, 3.797368e-06, 3.78343e-06, 
    3.887551e-06, 3.835828e-06, 3.94161e-06, 3.908388e-06, 3.992074e-06, 
    3.936429e-06, 4.003335e-06, 3.990468e-06, 4.029258e-06, 4.018129e-06, 
    4.067907e-06, 4.034398e-06, 4.093818e-06, 4.059896e-06, 4.065193e-06, 
    4.033294e-06, 3.846217e-06, 3.881094e-06, 3.844154e-06, 3.849118e-06, 
    3.846891e-06, 3.81985e-06, 3.806251e-06, 3.777851e-06, 3.783001e-06, 
    3.803865e-06, 3.851351e-06, 3.835206e-06, 3.87596e-06, 3.875038e-06, 
    3.920619e-06, 3.900039e-06, 3.976995e-06, 3.955059e-06, 4.018593e-06, 
    4.002574e-06, 4.01784e-06, 4.013209e-06, 4.0179e-06, 3.994417e-06, 
    4.004471e-06, 3.983835e-06, 3.903889e-06, 3.927311e-06, 3.85763e-06, 
    3.815984e-06, 3.78844e-06, 3.768944e-06, 3.771698e-06, 3.776949e-06, 
    3.803987e-06, 3.829487e-06, 3.848968e-06, 3.862023e-06, 3.874905e-06, 
    3.914e-06, 3.934769e-06, 3.981435e-06, 3.973e-06, 3.987298e-06, 
    4.000982e-06, 4.023997e-06, 4.020206e-06, 4.030358e-06, 3.986923e-06, 
    4.015767e-06, 3.968197e-06, 3.981183e-06, 3.878397e-06, 3.839559e-06, 
    3.823091e-06, 3.808711e-06, 3.773815e-06, 3.797898e-06, 3.788396e-06, 
    3.811022e-06, 3.825427e-06, 3.8183e-06, 3.86238e-06, 3.845217e-06, 
    3.936001e-06, 3.896786e-06, 3.999385e-06, 3.974731e-06, 4.005304e-06, 
    3.989692e-06, 4.016458e-06, 3.992365e-06, 4.034141e-06, 4.04326e-06, 
    4.037027e-06, 4.060998e-06, 3.991031e-06, 4.017838e-06, 3.818099e-06, 
    3.819261e-06, 3.824678e-06, 3.800893e-06, 3.799441e-06, 3.777709e-06, 
    3.797045e-06, 3.805291e-06, 3.826263e-06, 3.838689e-06, 3.850519e-06, 
    3.876583e-06, 3.905779e-06, 3.946765e-06, 3.976327e-06, 3.996194e-06, 
    3.984008e-06, 3.994766e-06, 3.98274e-06, 3.977109e-06, 4.039841e-06, 
    4.004564e-06, 4.057546e-06, 4.054607e-06, 4.030599e-06, 4.054938e-06, 
    3.820077e-06, 3.813393e-06, 3.790218e-06, 3.808349e-06, 3.775346e-06, 
    3.793803e-06, 3.804432e-06, 3.845572e-06, 3.85464e-06, 3.863052e-06, 
    3.879692e-06, 3.901092e-06, 3.938751e-06, 3.971646e-06, 4.001779e-06, 
    3.999568e-06, 4.000347e-06, 4.007089e-06, 3.990395e-06, 4.009833e-06, 
    4.013097e-06, 4.004562e-06, 4.054214e-06, 4.040002e-06, 4.054545e-06, 
    4.045289e-06, 3.815565e-06, 3.826819e-06, 3.820736e-06, 3.832178e-06, 
    3.824115e-06, 3.860023e-06, 3.870817e-06, 3.9215e-06, 3.900669e-06, 
    3.933848e-06, 3.904035e-06, 3.90931e-06, 3.934927e-06, 3.905644e-06, 
    3.969827e-06, 3.92626e-06, 4.007351e-06, 3.963663e-06, 4.010095e-06, 
    4.001649e-06, 4.015639e-06, 4.028184e-06, 4.043994e-06, 4.073228e-06, 
    4.066451e-06, 4.090953e-06, 3.843625e-06, 3.85827e-06, 3.856982e-06, 
    3.872334e-06, 3.883703e-06, 3.908399e-06, 3.948143e-06, 3.933179e-06, 
    3.960673e-06, 3.966202e-06, 3.924439e-06, 3.950056e-06, 3.868087e-06, 
    3.881278e-06, 3.873423e-06, 3.844778e-06, 3.936621e-06, 3.88937e-06, 
    3.976816e-06, 3.951077e-06, 4.026394e-06, 3.98886e-06, 4.062722e-06, 
    4.094465e-06, 4.124448e-06, 4.159587e-06, 3.866276e-06, 3.856313e-06, 
    3.874162e-06, 3.898911e-06, 3.921941e-06, 3.952644e-06, 3.955793e-06, 
    3.961557e-06, 3.976509e-06, 3.989097e-06, 3.963378e-06, 3.992256e-06, 
    3.884335e-06, 3.940735e-06, 3.852547e-06, 3.879009e-06, 3.897451e-06, 
    3.889359e-06, 3.93147e-06, 3.941423e-06, 3.981975e-06, 3.960991e-06, 
    4.086618e-06, 4.030833e-06, 4.186435e-06, 4.142701e-06, 3.852834e-06, 
    3.866243e-06, 3.913062e-06, 3.890756e-06, 3.954699e-06, 3.970506e-06, 
    3.983377e-06, 3.999852e-06, 4.001635e-06, 4.011412e-06, 3.995395e-06, 
    4.01078e-06, 3.952709e-06, 3.978616e-06, 3.907701e-06, 3.924909e-06, 
    3.91699e-06, 3.908309e-06, 3.935128e-06, 3.963782e-06, 3.964399e-06, 
    3.973606e-06, 3.999591e-06, 3.954959e-06, 4.093834e-06, 4.007822e-06, 
    3.880887e-06, 3.906807e-06, 3.91052e-06, 3.900466e-06, 3.968919e-06, 
    3.944057e-06, 4.011174e-06, 3.992988e-06, 4.022805e-06, 4.007976e-06, 
    4.005796e-06, 3.98679e-06, 3.974976e-06, 3.945195e-06, 3.921034e-06, 
    3.901924e-06, 3.906364e-06, 3.92737e-06, 3.965538e-06, 4.001794e-06, 
    3.99384e-06, 4.020535e-06, 3.950047e-06, 3.979538e-06, 3.968127e-06, 
    3.99791e-06, 3.93278e-06, 3.9882e-06, 3.918666e-06, 3.924742e-06, 
    3.943564e-06, 3.981539e-06, 3.989967e-06, 3.998968e-06, 3.993413e-06, 
    3.96651e-06, 3.962112e-06, 3.943107e-06, 3.937865e-06, 3.923419e-06, 
    3.911475e-06, 3.922386e-06, 3.933858e-06, 3.966523e-06, 3.996056e-06, 
    4.028363e-06, 4.036287e-06, 4.074193e-06, 4.043319e-06, 4.094315e-06, 
    4.050933e-06, 4.126156e-06, 3.991428e-06, 4.049668e-06, 3.944423e-06, 
    3.955705e-06, 3.976143e-06, 4.023197e-06, 3.997769e-06, 4.027515e-06, 
    3.96194e-06, 3.928093e-06, 3.919361e-06, 3.903084e-06, 3.919734e-06, 
    3.918379e-06, 3.934337e-06, 3.929206e-06, 3.96761e-06, 3.946961e-06, 
    4.005741e-06, 4.027281e-06, 4.088381e-06, 4.126025e-06, 4.1645e-06, 
    4.181531e-06, 4.186721e-06, 4.188891e-06,
  3.868069e-06, 3.904865e-06, 3.897699e-06, 3.927474e-06, 3.910944e-06, 
    3.93046e-06, 3.875516e-06, 3.906329e-06, 3.886645e-06, 3.871375e-06, 
    3.985568e-06, 3.928805e-06, 4.04495e-06, 4.008443e-06, 4.100456e-06, 
    4.039258e-06, 4.11285e-06, 4.098686e-06, 4.14139e-06, 4.129135e-06, 
    4.183986e-06, 4.147053e-06, 4.212558e-06, 4.175152e-06, 4.180993e-06, 
    4.145837e-06, 3.940198e-06, 3.978479e-06, 3.937935e-06, 3.943382e-06, 
    3.940937e-06, 3.911285e-06, 3.896382e-06, 3.865264e-06, 3.870904e-06, 
    3.893765e-06, 3.945832e-06, 3.928121e-06, 3.972833e-06, 3.971821e-06, 
    4.021879e-06, 3.999271e-06, 4.083861e-06, 4.059733e-06, 4.129646e-06, 
    4.112009e-06, 4.128816e-06, 4.123717e-06, 4.128883e-06, 4.103032e-06, 
    4.114098e-06, 4.091386e-06, 4.003501e-06, 4.029233e-06, 3.95272e-06, 
    3.907053e-06, 3.876864e-06, 3.85551e-06, 3.858526e-06, 3.864277e-06, 
    3.893899e-06, 3.92185e-06, 3.943215e-06, 3.957538e-06, 3.971675e-06, 
    4.014613e-06, 4.037431e-06, 4.088748e-06, 4.079465e-06, 4.095198e-06, 
    4.110257e-06, 4.135597e-06, 4.131422e-06, 4.142604e-06, 4.094783e-06, 
    4.126535e-06, 4.074181e-06, 4.088468e-06, 3.975519e-06, 3.932895e-06, 
    3.914842e-06, 3.899076e-06, 3.860845e-06, 3.887227e-06, 3.876817e-06, 
    3.901606e-06, 3.917397e-06, 3.909584e-06, 3.95793e-06, 3.9391e-06, 
    4.038785e-06, 3.9957e-06, 4.108499e-06, 4.081369e-06, 4.115014e-06, 
    4.09783e-06, 4.127296e-06, 4.100772e-06, 4.14677e-06, 4.156818e-06, 
    4.149951e-06, 4.176364e-06, 4.099304e-06, 4.128816e-06, 3.909365e-06, 
    3.910638e-06, 3.916576e-06, 3.890509e-06, 3.888917e-06, 3.865109e-06, 
    3.88629e-06, 3.895327e-06, 3.918314e-06, 3.931941e-06, 3.944916e-06, 
    3.973517e-06, 4.005577e-06, 4.050617e-06, 4.083126e-06, 4.104986e-06, 
    4.091575e-06, 4.103414e-06, 4.09018e-06, 4.083985e-06, 4.153052e-06, 
    4.114201e-06, 4.17256e-06, 4.169321e-06, 4.14287e-06, 4.169685e-06, 
    3.911533e-06, 3.904205e-06, 3.878812e-06, 3.898677e-06, 3.86252e-06, 
    3.882739e-06, 3.894387e-06, 3.939492e-06, 3.949437e-06, 3.958668e-06, 
    3.97693e-06, 4.000427e-06, 4.041807e-06, 4.077978e-06, 4.111133e-06, 
    4.1087e-06, 4.109557e-06, 4.116979e-06, 4.098604e-06, 4.12e-06, 
    4.123596e-06, 4.114197e-06, 4.168886e-06, 4.153227e-06, 4.169251e-06, 
    4.159052e-06, 3.906586e-06, 3.918925e-06, 3.912255e-06, 3.924802e-06, 
    3.91596e-06, 3.955347e-06, 3.967193e-06, 4.02285e-06, 3.999964e-06, 
    4.036418e-06, 4.00366e-06, 4.009455e-06, 4.037609e-06, 4.005427e-06, 
    4.075979e-06, 4.028081e-06, 4.117268e-06, 4.069202e-06, 4.120289e-06, 
    4.11099e-06, 4.126392e-06, 4.14021e-06, 4.157625e-06, 4.18985e-06, 
    4.182377e-06, 4.209396e-06, 3.937354e-06, 3.953422e-06, 3.952007e-06, 
    3.968853e-06, 3.981334e-06, 4.008452e-06, 4.05213e-06, 4.035679e-06, 
    4.065906e-06, 4.071987e-06, 4.026075e-06, 4.054234e-06, 3.964194e-06, 
    3.978675e-06, 3.97005e-06, 3.93862e-06, 4.039466e-06, 3.987558e-06, 
    4.083663e-06, 4.055355e-06, 4.138238e-06, 4.096918e-06, 4.178266e-06, 
    4.213275e-06, 4.246354e-06, 4.285165e-06, 3.962205e-06, 3.951272e-06, 
    3.970859e-06, 3.998035e-06, 4.023331e-06, 4.057079e-06, 4.06054e-06, 
    4.06688e-06, 4.083324e-06, 4.097175e-06, 4.068885e-06, 4.100651e-06, 
    3.982036e-06, 4.043987e-06, 3.947142e-06, 3.976184e-06, 3.996431e-06, 
    3.987544e-06, 4.033801e-06, 4.04474e-06, 4.089341e-06, 4.066256e-06, 
    4.20462e-06, 4.14313e-06, 4.314832e-06, 4.266512e-06, 3.947456e-06, 
    3.962168e-06, 4.013577e-06, 3.989077e-06, 4.059337e-06, 4.076721e-06, 
    4.090881e-06, 4.109014e-06, 4.110975e-06, 4.121739e-06, 4.104107e-06, 
    4.121042e-06, 4.057151e-06, 4.085643e-06, 4.007685e-06, 4.026593e-06, 
    4.017889e-06, 4.008353e-06, 4.037821e-06, 4.069329e-06, 4.070004e-06, 
    4.080133e-06, 4.108738e-06, 4.059623e-06, 4.212587e-06, 4.117798e-06, 
    3.978241e-06, 4.006708e-06, 4.010783e-06, 3.999739e-06, 4.074977e-06, 
    4.047637e-06, 4.121477e-06, 4.101458e-06, 4.134284e-06, 4.117956e-06, 
    4.115556e-06, 4.094637e-06, 4.081639e-06, 4.048889e-06, 4.022335e-06, 
    4.00134e-06, 4.006217e-06, 4.029297e-06, 4.07126e-06, 4.111152e-06, 
    4.102397e-06, 4.131784e-06, 4.054223e-06, 4.086659e-06, 4.074107e-06, 
    4.106875e-06, 4.035242e-06, 4.0962e-06, 4.019731e-06, 4.026408e-06, 
    4.047095e-06, 4.088863e-06, 4.098133e-06, 4.10804e-06, 4.101926e-06, 
    4.072328e-06, 4.06749e-06, 4.046592e-06, 4.040831e-06, 4.024954e-06, 
    4.011831e-06, 4.02382e-06, 4.036428e-06, 4.072341e-06, 4.104837e-06, 
    4.140406e-06, 4.149134e-06, 4.19092e-06, 4.156888e-06, 4.213117e-06, 
    4.165287e-06, 4.248252e-06, 4.099748e-06, 4.163885e-06, 4.048038e-06, 
    4.060444e-06, 4.082926e-06, 4.13472e-06, 4.106721e-06, 4.139475e-06, 
    4.0673e-06, 4.030094e-06, 4.020495e-06, 4.002614e-06, 4.020904e-06, 
    4.019415e-06, 4.036951e-06, 4.031312e-06, 4.073536e-06, 4.050829e-06, 
    4.115496e-06, 4.139216e-06, 4.20656e-06, 4.2481e-06, 4.290588e-06, 
    4.309409e-06, 4.315146e-06, 4.317545e-06,
  4.120389e-06, 4.15886e-06, 4.151365e-06, 4.182512e-06, 4.165217e-06, 
    4.185637e-06, 4.128171e-06, 4.160392e-06, 4.139806e-06, 4.123843e-06, 
    4.243343e-06, 4.183905e-06, 4.305588e-06, 4.267306e-06, 4.363847e-06, 
    4.29962e-06, 4.376864e-06, 4.361985e-06, 4.406853e-06, 4.393972e-06, 
    4.451656e-06, 4.412806e-06, 4.481728e-06, 4.442359e-06, 4.448505e-06, 
    4.411528e-06, 4.195826e-06, 4.235917e-06, 4.193458e-06, 4.19916e-06, 
    4.1966e-06, 4.165574e-06, 4.14999e-06, 4.117456e-06, 4.123351e-06, 
    4.147251e-06, 4.201725e-06, 4.183187e-06, 4.229994e-06, 4.228934e-06, 
    4.281391e-06, 4.257693e-06, 4.346419e-06, 4.321093e-06, 4.394509e-06, 
    4.375979e-06, 4.393638e-06, 4.388279e-06, 4.393708e-06, 4.366549e-06, 
    4.378173e-06, 4.354319e-06, 4.262126e-06, 4.289103e-06, 4.208935e-06, 
    4.161152e-06, 4.129582e-06, 4.107264e-06, 4.110415e-06, 4.116426e-06, 
    4.147392e-06, 4.176625e-06, 4.198983e-06, 4.213978e-06, 4.228782e-06, 
    4.273779e-06, 4.297702e-06, 4.351551e-06, 4.341803e-06, 4.358323e-06, 
    4.374137e-06, 4.400765e-06, 4.396376e-06, 4.40813e-06, 4.357886e-06, 
    4.391242e-06, 4.336256e-06, 4.351255e-06, 4.232817e-06, 4.188183e-06, 
    4.169299e-06, 4.152805e-06, 4.112839e-06, 4.140416e-06, 4.129532e-06, 
    4.15545e-06, 4.171968e-06, 4.163793e-06, 4.214388e-06, 4.194677e-06, 
    4.299122e-06, 4.253953e-06, 4.372291e-06, 4.343803e-06, 4.379136e-06, 
    4.361085e-06, 4.39204e-06, 4.364175e-06, 4.412509e-06, 4.423076e-06, 
    4.415854e-06, 4.443632e-06, 4.362633e-06, 4.393638e-06, 4.163565e-06, 
    4.164897e-06, 4.171108e-06, 4.143847e-06, 4.142182e-06, 4.117294e-06, 
    4.139435e-06, 4.148885e-06, 4.172926e-06, 4.187185e-06, 4.200765e-06, 
    4.230712e-06, 4.264304e-06, 4.311531e-06, 4.345646e-06, 4.368601e-06, 
    4.354516e-06, 4.36695e-06, 4.353053e-06, 4.346547e-06, 4.419115e-06, 
    4.378282e-06, 4.439631e-06, 4.436223e-06, 4.40841e-06, 4.436607e-06, 
    4.165833e-06, 4.158167e-06, 4.131617e-06, 4.152387e-06, 4.114589e-06, 
    4.135723e-06, 4.147903e-06, 4.195089e-06, 4.205496e-06, 4.215161e-06, 
    4.234286e-06, 4.258904e-06, 4.302289e-06, 4.340243e-06, 4.375058e-06, 
    4.372502e-06, 4.373402e-06, 4.3812e-06, 4.361899e-06, 4.384374e-06, 
    4.388153e-06, 4.378277e-06, 4.435766e-06, 4.419298e-06, 4.43615e-06, 
    4.425423e-06, 4.160658e-06, 4.173565e-06, 4.166588e-06, 4.179715e-06, 
    4.170465e-06, 4.211686e-06, 4.224091e-06, 4.282411e-06, 4.258419e-06, 
    4.296638e-06, 4.262292e-06, 4.268367e-06, 4.297891e-06, 4.264144e-06, 
    4.338146e-06, 4.287897e-06, 4.381503e-06, 4.331037e-06, 4.384678e-06, 
    4.374907e-06, 4.39109e-06, 4.405613e-06, 4.423922e-06, 4.457824e-06, 
    4.44996e-06, 4.478396e-06, 4.19285e-06, 4.20967e-06, 4.208187e-06, 
    4.225827e-06, 4.238901e-06, 4.267315e-06, 4.313118e-06, 4.29586e-06, 
    4.327571e-06, 4.333954e-06, 4.285789e-06, 4.315326e-06, 4.220949e-06, 
    4.236117e-06, 4.227081e-06, 4.194176e-06, 4.299835e-06, 4.245422e-06, 
    4.346211e-06, 4.316501e-06, 4.403541e-06, 4.36013e-06, 4.445634e-06, 
    4.482485e-06, 4.517323e-06, 4.558243e-06, 4.218866e-06, 4.207418e-06, 
    4.227927e-06, 4.2564e-06, 4.282913e-06, 4.318309e-06, 4.32194e-06, 
    4.328594e-06, 4.345854e-06, 4.360398e-06, 4.3307e-06, 4.364048e-06, 
    4.239641e-06, 4.304577e-06, 4.203096e-06, 4.233509e-06, 4.254718e-06, 
    4.245405e-06, 4.29389e-06, 4.305364e-06, 4.352173e-06, 4.327938e-06, 
    4.473375e-06, 4.408686e-06, 4.58954e-06, 4.538573e-06, 4.203423e-06, 
    4.218826e-06, 4.272688e-06, 4.247011e-06, 4.320678e-06, 4.338924e-06, 
    4.353788e-06, 4.372833e-06, 4.374891e-06, 4.386202e-06, 4.367677e-06, 
    4.385469e-06, 4.318385e-06, 4.348289e-06, 4.266511e-06, 4.286333e-06, 
    4.277207e-06, 4.26721e-06, 4.298107e-06, 4.331167e-06, 4.331873e-06, 
    4.342506e-06, 4.372554e-06, 4.320978e-06, 4.481768e-06, 4.38207e-06, 
    4.235659e-06, 4.26549e-06, 4.269758e-06, 4.258182e-06, 4.337092e-06, 
    4.308404e-06, 4.385925e-06, 4.364895e-06, 4.399383e-06, 4.382226e-06, 
    4.379705e-06, 4.357733e-06, 4.344085e-06, 4.309717e-06, 4.281869e-06, 
    4.25986e-06, 4.264972e-06, 4.289169e-06, 4.333193e-06, 4.375079e-06, 
    4.365884e-06, 4.396757e-06, 4.315312e-06, 4.349357e-06, 4.336181e-06, 
    4.370585e-06, 4.295403e-06, 4.359383e-06, 4.279137e-06, 4.286138e-06, 
    4.307836e-06, 4.351673e-06, 4.361404e-06, 4.371811e-06, 4.365387e-06, 
    4.334314e-06, 4.329234e-06, 4.307307e-06, 4.301265e-06, 4.284613e-06, 
    4.270856e-06, 4.283425e-06, 4.296648e-06, 4.334326e-06, 4.368445e-06, 
    4.40582e-06, 4.414994e-06, 4.458955e-06, 4.423153e-06, 4.482327e-06, 
    4.431993e-06, 4.519331e-06, 4.363105e-06, 4.430513e-06, 4.308824e-06, 
    4.321839e-06, 4.34544e-06, 4.399846e-06, 4.370424e-06, 4.404844e-06, 
    4.329036e-06, 4.290006e-06, 4.279939e-06, 4.261196e-06, 4.280368e-06, 
    4.278807e-06, 4.297195e-06, 4.291281e-06, 4.33558e-06, 4.311752e-06, 
    4.379642e-06, 4.404571e-06, 4.475412e-06, 4.519166e-06, 4.563958e-06, 
    4.583816e-06, 4.589871e-06, 4.592403e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.77824, 5.778221, 5.778224, 5.778209, 5.778217, 5.778207, 5.778236, 
    5.77822, 5.77823, 5.778238, 5.778179, 5.778208, 5.778149, 5.778167, 
    5.77812, 5.778152, 5.778114, 5.778121, 5.7781, 5.778106, 5.778078, 
    5.778097, 5.778064, 5.778082, 5.77808, 5.778097, 5.778203, 5.778183, 
    5.778203, 5.778201, 5.778202, 5.778217, 5.778225, 5.778241, 5.778238, 
    5.778226, 5.7782, 5.778209, 5.778185, 5.778186, 5.77816, 5.778172, 
    5.778129, 5.778141, 5.778105, 5.778114, 5.778106, 5.778108, 5.778106, 
    5.778119, 5.778113, 5.778125, 5.77817, 5.778156, 5.778196, 5.77822, 
    5.778235, 5.778246, 5.778245, 5.778242, 5.778226, 5.778212, 5.778201, 
    5.778193, 5.778186, 5.778164, 5.778152, 5.778126, 5.778131, 5.778123, 
    5.778115, 5.778102, 5.778104, 5.778099, 5.778123, 5.778107, 5.778133, 
    5.778126, 5.778184, 5.778206, 5.778215, 5.778224, 5.778244, 5.77823, 
    5.778235, 5.778223, 5.778214, 5.778218, 5.778193, 5.778203, 5.778152, 
    5.778174, 5.778116, 5.77813, 5.778113, 5.778121, 5.778107, 5.77812, 
    5.778097, 5.778091, 5.778095, 5.778082, 5.778121, 5.778106, 5.778218, 
    5.778218, 5.778214, 5.778228, 5.778229, 5.778242, 5.77823, 5.778226, 
    5.778214, 5.778207, 5.7782, 5.778185, 5.778169, 5.778145, 5.778129, 
    5.778118, 5.778125, 5.778119, 5.778125, 5.778129, 5.778093, 5.778113, 
    5.778084, 5.778085, 5.778099, 5.778085, 5.778217, 5.778221, 5.778234, 
    5.778224, 5.778243, 5.778232, 5.778226, 5.778203, 5.778198, 5.778193, 
    5.778183, 5.778171, 5.77815, 5.778131, 5.778115, 5.778116, 5.778116, 
    5.778112, 5.778121, 5.77811, 5.778109, 5.778113, 5.778086, 5.778093, 
    5.778085, 5.77809, 5.77822, 5.778214, 5.778217, 5.77821, 5.778215, 
    5.778194, 5.778188, 5.77816, 5.778172, 5.778153, 5.77817, 5.778167, 
    5.778152, 5.778169, 5.778132, 5.778157, 5.778111, 5.778136, 5.77811, 
    5.778115, 5.778107, 5.7781, 5.778091, 5.778075, 5.778079, 5.778065, 
    5.778204, 5.778195, 5.778196, 5.778188, 5.778181, 5.778167, 5.778145, 
    5.778153, 5.778138, 5.778135, 5.778158, 5.778144, 5.77819, 5.778183, 
    5.778187, 5.778203, 5.778151, 5.778178, 5.778129, 5.778143, 5.778101, 
    5.778122, 5.778081, 5.778063, 5.778047, 5.778027, 5.778191, 5.778197, 
    5.778186, 5.778172, 5.77816, 5.778142, 5.778141, 5.778137, 5.778129, 
    5.778122, 5.778136, 5.77812, 5.778181, 5.778149, 5.778199, 5.778184, 
    5.778173, 5.778178, 5.778154, 5.778149, 5.778126, 5.778138, 5.778068, 
    5.778099, 5.778013, 5.778037, 5.778199, 5.778191, 5.778164, 5.778177, 
    5.778141, 5.778132, 5.778125, 5.778116, 5.778115, 5.77811, 5.778118, 
    5.77811, 5.778142, 5.778128, 5.778168, 5.778158, 5.778162, 5.778167, 
    5.778152, 5.778136, 5.778136, 5.778131, 5.778116, 5.778141, 5.778063, 
    5.778111, 5.778183, 5.778168, 5.778166, 5.778172, 5.778133, 5.778147, 
    5.77811, 5.77812, 5.778103, 5.778111, 5.778112, 5.778123, 5.77813, 
    5.778146, 5.77816, 5.778171, 5.778168, 5.778156, 5.778135, 5.778115, 
    5.778119, 5.778104, 5.778144, 5.778127, 5.778133, 5.778117, 5.778153, 
    5.778122, 5.778162, 5.778158, 5.778147, 5.778126, 5.778121, 5.778116, 
    5.77812, 5.778134, 5.778137, 5.778148, 5.778151, 5.778159, 5.778165, 
    5.778159, 5.778153, 5.778134, 5.778118, 5.7781, 5.778095, 5.778074, 
    5.778091, 5.778063, 5.778087, 5.778046, 5.778121, 5.778088, 5.778147, 
    5.778141, 5.778129, 5.778103, 5.778117, 5.7781, 5.778137, 5.778156, 
    5.778161, 5.77817, 5.778161, 5.778162, 5.778152, 5.778155, 5.778134, 
    5.778145, 5.778112, 5.7781, 5.778067, 5.778046, 5.778025, 5.778015, 
    5.778012, 5.778011 ;

 SOIL1C_TO_SOIL2C =
  3.099197e-08, 3.112855e-08, 3.1102e-08, 3.121216e-08, 3.115106e-08, 
    3.122319e-08, 3.101967e-08, 3.113397e-08, 3.1061e-08, 3.100427e-08, 
    3.142594e-08, 3.121708e-08, 3.164294e-08, 3.150972e-08, 3.184439e-08, 
    3.162221e-08, 3.18892e-08, 3.183799e-08, 3.199213e-08, 3.194797e-08, 
    3.214512e-08, 3.201251e-08, 3.224732e-08, 3.211345e-08, 3.213439e-08, 
    3.200814e-08, 3.125912e-08, 3.139994e-08, 3.125077e-08, 3.127085e-08, 
    3.126184e-08, 3.115231e-08, 3.109712e-08, 3.098154e-08, 3.100252e-08, 
    3.108741e-08, 3.127988e-08, 3.121455e-08, 3.137922e-08, 3.13755e-08, 
    3.155882e-08, 3.147616e-08, 3.17843e-08, 3.169673e-08, 3.194982e-08, 
    3.188616e-08, 3.194683e-08, 3.192843e-08, 3.194706e-08, 3.185371e-08, 
    3.189371e-08, 3.181157e-08, 3.149164e-08, 3.158566e-08, 3.130525e-08, 
    3.113665e-08, 3.102468e-08, 3.094522e-08, 3.095645e-08, 3.097787e-08, 
    3.108791e-08, 3.119139e-08, 3.127024e-08, 3.132299e-08, 3.137496e-08, 
    3.153227e-08, 3.161555e-08, 3.180201e-08, 3.176837e-08, 3.182537e-08, 
    3.187983e-08, 3.197126e-08, 3.195622e-08, 3.19965e-08, 3.182387e-08, 
    3.19386e-08, 3.17492e-08, 3.1801e-08, 3.138907e-08, 3.123218e-08, 
    3.116547e-08, 3.110711e-08, 3.096509e-08, 3.106316e-08, 3.10245e-08, 
    3.111648e-08, 3.117493e-08, 3.114602e-08, 3.132443e-08, 3.125507e-08, 
    3.162048e-08, 3.146308e-08, 3.187348e-08, 3.177527e-08, 3.189702e-08, 
    3.18349e-08, 3.194134e-08, 3.184554e-08, 3.20115e-08, 3.204763e-08, 
    3.202294e-08, 3.21178e-08, 3.184023e-08, 3.194682e-08, 3.114521e-08, 
    3.114993e-08, 3.117189e-08, 3.107534e-08, 3.106943e-08, 3.098096e-08, 
    3.105968e-08, 3.109321e-08, 3.117832e-08, 3.122866e-08, 3.127651e-08, 
    3.138173e-08, 3.149924e-08, 3.166357e-08, 3.178164e-08, 3.186078e-08, 
    3.181225e-08, 3.18551e-08, 3.18072e-08, 3.178475e-08, 3.203409e-08, 
    3.189408e-08, 3.210416e-08, 3.209253e-08, 3.199746e-08, 3.209384e-08, 
    3.115323e-08, 3.112611e-08, 3.103191e-08, 3.110563e-08, 3.097133e-08, 
    3.10465e-08, 3.108972e-08, 3.125651e-08, 3.129317e-08, 3.132714e-08, 
    3.139426e-08, 3.148039e-08, 3.163149e-08, 3.176297e-08, 3.1883e-08, 
    3.187421e-08, 3.18773e-08, 3.190411e-08, 3.18377e-08, 3.191502e-08, 
    3.192799e-08, 3.189407e-08, 3.209098e-08, 3.203472e-08, 3.209228e-08, 
    3.205566e-08, 3.113493e-08, 3.118058e-08, 3.115591e-08, 3.120229e-08, 
    3.116961e-08, 3.131492e-08, 3.135849e-08, 3.156236e-08, 3.14787e-08, 
    3.161186e-08, 3.149222e-08, 3.151342e-08, 3.161619e-08, 3.149869e-08, 
    3.175572e-08, 3.158145e-08, 3.190516e-08, 3.173112e-08, 3.191606e-08, 
    3.188248e-08, 3.193808e-08, 3.198788e-08, 3.205053e-08, 3.216612e-08, 
    3.213936e-08, 3.223603e-08, 3.124863e-08, 3.130784e-08, 3.130263e-08, 
    3.13646e-08, 3.141042e-08, 3.150976e-08, 3.166907e-08, 3.160917e-08, 
    3.171916e-08, 3.174124e-08, 3.157414e-08, 3.167673e-08, 3.134747e-08, 
    3.140066e-08, 3.136899e-08, 3.12533e-08, 3.162296e-08, 3.143325e-08, 
    3.178359e-08, 3.168081e-08, 3.198078e-08, 3.183159e-08, 3.212462e-08, 
    3.224988e-08, 3.23678e-08, 3.250558e-08, 3.134016e-08, 3.129993e-08, 
    3.137197e-08, 3.147163e-08, 3.156412e-08, 3.168708e-08, 3.169966e-08, 
    3.172269e-08, 3.178236e-08, 3.183253e-08, 3.172997e-08, 3.18451e-08, 
    3.141299e-08, 3.163943e-08, 3.128471e-08, 3.139152e-08, 3.146576e-08, 
    3.14332e-08, 3.160232e-08, 3.164218e-08, 3.180416e-08, 3.172043e-08, 
    3.221896e-08, 3.199839e-08, 3.26105e-08, 3.243943e-08, 3.128587e-08, 
    3.134002e-08, 3.152849e-08, 3.143882e-08, 3.169529e-08, 3.175841e-08, 
    3.180974e-08, 3.187534e-08, 3.188243e-08, 3.19213e-08, 3.18576e-08, 
    3.191878e-08, 3.168734e-08, 3.179077e-08, 3.150695e-08, 3.157603e-08, 
    3.154425e-08, 3.150939e-08, 3.161697e-08, 3.173158e-08, 3.173404e-08, 
    3.177079e-08, 3.187433e-08, 3.169633e-08, 3.224742e-08, 3.190706e-08, 
    3.139907e-08, 3.150337e-08, 3.151828e-08, 3.147787e-08, 3.175209e-08, 
    3.165272e-08, 3.192035e-08, 3.184802e-08, 3.196653e-08, 3.190764e-08, 
    3.189898e-08, 3.182334e-08, 3.177625e-08, 3.165728e-08, 3.156049e-08, 
    3.148374e-08, 3.150158e-08, 3.158589e-08, 3.17386e-08, 3.188307e-08, 
    3.185142e-08, 3.195753e-08, 3.167669e-08, 3.179444e-08, 3.174893e-08, 
    3.186761e-08, 3.160757e-08, 3.182899e-08, 3.155098e-08, 3.157535e-08, 
    3.165075e-08, 3.180243e-08, 3.1836e-08, 3.187182e-08, 3.184972e-08, 
    3.174247e-08, 3.172491e-08, 3.164892e-08, 3.162794e-08, 3.157005e-08, 
    3.152211e-08, 3.156591e-08, 3.16119e-08, 3.174252e-08, 3.186024e-08, 
    3.198858e-08, 3.202e-08, 3.216995e-08, 3.204788e-08, 3.224931e-08, 
    3.207804e-08, 3.237454e-08, 3.184183e-08, 3.207301e-08, 3.165419e-08, 
    3.169931e-08, 3.178091e-08, 3.19681e-08, 3.186705e-08, 3.198523e-08, 
    3.172422e-08, 3.15888e-08, 3.155377e-08, 3.14884e-08, 3.155526e-08, 
    3.154982e-08, 3.16138e-08, 3.159325e-08, 3.174686e-08, 3.166435e-08, 
    3.189876e-08, 3.19843e-08, 3.22259e-08, 3.2374e-08, 3.252478e-08, 
    3.259135e-08, 3.261161e-08, 3.262008e-08 ;

 SOIL1C_TO_SOIL3C =
  3.675989e-10, 3.692194e-10, 3.689044e-10, 3.702115e-10, 3.694864e-10, 
    3.703423e-10, 3.679275e-10, 3.692837e-10, 3.684179e-10, 3.677448e-10, 
    3.727481e-10, 3.702698e-10, 3.753229e-10, 3.737421e-10, 3.777133e-10, 
    3.750769e-10, 3.782449e-10, 3.776373e-10, 3.794663e-10, 3.789423e-10, 
    3.812817e-10, 3.797082e-10, 3.824945e-10, 3.80906e-10, 3.811544e-10, 
    3.796563e-10, 3.707686e-10, 3.724395e-10, 3.706696e-10, 3.709079e-10, 
    3.708009e-10, 3.695014e-10, 3.688465e-10, 3.674751e-10, 3.67724e-10, 
    3.687313e-10, 3.71015e-10, 3.702398e-10, 3.721936e-10, 3.721495e-10, 
    3.743247e-10, 3.73344e-10, 3.770003e-10, 3.759611e-10, 3.789642e-10, 
    3.782089e-10, 3.789287e-10, 3.787105e-10, 3.789316e-10, 3.778239e-10, 
    3.782984e-10, 3.773238e-10, 3.735276e-10, 3.746432e-10, 3.71316e-10, 
    3.693155e-10, 3.679869e-10, 3.670441e-10, 3.671774e-10, 3.674315e-10, 
    3.687372e-10, 3.69965e-10, 3.709006e-10, 3.715265e-10, 3.721432e-10, 
    3.740097e-10, 3.749979e-10, 3.772104e-10, 3.768112e-10, 3.774875e-10, 
    3.781338e-10, 3.792188e-10, 3.790402e-10, 3.795182e-10, 3.774697e-10, 
    3.788311e-10, 3.765837e-10, 3.771984e-10, 3.723106e-10, 3.70449e-10, 
    3.696575e-10, 3.689649e-10, 3.672799e-10, 3.684435e-10, 3.679848e-10, 
    3.690762e-10, 3.697697e-10, 3.694267e-10, 3.715436e-10, 3.707206e-10, 
    3.750564e-10, 3.731888e-10, 3.780584e-10, 3.768931e-10, 3.783378e-10, 
    3.776006e-10, 3.788637e-10, 3.777269e-10, 3.796961e-10, 3.801249e-10, 
    3.798319e-10, 3.809575e-10, 3.776639e-10, 3.789287e-10, 3.694171e-10, 
    3.69473e-10, 3.697336e-10, 3.68588e-10, 3.68518e-10, 3.674682e-10, 
    3.684023e-10, 3.688001e-10, 3.698099e-10, 3.704072e-10, 3.70975e-10, 
    3.722234e-10, 3.736178e-10, 3.755677e-10, 3.769687e-10, 3.779077e-10, 
    3.773319e-10, 3.778403e-10, 3.77272e-10, 3.770056e-10, 3.799642e-10, 
    3.783029e-10, 3.807956e-10, 3.806577e-10, 3.795295e-10, 3.806733e-10, 
    3.695123e-10, 3.691904e-10, 3.680728e-10, 3.689474e-10, 3.673539e-10, 
    3.682459e-10, 3.687587e-10, 3.707377e-10, 3.711726e-10, 3.715758e-10, 
    3.723722e-10, 3.733941e-10, 3.751871e-10, 3.767471e-10, 3.781714e-10, 
    3.78067e-10, 3.781038e-10, 3.78422e-10, 3.776338e-10, 3.785513e-10, 
    3.787053e-10, 3.783027e-10, 3.806392e-10, 3.799717e-10, 3.806548e-10, 
    3.802202e-10, 3.692951e-10, 3.698367e-10, 3.69544e-10, 3.700944e-10, 
    3.697066e-10, 3.714307e-10, 3.719477e-10, 3.743668e-10, 3.73374e-10, 
    3.749541e-10, 3.735346e-10, 3.737861e-10, 3.750055e-10, 3.736113e-10, 
    3.766611e-10, 3.745933e-10, 3.784343e-10, 3.763692e-10, 3.785637e-10, 
    3.781652e-10, 3.78825e-10, 3.794159e-10, 3.801593e-10, 3.81531e-10, 
    3.812133e-10, 3.823605e-10, 3.706442e-10, 3.713467e-10, 3.712849e-10, 
    3.720202e-10, 3.725639e-10, 3.737426e-10, 3.75633e-10, 3.749221e-10, 
    3.762272e-10, 3.764893e-10, 3.745065e-10, 3.757238e-10, 3.718169e-10, 
    3.724481e-10, 3.720723e-10, 3.706996e-10, 3.750859e-10, 3.728347e-10, 
    3.769918e-10, 3.757722e-10, 3.793316e-10, 3.775614e-10, 3.810385e-10, 
    3.825249e-10, 3.839241e-10, 3.855591e-10, 3.717302e-10, 3.712528e-10, 
    3.721076e-10, 3.732902e-10, 3.743876e-10, 3.758466e-10, 3.759959e-10, 
    3.762692e-10, 3.769772e-10, 3.775725e-10, 3.763556e-10, 3.777217e-10, 
    3.725943e-10, 3.752813e-10, 3.710723e-10, 3.723396e-10, 3.732205e-10, 
    3.728342e-10, 3.748409e-10, 3.753139e-10, 3.772359e-10, 3.762423e-10, 
    3.82158e-10, 3.795406e-10, 3.868041e-10, 3.847741e-10, 3.710861e-10, 
    3.717286e-10, 3.739649e-10, 3.729008e-10, 3.75944e-10, 3.766931e-10, 
    3.773021e-10, 3.780805e-10, 3.781646e-10, 3.786258e-10, 3.7787e-10, 
    3.78596e-10, 3.758497e-10, 3.770769e-10, 3.737093e-10, 3.745289e-10, 
    3.741519e-10, 3.737383e-10, 3.750148e-10, 3.763747e-10, 3.764039e-10, 
    3.768399e-10, 3.780685e-10, 3.759563e-10, 3.824956e-10, 3.784569e-10, 
    3.724293e-10, 3.736668e-10, 3.738437e-10, 3.733643e-10, 3.76618e-10, 
    3.75439e-10, 3.786146e-10, 3.777563e-10, 3.791626e-10, 3.784638e-10, 
    3.78361e-10, 3.774635e-10, 3.769047e-10, 3.754931e-10, 3.743445e-10, 
    3.734338e-10, 3.736456e-10, 3.74646e-10, 3.764579e-10, 3.781722e-10, 
    3.777967e-10, 3.790557e-10, 3.757233e-10, 3.771206e-10, 3.765805e-10, 
    3.779888e-10, 3.749032e-10, 3.775305e-10, 3.742317e-10, 3.745209e-10, 
    3.754156e-10, 3.772153e-10, 3.776136e-10, 3.780387e-10, 3.777764e-10, 
    3.765039e-10, 3.762955e-10, 3.753939e-10, 3.751449e-10, 3.744579e-10, 
    3.738892e-10, 3.744088e-10, 3.749545e-10, 3.765045e-10, 3.779013e-10, 
    3.794243e-10, 3.79797e-10, 3.815764e-10, 3.801278e-10, 3.825181e-10, 
    3.804857e-10, 3.840041e-10, 3.776829e-10, 3.804261e-10, 3.754563e-10, 
    3.759917e-10, 3.769601e-10, 3.791812e-10, 3.779821e-10, 3.793845e-10, 
    3.762873e-10, 3.746805e-10, 3.742648e-10, 3.734892e-10, 3.742825e-10, 
    3.74218e-10, 3.749772e-10, 3.747332e-10, 3.76556e-10, 3.755769e-10, 
    3.783584e-10, 3.793734e-10, 3.822403e-10, 3.839978e-10, 3.85787e-10, 
    3.865769e-10, 3.868173e-10, 3.869178e-10 ;

 SOIL1C_vr =
  19.98109, 19.98104, 19.98105, 19.98101, 19.98103, 19.981, 19.98108, 
    19.98104, 19.98107, 19.98109, 19.98093, 19.98101, 19.98085, 19.9809, 
    19.98077, 19.98085, 19.98075, 19.98077, 19.98071, 19.98073, 19.98066, 
    19.98071, 19.98062, 19.98067, 19.98066, 19.98071, 19.98099, 19.98094, 
    19.981, 19.98099, 19.98099, 19.98103, 19.98105, 19.9811, 19.98109, 
    19.98106, 19.98098, 19.98101, 19.98095, 19.98095, 19.98088, 19.98091, 
    19.98079, 19.98083, 19.98073, 19.98075, 19.98073, 19.98074, 19.98073, 
    19.98077, 19.98075, 19.98078, 19.9809, 19.98087, 19.98097, 19.98104, 
    19.98108, 19.98111, 19.98111, 19.9811, 19.98106, 19.98102, 19.98099, 
    19.98097, 19.98095, 19.98089, 19.98086, 19.98079, 19.9808, 19.98078, 
    19.98076, 19.98072, 19.98073, 19.98071, 19.98078, 19.98074, 19.98081, 
    19.98079, 19.98094, 19.981, 19.98103, 19.98105, 19.9811, 19.98107, 
    19.98108, 19.98104, 19.98102, 19.98103, 19.98097, 19.98099, 19.98086, 
    19.98092, 19.98076, 19.9808, 19.98075, 19.98077, 19.98073, 19.98077, 
    19.98071, 19.98069, 19.9807, 19.98067, 19.98077, 19.98073, 19.98104, 
    19.98103, 19.98102, 19.98106, 19.98106, 19.9811, 19.98107, 19.98105, 
    19.98102, 19.981, 19.98099, 19.98095, 19.9809, 19.98084, 19.98079, 
    19.98076, 19.98078, 19.98077, 19.98079, 19.98079, 19.9807, 19.98075, 
    19.98067, 19.98068, 19.98071, 19.98068, 19.98103, 19.98104, 19.98108, 
    19.98105, 19.9811, 19.98107, 19.98106, 19.98099, 19.98098, 19.98097, 
    19.98094, 19.98091, 19.98085, 19.9808, 19.98076, 19.98076, 19.98076, 
    19.98075, 19.98077, 19.98075, 19.98074, 19.98075, 19.98068, 19.9807, 
    19.98068, 19.98069, 19.98104, 19.98102, 19.98103, 19.98101, 19.98103, 
    19.98097, 19.98095, 19.98088, 19.98091, 19.98086, 19.9809, 19.9809, 
    19.98086, 19.9809, 19.9808, 19.98087, 19.98075, 19.98081, 19.98074, 
    19.98076, 19.98074, 19.98072, 19.98069, 19.98065, 19.98066, 19.98062, 
    19.981, 19.98097, 19.98097, 19.98095, 19.98093, 19.9809, 19.98084, 
    19.98086, 19.98082, 19.98081, 19.98087, 19.98083, 19.98096, 19.98094, 
    19.98095, 19.98099, 19.98085, 19.98093, 19.98079, 19.98083, 19.98072, 
    19.98078, 19.98067, 19.98062, 19.98058, 19.98052, 19.98096, 19.98098, 
    19.98095, 19.98091, 19.98088, 19.98083, 19.98083, 19.98082, 19.98079, 
    19.98078, 19.98081, 19.98077, 19.98093, 19.98085, 19.98098, 19.98094, 
    19.98091, 19.98093, 19.98086, 19.98085, 19.98079, 19.98082, 19.98063, 
    19.98071, 19.98048, 19.98055, 19.98098, 19.98096, 19.98089, 19.98092, 
    19.98083, 19.9808, 19.98078, 19.98076, 19.98076, 19.98074, 19.98077, 
    19.98074, 19.98083, 19.98079, 19.9809, 19.98087, 19.98088, 19.9809, 
    19.98086, 19.98081, 19.98081, 19.9808, 19.98076, 19.98083, 19.98062, 
    19.98075, 19.98094, 19.9809, 19.98089, 19.98091, 19.98081, 19.98084, 
    19.98074, 19.98077, 19.98072, 19.98075, 19.98075, 19.98078, 19.9808, 
    19.98084, 19.98088, 19.98091, 19.9809, 19.98087, 19.98081, 19.98076, 
    19.98077, 19.98073, 19.98083, 19.98079, 19.98081, 19.98076, 19.98086, 
    19.98078, 19.98088, 19.98087, 19.98084, 19.98079, 19.98077, 19.98076, 
    19.98077, 19.98081, 19.98082, 19.98084, 19.98085, 19.98088, 19.98089, 
    19.98088, 19.98086, 19.98081, 19.98076, 19.98072, 19.98071, 19.98065, 
    19.98069, 19.98062, 19.98068, 19.98057, 19.98077, 19.98068, 19.98084, 
    19.98083, 19.98079, 19.98072, 19.98076, 19.98072, 19.98082, 19.98087, 
    19.98088, 19.98091, 19.98088, 19.98088, 19.98086, 19.98087, 19.98081, 
    19.98084, 19.98075, 19.98072, 19.98063, 19.98057, 19.98052, 19.98049, 
    19.98048, 19.98048,
  19.98328, 19.98321, 19.98323, 19.98318, 19.9832, 19.98317, 19.98326, 
    19.98321, 19.98325, 19.98327, 19.98308, 19.98317, 19.98298, 19.98304, 
    19.98288, 19.98298, 19.98286, 19.98288, 19.98281, 19.98283, 19.98274, 
    19.9828, 19.98269, 19.98276, 19.98275, 19.98281, 19.98315, 19.98309, 
    19.98316, 19.98315, 19.98315, 19.9832, 19.98323, 19.98328, 19.98327, 
    19.98323, 19.98314, 19.98317, 19.9831, 19.9831, 19.98301, 19.98305, 
    19.98291, 19.98295, 19.98283, 19.98286, 19.98283, 19.98284, 19.98283, 
    19.98288, 19.98286, 19.98289, 19.98304, 19.983, 19.98313, 19.98321, 
    19.98326, 19.9833, 19.98329, 19.98328, 19.98323, 19.98318, 19.98315, 
    19.98312, 19.9831, 19.98303, 19.98299, 19.9829, 19.98292, 19.98289, 
    19.98286, 19.98282, 19.98283, 19.98281, 19.98289, 19.98284, 19.98293, 
    19.9829, 19.98309, 19.98317, 19.9832, 19.98322, 19.98329, 19.98324, 
    19.98326, 19.98322, 19.98319, 19.98321, 19.98312, 19.98315, 19.98298, 
    19.98306, 19.98287, 19.98291, 19.98286, 19.98289, 19.98284, 19.98288, 
    19.9828, 19.98279, 19.9828, 19.98275, 19.98288, 19.98283, 19.98321, 
    19.9832, 19.98319, 19.98324, 19.98324, 19.98328, 19.98325, 19.98323, 
    19.98319, 19.98317, 19.98314, 19.9831, 19.98304, 19.98297, 19.98291, 
    19.98287, 19.98289, 19.98288, 19.9829, 19.98291, 19.98279, 19.98286, 
    19.98276, 19.98277, 19.98281, 19.98277, 19.9832, 19.98322, 19.98326, 
    19.98322, 19.98329, 19.98325, 19.98323, 19.98315, 19.98314, 19.98312, 
    19.98309, 19.98305, 19.98298, 19.98292, 19.98286, 19.98287, 19.98286, 
    19.98285, 19.98288, 19.98285, 19.98284, 19.98286, 19.98277, 19.98279, 
    19.98277, 19.98278, 19.98321, 19.98319, 19.9832, 19.98318, 19.98319, 
    19.98313, 19.98311, 19.98301, 19.98305, 19.98299, 19.98304, 19.98303, 
    19.98299, 19.98304, 19.98292, 19.983, 19.98285, 19.98293, 19.98285, 
    19.98286, 19.98284, 19.98281, 19.98278, 19.98273, 19.98274, 19.9827, 
    19.98316, 19.98313, 19.98313, 19.9831, 19.98308, 19.98304, 19.98296, 
    19.98299, 19.98294, 19.98293, 19.98301, 19.98296, 19.98311, 19.98309, 
    19.9831, 19.98316, 19.98298, 19.98307, 19.98291, 19.98296, 19.98282, 
    19.98289, 19.98275, 19.98269, 19.98264, 19.98257, 19.98312, 19.98313, 
    19.9831, 19.98305, 19.98301, 19.98295, 19.98295, 19.98294, 19.98291, 
    19.98289, 19.98293, 19.98288, 19.98308, 19.98298, 19.98314, 19.98309, 
    19.98306, 19.98307, 19.98299, 19.98298, 19.9829, 19.98294, 19.98271, 
    19.98281, 19.98252, 19.9826, 19.98314, 19.98312, 19.98303, 19.98307, 
    19.98295, 19.98292, 19.9829, 19.98287, 19.98286, 19.98285, 19.98287, 
    19.98285, 19.98295, 19.98291, 19.98304, 19.98301, 19.98302, 19.98304, 
    19.98299, 19.98293, 19.98293, 19.98291, 19.98287, 19.98295, 19.98269, 
    19.98285, 19.98309, 19.98304, 19.98303, 19.98305, 19.98292, 19.98297, 
    19.98285, 19.98288, 19.98282, 19.98285, 19.98285, 19.98289, 19.98291, 
    19.98297, 19.98301, 19.98305, 19.98304, 19.983, 19.98293, 19.98286, 
    19.98288, 19.98283, 19.98296, 19.9829, 19.98293, 19.98287, 19.98299, 
    19.98289, 19.98302, 19.98301, 19.98297, 19.9829, 19.98288, 19.98287, 
    19.98288, 19.98293, 19.98294, 19.98297, 19.98298, 19.98301, 19.98303, 
    19.98301, 19.98299, 19.98293, 19.98287, 19.98281, 19.9828, 19.98273, 
    19.98279, 19.98269, 19.98277, 19.98264, 19.98288, 19.98277, 19.98297, 
    19.98295, 19.98291, 19.98282, 19.98287, 19.98281, 19.98294, 19.983, 
    19.98302, 19.98305, 19.98302, 19.98302, 19.98299, 19.983, 19.98293, 
    19.98296, 19.98285, 19.98281, 19.9827, 19.98264, 19.98256, 19.98253, 
    19.98252, 19.98252,
  19.98426, 19.98419, 19.9842, 19.98414, 19.98418, 19.98414, 19.98424, 
    19.98418, 19.98422, 19.98425, 19.98404, 19.98414, 19.98392, 19.98399, 
    19.98382, 19.98393, 19.9838, 19.98383, 19.98375, 19.98377, 19.98367, 
    19.98374, 19.98362, 19.98368, 19.98368, 19.98374, 19.98412, 19.98405, 
    19.98413, 19.98411, 19.98412, 19.98417, 19.9842, 19.98426, 19.98425, 
    19.98421, 19.98411, 19.98414, 19.98406, 19.98406, 19.98397, 19.98401, 
    19.98385, 19.9839, 19.98377, 19.9838, 19.98377, 19.98378, 19.98377, 
    19.98382, 19.9838, 19.98384, 19.984, 19.98395, 19.9841, 19.98418, 
    19.98424, 19.98428, 19.98428, 19.98426, 19.98421, 19.98416, 19.98412, 
    19.98409, 19.98406, 19.98398, 19.98394, 19.98384, 19.98386, 19.98383, 
    19.9838, 19.98376, 19.98376, 19.98375, 19.98383, 19.98377, 19.98387, 
    19.98384, 19.98405, 19.98413, 19.98417, 19.9842, 19.98427, 19.98422, 
    19.98424, 19.98419, 19.98416, 19.98418, 19.98409, 19.98412, 19.98394, 
    19.98402, 19.98381, 19.98386, 19.9838, 19.98383, 19.98377, 19.98382, 
    19.98374, 19.98372, 19.98373, 19.98368, 19.98382, 19.98377, 19.98418, 
    19.98418, 19.98417, 19.98421, 19.98422, 19.98426, 19.98422, 19.98421, 
    19.98416, 19.98414, 19.98411, 19.98406, 19.984, 19.98391, 19.98385, 
    19.98381, 19.98384, 19.98382, 19.98384, 19.98385, 19.98372, 19.9838, 
    19.98369, 19.9837, 19.98374, 19.9837, 19.98417, 19.98419, 19.98424, 
    19.9842, 19.98427, 19.98423, 19.98421, 19.98412, 19.9841, 19.98409, 
    19.98405, 19.98401, 19.98393, 19.98386, 19.9838, 19.98381, 19.9838, 
    19.98379, 19.98383, 19.98379, 19.98378, 19.9838, 19.9837, 19.98372, 
    19.9837, 19.98372, 19.98418, 19.98416, 19.98417, 19.98415, 19.98417, 
    19.98409, 19.98407, 19.98396, 19.98401, 19.98394, 19.984, 19.98399, 
    19.98394, 19.984, 19.98387, 19.98396, 19.98379, 19.98388, 19.98379, 
    19.9838, 19.98377, 19.98375, 19.98372, 19.98366, 19.98367, 19.98362, 
    19.98413, 19.9841, 19.9841, 19.98407, 19.98404, 19.98399, 19.98391, 
    19.98394, 19.98389, 19.98388, 19.98396, 19.98391, 19.98408, 19.98405, 
    19.98406, 19.98412, 19.98393, 19.98403, 19.98385, 19.98391, 19.98375, 
    19.98383, 19.98368, 19.98362, 19.98356, 19.98349, 19.98408, 19.9841, 
    19.98406, 19.98401, 19.98396, 19.9839, 19.9839, 19.98388, 19.98385, 
    19.98383, 19.98388, 19.98382, 19.98404, 19.98393, 19.98411, 19.98405, 
    19.98401, 19.98403, 19.98395, 19.98392, 19.98384, 19.98388, 19.98363, 
    19.98374, 19.98343, 19.98352, 19.98411, 19.98408, 19.98398, 19.98403, 
    19.9839, 19.98387, 19.98384, 19.98381, 19.9838, 19.98378, 19.98382, 
    19.98378, 19.9839, 19.98385, 19.98399, 19.98396, 19.98397, 19.98399, 
    19.98394, 19.98388, 19.98388, 19.98386, 19.98381, 19.9839, 19.98362, 
    19.98379, 19.98405, 19.984, 19.98399, 19.98401, 19.98387, 19.98392, 
    19.98378, 19.98382, 19.98376, 19.98379, 19.9838, 19.98383, 19.98386, 
    19.98392, 19.98397, 19.984, 19.984, 19.98395, 19.98388, 19.9838, 
    19.98382, 19.98376, 19.98391, 19.98385, 19.98387, 19.98381, 19.98394, 
    19.98383, 19.98397, 19.98396, 19.98392, 19.98384, 19.98383, 19.98381, 
    19.98382, 19.98387, 19.98388, 19.98392, 19.98393, 19.98396, 19.98399, 
    19.98396, 19.98394, 19.98387, 19.98381, 19.98375, 19.98373, 19.98366, 
    19.98372, 19.98362, 19.9837, 19.98355, 19.98382, 19.98371, 19.98392, 
    19.9839, 19.98385, 19.98376, 19.98381, 19.98375, 19.98388, 19.98395, 
    19.98397, 19.984, 19.98397, 19.98397, 19.98394, 19.98395, 19.98387, 
    19.98391, 19.9838, 19.98375, 19.98363, 19.98355, 19.98348, 19.98344, 
    19.98343, 19.98343,
  19.98501, 19.98494, 19.98495, 19.98489, 19.98492, 19.98489, 19.98499, 
    19.98493, 19.98497, 19.985, 19.98478, 19.98489, 19.98467, 19.98474, 
    19.98456, 19.98468, 19.98454, 19.98457, 19.98449, 19.98451, 19.98441, 
    19.98448, 19.98435, 19.98442, 19.98441, 19.98448, 19.98487, 19.98479, 
    19.98487, 19.98486, 19.98487, 19.98492, 19.98495, 19.98501, 19.985, 
    19.98496, 19.98486, 19.98489, 19.9848, 19.98481, 19.98471, 19.98475, 
    19.98459, 19.98464, 19.98451, 19.98454, 19.98451, 19.98452, 19.98451, 
    19.98456, 19.98454, 19.98458, 19.98475, 19.9847, 19.98484, 19.98493, 
    19.98499, 19.98503, 19.98503, 19.98501, 19.98496, 19.9849, 19.98486, 
    19.98483, 19.98481, 19.98473, 19.98468, 19.98458, 19.9846, 19.98457, 
    19.98454, 19.9845, 19.9845, 19.98448, 19.98457, 19.98451, 19.98461, 
    19.98458, 19.9848, 19.98488, 19.98492, 19.98495, 19.98502, 19.98497, 
    19.98499, 19.98494, 19.98491, 19.98493, 19.98483, 19.98487, 19.98468, 
    19.98476, 19.98455, 19.9846, 19.98454, 19.98457, 19.98451, 19.98456, 
    19.98448, 19.98446, 19.98447, 19.98442, 19.98457, 19.98451, 19.98493, 
    19.98492, 19.98491, 19.98496, 19.98497, 19.98501, 19.98497, 19.98495, 
    19.98491, 19.98488, 19.98486, 19.9848, 19.98474, 19.98466, 19.9846, 
    19.98455, 19.98458, 19.98456, 19.98458, 19.98459, 19.98446, 19.98454, 
    19.98443, 19.98443, 19.98448, 19.98443, 19.98492, 19.98494, 19.98499, 
    19.98495, 19.98502, 19.98498, 19.98496, 19.98487, 19.98485, 19.98483, 
    19.9848, 19.98475, 19.98467, 19.98461, 19.98454, 19.98455, 19.98454, 
    19.98453, 19.98457, 19.98453, 19.98452, 19.98454, 19.98443, 19.98446, 
    19.98443, 19.98445, 19.98493, 19.98491, 19.98492, 19.9849, 19.98491, 
    19.98484, 19.98482, 19.98471, 19.98475, 19.98468, 19.98475, 19.98474, 
    19.98468, 19.98474, 19.98461, 19.9847, 19.98453, 19.98462, 19.98453, 
    19.98454, 19.98451, 19.98449, 19.98446, 19.9844, 19.98441, 19.98436, 
    19.98487, 19.98484, 19.98484, 19.98481, 19.98479, 19.98474, 19.98465, 
    19.98469, 19.98463, 19.98462, 19.9847, 19.98465, 19.98482, 19.98479, 
    19.98481, 19.98487, 19.98468, 19.98478, 19.98459, 19.98465, 19.98449, 
    19.98457, 19.98442, 19.98435, 19.98429, 19.98422, 19.98483, 19.98485, 
    19.98481, 19.98476, 19.98471, 19.98464, 19.98464, 19.98463, 19.98459, 
    19.98457, 19.98462, 19.98456, 19.98479, 19.98467, 19.98485, 19.9848, 
    19.98476, 19.98478, 19.98469, 19.98467, 19.98458, 19.98463, 19.98437, 
    19.98448, 19.98417, 19.98425, 19.98485, 19.98483, 19.98473, 19.98477, 
    19.98464, 19.98461, 19.98458, 19.98455, 19.98454, 19.98452, 19.98456, 
    19.98452, 19.98464, 19.98459, 19.98474, 19.9847, 19.98472, 19.98474, 
    19.98468, 19.98462, 19.98462, 19.9846, 19.98455, 19.98464, 19.98435, 
    19.98453, 19.98479, 19.98474, 19.98473, 19.98475, 19.98461, 19.98466, 
    19.98452, 19.98456, 19.9845, 19.98453, 19.98454, 19.98457, 19.9846, 
    19.98466, 19.98471, 19.98475, 19.98474, 19.9847, 19.98462, 19.98454, 
    19.98456, 19.9845, 19.98465, 19.98459, 19.98461, 19.98455, 19.98469, 
    19.98457, 19.98472, 19.9847, 19.98466, 19.98458, 19.98457, 19.98455, 
    19.98456, 19.98462, 19.98462, 19.98466, 19.98468, 19.9847, 19.98473, 
    19.98471, 19.98468, 19.98462, 19.98455, 19.98449, 19.98447, 19.98439, 
    19.98446, 19.98435, 19.98444, 19.98429, 19.98456, 19.98444, 19.98466, 
    19.98464, 19.9846, 19.9845, 19.98455, 19.98449, 19.98462, 19.9847, 
    19.98471, 19.98475, 19.98471, 19.98472, 19.98468, 19.98469, 19.98461, 
    19.98466, 19.98454, 19.98449, 19.98436, 19.98429, 19.98421, 19.98417, 
    19.98416, 19.98416,
  19.98609, 19.98602, 19.98603, 19.98598, 19.98601, 19.98598, 19.98607, 
    19.98602, 19.98605, 19.98608, 19.98588, 19.98598, 19.98577, 19.98584, 
    19.98568, 19.98579, 19.98566, 19.98568, 19.98561, 19.98563, 19.98554, 
    19.9856, 19.98549, 19.98555, 19.98554, 19.9856, 19.98596, 19.98589, 
    19.98596, 19.98595, 19.98596, 19.98601, 19.98603, 19.98609, 19.98608, 
    19.98604, 19.98595, 19.98598, 19.9859, 19.9859, 19.98582, 19.98586, 
    19.98571, 19.98575, 19.98563, 19.98566, 19.98563, 19.98564, 19.98563, 
    19.98568, 19.98566, 19.98569, 19.98585, 19.9858, 19.98594, 19.98602, 
    19.98607, 19.98611, 19.9861, 19.98609, 19.98604, 19.98599, 19.98595, 
    19.98593, 19.9859, 19.98583, 19.98579, 19.9857, 19.98572, 19.98569, 
    19.98566, 19.98562, 19.98563, 19.98561, 19.98569, 19.98564, 19.98573, 
    19.9857, 19.9859, 19.98597, 19.986, 19.98603, 19.9861, 19.98605, 
    19.98607, 19.98603, 19.986, 19.98601, 19.98593, 19.98596, 19.98579, 
    19.98586, 19.98567, 19.98571, 19.98565, 19.98568, 19.98563, 19.98568, 
    19.9856, 19.98558, 19.98559, 19.98555, 19.98568, 19.98563, 19.98601, 
    19.98601, 19.986, 19.98605, 19.98605, 19.98609, 19.98605, 19.98604, 
    19.986, 19.98597, 19.98595, 19.9859, 19.98584, 19.98577, 19.98571, 
    19.98567, 19.98569, 19.98567, 19.9857, 19.98571, 19.98559, 19.98566, 
    19.98556, 19.98556, 19.98561, 19.98556, 19.98601, 19.98602, 19.98607, 
    19.98603, 19.9861, 19.98606, 19.98604, 19.98596, 19.98594, 19.98593, 
    19.98589, 19.98585, 19.98578, 19.98572, 19.98566, 19.98567, 19.98566, 
    19.98565, 19.98568, 19.98565, 19.98564, 19.98566, 19.98556, 19.98559, 
    19.98556, 19.98558, 19.98602, 19.986, 19.98601, 19.98598, 19.986, 
    19.98593, 19.98591, 19.98581, 19.98585, 19.98579, 19.98585, 19.98584, 
    19.98579, 19.98584, 19.98572, 19.98581, 19.98565, 19.98573, 19.98565, 
    19.98566, 19.98564, 19.98561, 19.98558, 19.98553, 19.98554, 19.98549, 
    19.98596, 19.98594, 19.98594, 19.98591, 19.98589, 19.98584, 19.98576, 
    19.98579, 19.98574, 19.98573, 19.98581, 19.98576, 19.98592, 19.98589, 
    19.98591, 19.98596, 19.98578, 19.98588, 19.98571, 19.98576, 19.98561, 
    19.98569, 19.98555, 19.98549, 19.98543, 19.98536, 19.98592, 19.98594, 
    19.9859, 19.98586, 19.98581, 19.98575, 19.98575, 19.98574, 19.98571, 
    19.98569, 19.98573, 19.98568, 19.98589, 19.98578, 19.98595, 19.9859, 
    19.98586, 19.98588, 19.9858, 19.98578, 19.9857, 19.98574, 19.9855, 
    19.98561, 19.98531, 19.9854, 19.98594, 19.98592, 19.98583, 19.98587, 
    19.98575, 19.98572, 19.9857, 19.98566, 19.98566, 19.98564, 19.98567, 
    19.98564, 19.98575, 19.9857, 19.98584, 19.98581, 19.98582, 19.98584, 
    19.98579, 19.98573, 19.98573, 19.98571, 19.98567, 19.98575, 19.98549, 
    19.98565, 19.98589, 19.98584, 19.98583, 19.98586, 19.98572, 19.98577, 
    19.98564, 19.98568, 19.98562, 19.98565, 19.98565, 19.98569, 19.98571, 
    19.98577, 19.98582, 19.98585, 19.98584, 19.9858, 19.98573, 19.98566, 
    19.98568, 19.98563, 19.98576, 19.9857, 19.98573, 19.98567, 19.98579, 
    19.98569, 19.98582, 19.98581, 19.98577, 19.9857, 19.98568, 19.98567, 
    19.98568, 19.98573, 19.98574, 19.98577, 19.98578, 19.98581, 19.98583, 
    19.98581, 19.98579, 19.98573, 19.98567, 19.98561, 19.9856, 19.98553, 
    19.98558, 19.98549, 19.98557, 19.98543, 19.98568, 19.98557, 19.98577, 
    19.98575, 19.98571, 19.98562, 19.98567, 19.98561, 19.98574, 19.9858, 
    19.98582, 19.98585, 19.98582, 19.98582, 19.98579, 19.9858, 19.98573, 
    19.98577, 19.98565, 19.98561, 19.9855, 19.98543, 19.98536, 19.98532, 
    19.98531, 19.98531,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.72228, 0.7222776, 0.7222781, 0.7222761, 0.7222772, 0.7222759, 0.7222795, 
    0.7222775, 0.7222788, 0.7222798, 0.7222724, 0.722276, 0.7222686, 
    0.7222709, 0.722265, 0.7222689, 0.7222642, 0.7222651, 0.7222624, 
    0.7222632, 0.7222598, 0.7222621, 0.722258, 0.7222603, 0.7222599, 
    0.7222621, 0.7222753, 0.7222728, 0.7222754, 0.7222751, 0.7222753, 
    0.7222772, 0.7222781, 0.7222801, 0.7222798, 0.7222783, 0.722275, 
    0.7222761, 0.7222732, 0.7222732, 0.72227, 0.7222715, 0.7222661, 
    0.7222676, 0.7222632, 0.7222643, 0.7222632, 0.7222635, 0.7222632, 
    0.7222648, 0.7222642, 0.7222656, 0.7222712, 0.7222695, 0.7222745, 
    0.7222775, 0.7222794, 0.7222808, 0.7222806, 0.7222803, 0.7222783, 
    0.7222765, 0.7222751, 0.7222742, 0.7222733, 0.7222705, 0.7222691, 
    0.7222658, 0.7222664, 0.7222654, 0.7222644, 0.7222628, 0.722263, 
    0.7222623, 0.7222654, 0.7222633, 0.7222667, 0.7222658, 0.722273, 
    0.7222758, 0.7222769, 0.7222779, 0.7222804, 0.7222787, 0.7222794, 
    0.7222778, 0.7222767, 0.7222773, 0.7222741, 0.7222754, 0.7222689, 
    0.7222717, 0.7222645, 0.7222663, 0.7222641, 0.7222652, 0.7222633, 
    0.722265, 0.7222621, 0.7222614, 0.7222619, 0.7222602, 0.7222651, 
    0.7222632, 0.7222773, 0.7222772, 0.7222768, 0.7222785, 0.7222787, 
    0.7222802, 0.7222788, 0.7222782, 0.7222767, 0.7222759, 0.722275, 
    0.7222732, 0.7222711, 0.7222682, 0.7222661, 0.7222647, 0.7222656, 
    0.7222648, 0.7222657, 0.7222661, 0.7222617, 0.7222642, 0.7222605, 
    0.7222607, 0.7222623, 0.7222607, 0.7222772, 0.7222776, 0.7222793, 
    0.722278, 0.7222803, 0.722279, 0.7222783, 0.7222753, 0.7222747, 
    0.7222741, 0.7222729, 0.7222714, 0.7222688, 0.7222664, 0.7222643, 
    0.7222645, 0.7222645, 0.722264, 0.7222651, 0.7222638, 0.7222636, 
    0.7222642, 0.7222607, 0.7222617, 0.7222607, 0.7222613, 0.7222775, 
    0.7222767, 0.7222771, 0.7222763, 0.7222769, 0.7222743, 0.7222735, 
    0.72227, 0.7222714, 0.7222691, 0.7222712, 0.7222708, 0.722269, 0.7222711, 
    0.7222666, 0.7222697, 0.7222639, 0.722267, 0.7222638, 0.7222643, 
    0.7222634, 0.7222625, 0.7222614, 0.7222593, 0.7222598, 0.7222582, 
    0.7222755, 0.7222744, 0.7222745, 0.7222735, 0.7222726, 0.7222709, 
    0.7222681, 0.7222692, 0.7222672, 0.7222669, 0.7222698, 0.722268, 
    0.7222738, 0.7222728, 0.7222733, 0.7222754, 0.7222689, 0.7222722, 
    0.7222661, 0.7222679, 0.7222626, 0.7222652, 0.7222601, 0.7222579, 
    0.7222558, 0.7222534, 0.7222739, 0.7222746, 0.7222733, 0.7222716, 
    0.72227, 0.7222678, 0.7222676, 0.7222672, 0.7222661, 0.7222652, 0.722267, 
    0.722265, 0.7222726, 0.7222686, 0.7222748, 0.722273, 0.7222717, 
    0.7222722, 0.7222693, 0.7222686, 0.7222657, 0.7222672, 0.7222584, 
    0.7222623, 0.7222516, 0.7222546, 0.7222748, 0.7222739, 0.7222705, 
    0.7222722, 0.7222676, 0.7222666, 0.7222656, 0.7222645, 0.7222643, 
    0.7222637, 0.7222648, 0.7222637, 0.7222677, 0.722266, 0.722271, 
    0.7222697, 0.7222703, 0.7222709, 0.722269, 0.722267, 0.722267, 0.7222663, 
    0.7222645, 0.7222676, 0.7222579, 0.7222639, 0.7222728, 0.722271, 
    0.7222707, 0.7222714, 0.7222666, 0.7222684, 0.7222637, 0.7222649, 
    0.7222629, 0.7222639, 0.7222641, 0.7222654, 0.7222662, 0.7222683, 
    0.72227, 0.7222713, 0.722271, 0.7222695, 0.7222669, 0.7222643, 0.7222649, 
    0.722263, 0.722268, 0.7222659, 0.7222667, 0.7222646, 0.7222692, 
    0.7222653, 0.7222702, 0.7222697, 0.7222684, 0.7222658, 0.7222652, 
    0.7222645, 0.7222649, 0.7222668, 0.7222671, 0.7222685, 0.7222688, 
    0.7222698, 0.7222707, 0.7222699, 0.7222691, 0.7222668, 0.7222648, 
    0.7222625, 0.7222619, 0.7222593, 0.7222614, 0.7222579, 0.7222609, 
    0.7222557, 0.7222651, 0.722261, 0.7222683, 0.7222676, 0.7222661, 
    0.7222629, 0.7222646, 0.7222626, 0.7222672, 0.7222695, 0.7222701, 
    0.7222713, 0.7222701, 0.7222702, 0.7222691, 0.7222694, 0.7222667, 
    0.7222682, 0.7222641, 0.7222626, 0.7222583, 0.7222557, 0.7222531, 
    0.7222519, 0.7222515, 0.7222514 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  3.083953e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 0, 5.139921e-21, 
    0, 1.541976e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 2.569961e-20, 
    -3.597945e-20, -1.541976e-20, 1.027984e-20, -2.055969e-20, -2.055969e-20, 
    -5.139921e-21, -2.055969e-20, -2.006177e-36, -1.027984e-20, 
    -5.139921e-21, -4.111937e-20, 2.055969e-20, -5.139921e-21, -3.597945e-20, 
    5.139921e-21, 2.055969e-20, 2.055969e-20, 0, -5.139921e-21, 
    -2.055969e-20, 2.055969e-20, -2.055969e-20, -2.569961e-20, -5.139921e-21, 
    -1.027984e-20, 2.055969e-20, 2.055969e-20, 1.541976e-20, 1.027984e-20, 
    -5.139921e-21, 3.597945e-20, -2.569961e-20, 5.139921e-21, 3.083953e-20, 
    5.139921e-21, 1.027984e-20, -1.027984e-20, -1.541976e-20, 2.569961e-20, 
    0, 0, 1.541976e-20, 0, -3.083953e-20, -1.027984e-20, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 1.541976e-20, -4.111937e-20, -3.083953e-20, 
    1.541976e-20, 2.055969e-20, -1.027984e-20, 1.541976e-20, 5.139921e-21, 
    -2.055969e-20, 2.569961e-20, -1.027984e-20, 1.027984e-20, -1.027984e-20, 
    1.541976e-20, 0, 1.541976e-20, 2.055969e-20, 0, -2.569961e-20, 
    -1.541976e-20, 3.083953e-20, -2.055969e-20, 2.006177e-36, -1.027984e-20, 
    -1.541976e-20, -5.139921e-21, 2.055969e-20, 3.083953e-20, 1.027984e-20, 
    -1.541976e-20, -5.139921e-21, 2.055969e-20, -2.055969e-20, -2.055969e-20, 
    -1.027984e-20, 2.055969e-20, 1.541976e-20, -2.055969e-20, 3.597945e-20, 
    1.541976e-20, -2.569961e-20, -3.597945e-20, -1.541976e-20, 2.055969e-20, 
    -5.139921e-21, -1.541976e-20, -1.027984e-20, -5.139921e-21, 
    -1.027984e-20, -1.027984e-20, -2.569961e-20, -2.006177e-36, 4.111937e-20, 
    2.055969e-20, -1.027984e-20, -1.027984e-20, 4.111937e-20, 1.027984e-20, 
    1.027984e-20, 2.006177e-36, -3.083953e-20, 5.139921e-21, -1.541976e-20, 
    2.055969e-20, 1.027984e-20, 1.541976e-20, -1.541976e-20, -1.027984e-20, 
    1.541976e-20, 1.027984e-20, 2.055969e-20, -1.541976e-20, 2.055969e-20, 
    5.139921e-21, 2.006177e-36, 1.027984e-20, 2.569961e-20, 5.139921e-21, 
    1.027984e-20, 2.055969e-20, 1.027984e-20, 2.055969e-20, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, -5.139921e-20, 5.139921e-21, 3.597945e-20, -2.569961e-20, 
    -1.027984e-20, 5.139921e-21, 2.569961e-20, 2.055969e-20, -1.541976e-20, 
    3.083953e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, 1.027984e-20, -1.027984e-20, -4.111937e-20, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 2.569961e-20, -2.055969e-20, -4.111937e-20, 
    -1.541976e-20, 1.541976e-20, -2.006177e-36, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, 0, -2.055969e-20, 
    1.541976e-20, 1.541976e-20, 1.541976e-20, 2.569961e-20, 3.597945e-20, 
    -5.139921e-21, 2.055969e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    1.027984e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, 3.083953e-20, -1.027984e-20, -2.055969e-20, 
    1.541976e-20, 1.027984e-20, -1.027984e-20, 2.006177e-36, 2.569961e-20, 
    -5.139921e-21, -3.597945e-20, -2.006177e-36, -1.027984e-20, 
    -1.027984e-20, 2.569961e-20, 1.541976e-20, -2.055969e-20, -1.541976e-20, 
    5.139921e-21, -1.027984e-20, 1.541976e-20, -2.006177e-36, 1.541976e-20, 
    1.027984e-20, -2.055969e-20, 3.597945e-20, 5.139921e-21, 4.625929e-20, 
    -1.541976e-20, 5.139921e-21, 3.083953e-20, 5.139921e-21, 5.139921e-21, 
    2.569961e-20, -2.569961e-20, -2.569961e-20, -5.139921e-21, -1.027984e-20, 
    -1.541976e-20, 5.139921e-21, -2.055969e-20, -1.027984e-20, 1.541976e-20, 
    2.569961e-20, -1.027984e-20, 5.139921e-21, -1.541976e-20, 1.541976e-20, 
    -3.083953e-20, 4.111937e-20, -1.027984e-20, 1.541976e-20, 2.569961e-20, 
    0, 2.006177e-36, -2.569961e-20, -1.027984e-20, -2.055969e-20, 
    1.541976e-20, 5.139921e-21, -3.597945e-20, -1.027984e-20, -2.569961e-20, 
    5.139921e-21, -1.027984e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, 
    0, 5.139921e-21, 1.027984e-20, 0, -1.541976e-20, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 0, 2.006177e-36, 1.541976e-20, 
    -5.139921e-20, -2.006177e-36, -3.083953e-20, -5.139921e-21, 3.083953e-20, 
    -3.597945e-20, -5.139921e-21, 1.541976e-20, 1.541976e-20, 2.055969e-20, 
    -4.111937e-20, -3.597945e-20, -1.541976e-20, 5.139921e-21, 2.055969e-20, 
    1.027984e-20, 2.055969e-20, -5.139921e-21, -1.027984e-20, 2.006177e-36, 
    -2.006177e-36, 1.027984e-20, 2.055969e-20, 2.055969e-20, 1.027984e-20, 
    2.055969e-20, 1.541976e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, 
    1.541976e-20, -2.055969e-20, -1.027984e-20, 0, -2.569961e-20, 
    1.027984e-20, -3.083953e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, -1.027984e-20, 1.541976e-20, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, -3.597945e-20, 
    5.139921e-21, 2.569961e-20, -2.569961e-20, 2.569961e-20, -2.569961e-20, 
    -5.139921e-21, -2.055969e-20, 0, -1.541976e-20, 3.597945e-20,
  -5.139921e-21, -2.569961e-20, -1.541976e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 0, -2.055969e-20, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 2.569961e-20, -2.006177e-36, 2.569961e-20, 
    2.569961e-20, 2.055969e-20, 1.541976e-20, 2.055969e-20, 1.541976e-20, 
    -1.027984e-20, 1.541976e-20, 0, -5.139921e-21, 0, 2.569961e-20, 
    1.027984e-20, -1.027984e-20, 5.139921e-21, 2.055969e-20, -5.139921e-21, 
    -2.055969e-20, 1.027984e-20, 0, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, 5.139921e-21, -2.006177e-36, -1.027984e-20, 3.083953e-20, 
    -5.139921e-21, 1.027984e-20, 5.139921e-21, -1.027984e-20, 0, 0, 
    5.139921e-21, 2.055969e-20, 1.541976e-20, -1.541976e-20, 0, 5.139921e-21, 
    5.139921e-21, 0, 1.541976e-20, 5.139921e-21, -2.055969e-20, 
    -5.139921e-21, -2.569961e-20, 3.083953e-20, -1.541976e-20, -1.541976e-20, 
    0, -1.027984e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -2.055969e-20, -1.541976e-20, -5.139921e-21, 1.027984e-20, -1.027984e-20, 
    0, 1.027984e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    1.541976e-20, 1.541976e-20, 1.027984e-20, -1.541976e-20, 0, 5.139921e-21, 
    5.139921e-21, -2.569961e-20, 3.083953e-20, 2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, -2.055969e-20, -1.027984e-20, 2.055969e-20, 
    -5.139921e-21, 1.027984e-20, 1.541976e-20, -1.027984e-20, 1.541976e-20, 
    0, 5.139921e-21, 1.541976e-20, -1.027984e-20, -1.541976e-20, 
    2.006177e-36, -5.139921e-21, 2.055969e-20, -1.027984e-20, 2.055969e-20, 
    3.083953e-20, -3.083953e-20, -1.027984e-20, 5.139921e-21, 0, 
    -1.027984e-20, -1.027984e-20, 3.597945e-20, 0, -1.541976e-20, 
    1.541976e-20, 0, 5.139921e-21, 0, -1.541976e-20, -1.027984e-20, 
    1.027984e-20, 3.083953e-20, -1.027984e-20, 5.139921e-21, 2.055969e-20, 
    -1.541976e-20, 0, 0, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -5.139921e-21, 0, -3.083953e-20, 1.541976e-20, -1.541976e-20, 
    2.569961e-20, -5.139921e-21, -5.139921e-21, 2.055969e-20, -5.139921e-21, 
    -1.541976e-20, -1.027984e-20, -3.083953e-20, 5.139921e-21, 2.569961e-20, 
    2.055969e-20, -1.027984e-20, 2.006177e-36, 0, 1.541976e-20, 0, 
    2.006177e-36, 1.541976e-20, 5.139921e-21, 0, 0, -5.139921e-21, 
    1.027984e-20, 2.055969e-20, -1.027984e-20, 1.541976e-20, -1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 5.139921e-21, 5.139921e-21, 1.541976e-20, 
    2.055969e-20, 5.139921e-21, 3.083953e-20, -1.541976e-20, 1.027984e-20, 
    1.541976e-20, 1.541976e-20, 1.027984e-20, -5.139921e-21, 1.541976e-20, 
    -1.027984e-20, 5.139921e-21, -3.597945e-20, -2.055969e-20, 1.027984e-20, 
    -2.569961e-20, 0, -2.569961e-20, -2.006177e-36, 1.027984e-20, 
    2.006177e-36, -1.541976e-20, 5.139921e-21, -1.541976e-20, -2.055969e-20, 
    -2.569961e-20, -2.055969e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    1.541976e-20, 1.027984e-20, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, -3.083953e-20, 1.541976e-20, 2.006177e-36, -1.027984e-20, 
    2.569961e-20, -1.541976e-20, 1.027984e-20, -1.541976e-20, -1.541976e-20, 
    3.597945e-20, 2.569961e-20, 2.006177e-36, -2.055969e-20, 0, 
    -1.027984e-20, 5.139921e-21, -2.055969e-20, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, 0, 0, -1.027984e-20, 0, 5.139921e-21, -1.541976e-20, 0, 
    1.541976e-20, -5.139921e-21, 5.139921e-21, -1.541976e-20, -1.541976e-20, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, 1.027984e-20, 
    0, -1.541976e-20, 0, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    2.055969e-20, -2.006177e-36, -1.541976e-20, 5.139921e-21, 2.055969e-20, 
    1.541976e-20, -5.139921e-21, 2.055969e-20, 5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 0, -1.541976e-20, 1.027984e-20, -1.541976e-20, 
    2.569961e-20, 1.541976e-20, -1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -1.541976e-20, 1.027984e-20, -3.083953e-20, 
    5.139921e-21, -2.055969e-20, -5.139921e-21, 0, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, -2.055969e-20, 1.027984e-20, -1.541976e-20, 
    0, 1.541976e-20, 0, -2.569961e-20, -1.541976e-20, -1.027984e-20, 0, 
    5.139921e-21, -2.569961e-20, -1.027984e-20, 0, -2.055969e-20, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, -1.541976e-20, 
    0, 2.569961e-20, 2.569961e-20, -5.139921e-21, 1.027984e-20, 
    -2.569961e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, -1.541976e-20, 
    2.006177e-36, 0, -2.006177e-36, 1.027984e-20, 5.139921e-21, 3.083953e-20, 
    -3.083953e-20, 5.139921e-21, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    -2.055969e-20, 5.139921e-21, 3.083953e-20, -1.541976e-20, 1.541976e-20, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, -1.027984e-20, -1.541976e-20, 
    5.139921e-21, -5.139921e-21, 5.139921e-21,
  -1.027984e-20, -1.027984e-20, -5.139921e-21, 1.541976e-20, 2.569961e-20, 
    1.027984e-20, -1.541976e-20, -5.139921e-21, 3.083953e-20, -1.027984e-20, 
    1.541976e-20, -1.027984e-20, 5.139921e-21, 2.055969e-20, 0, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -5.139921e-20, -2.055969e-20, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, 1.027984e-20, -1.027984e-20, 2.006177e-36, 
    0, 0, 1.027984e-20, 1.027984e-20, -1.027984e-20, 2.006177e-36, 
    -2.569961e-20, -1.541976e-20, 5.139921e-21, 1.541976e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 0, -2.569961e-20, 0, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    -1.027984e-20, 5.139921e-21, -1.027984e-20, 2.569961e-20, -1.541976e-20, 
    1.027984e-20, 2.006177e-36, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -3.597945e-20, -5.139921e-21, -1.027984e-20, 2.006177e-36, 1.027984e-20, 
    -1.027984e-20, 2.055969e-20, 1.541976e-20, -1.027984e-20, 0, 
    1.541976e-20, 2.055969e-20, -1.027984e-20, 1.541976e-20, -5.139921e-21, 
    -1.541976e-20, -1.027984e-20, -1.027984e-20, -1.027984e-20, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, -5.139921e-21, 1.027984e-20, 1.541976e-20, 
    3.083953e-20, 2.569961e-20, -2.006177e-36, 2.569961e-20, 2.569961e-20, 
    -2.569961e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 0, 0, 
    -1.027984e-20, -5.139921e-21, 5.139921e-21, -4.111937e-20, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, 1.541976e-20, -5.139921e-21, -2.006177e-36, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, -2.569961e-20, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -2.055969e-20, 1.027984e-20, -1.541976e-20, 
    -2.569961e-20, 2.006177e-36, -4.625929e-20, -1.027984e-20, -3.597945e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, -1.541976e-20, 2.006177e-36, 5.139921e-21, -1.027984e-20, 
    -1.541976e-20, 5.139921e-21, 3.597945e-20, 2.006177e-36, -1.027984e-20, 
    -3.597945e-20, 3.083953e-20, 1.027984e-20, -1.541976e-20, -1.027984e-20, 
    -1.027984e-20, 2.006177e-36, 3.083953e-20, 2.569961e-20, -3.083953e-20, 
    1.027984e-20, -5.139921e-21, 2.055969e-20, -3.083953e-20, 2.055969e-20, 
    -2.055969e-20, 1.541976e-20, -1.541976e-20, 5.139921e-21, -2.055969e-20, 
    -1.027984e-20, 2.569961e-20, -1.027984e-20, -1.027984e-20, -2.569961e-20, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 0, 
    1.027984e-20, -3.083953e-20, -1.027984e-20, 5.139921e-21, -2.006177e-36, 
    -1.027984e-20, -5.139921e-21, -5.139921e-21, 2.569961e-20, 0, 
    1.541976e-20, -1.027984e-20, 5.139921e-21, 2.569961e-20, 3.597945e-20, 
    -2.055969e-20, -1.541976e-20, 1.027984e-20, -2.055969e-20, 0, 
    2.006177e-36, 5.139921e-21, -3.083953e-20, 2.006177e-36, 5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 2.569961e-20, -5.139921e-21, -1.027984e-20, 
    3.597945e-20, 5.139921e-21, -1.541976e-20, 1.027984e-20, 1.027984e-20, 
    -1.541976e-20, 2.055969e-20, -2.055969e-20, 2.055969e-20, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, -1.541976e-20, -3.083953e-20, 5.139921e-21, 
    -2.055969e-20, 1.027984e-20, 1.027984e-20, -2.055969e-20, -2.006177e-36, 
    -1.027984e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -3.083953e-20, 5.139921e-21, 0, -1.027984e-20, 0, -2.055969e-20, 
    -4.111937e-20, 3.597945e-20, 2.006177e-36, -1.027984e-20, -5.139921e-21, 
    1.541976e-20, -2.055969e-20, 1.541976e-20, -3.083953e-20, -1.027984e-20, 
    -1.541976e-20, 2.006177e-36, -5.139921e-21, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 1.541976e-20, 5.139921e-21, 1.027984e-20, 
    2.569961e-20, 5.139921e-21, 1.027984e-20, 0, -1.027984e-20, 
    -2.055969e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    2.055969e-20, 5.139921e-21, -1.027984e-20, -1.027984e-20, 0, 
    1.027984e-20, 1.541976e-20, 3.083953e-20, 1.027984e-20, -2.006177e-36, 
    1.541976e-20, -5.139921e-21, -1.541976e-20, 2.006177e-36, 2.569961e-20, 
    -2.006177e-36, -1.027984e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, -1.027984e-20, -2.055969e-20, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, 1.027984e-20, 0, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, 1.541976e-20, 1.541976e-20, 
    1.027984e-20, -2.569961e-20, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    0, -1.541976e-20, -1.541976e-20, -1.027984e-20, -1.027984e-20, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, -1.027984e-20, 1.541976e-20, 
    1.541976e-20, -1.027984e-20, 3.597945e-20, 3.083953e-20, -2.055969e-20, 
    -2.055969e-20, 2.055969e-20, 1.541976e-20, -2.055969e-20, 4.111937e-20, 
    1.027984e-20, 1.541976e-20, -1.027984e-20, -2.569961e-20, 1.541976e-20, 
    -5.139921e-21, -1.541976e-20, 1.541976e-20, 1.027984e-20, 1.027984e-20, 
    1.027984e-20, 1.541976e-20, 2.569961e-20, -1.027984e-20, 2.055969e-20, 
    1.027984e-20, 1.027984e-20, -1.541976e-20, -1.541976e-20, 5.139921e-21, 
    5.139921e-21, -1.027984e-20, -5.139921e-21,
  1.027984e-20, -2.055969e-20, -2.055969e-20, 1.541976e-20, 5.139921e-21, 
    -5.139921e-21, 0, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, -2.569961e-20, 5.139921e-21, 2.055969e-20, 
    1.541976e-20, -1.027984e-20, -1.027984e-20, -2.569961e-20, 1.027984e-20, 
    0, 2.055969e-20, 3.083953e-20, -5.139921e-21, -2.569961e-20, 
    5.139921e-21, -4.625929e-20, 2.055969e-20, -1.541976e-20, 2.569961e-20, 
    -1.541976e-20, 1.541976e-20, 0, 2.006177e-36, -2.006177e-36, 
    -5.139921e-21, -2.006177e-36, -5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -2.006177e-36, -1.541976e-20, 1.027984e-20, 0, 
    -1.027984e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, 
    -2.055969e-20, 4.111937e-20, 5.139921e-21, -5.139921e-21, 2.006177e-36, 
    -4.111937e-20, -2.055969e-20, -1.541976e-20, 2.055969e-20, 1.027984e-20, 
    2.569961e-20, -3.597945e-20, 2.006177e-36, 5.139921e-21, 2.569961e-20, 
    2.055969e-20, 1.027984e-20, -5.139921e-21, 0, 0, 2.569961e-20, 
    -5.139921e-21, -1.027984e-20, 1.027984e-20, -5.139921e-21, 1.541976e-20, 
    -2.055969e-20, 1.027984e-20, 2.569961e-20, 0, -2.569961e-20, 
    1.541976e-20, -2.055969e-20, 5.139921e-21, 1.027984e-20, -1.541976e-20, 
    1.541976e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 0, 
    -2.569961e-20, -1.541976e-20, -2.569961e-20, -1.541976e-20, 1.541976e-20, 
    2.569961e-20, 3.083953e-20, -4.111937e-20, -5.139921e-21, 5.139921e-21, 
    -2.006177e-36, -1.541976e-20, 2.055969e-20, 2.055969e-20, 0, 
    1.027984e-20, 1.541976e-20, -2.055969e-20, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, -3.597945e-20, -2.006177e-36, 
    -1.541976e-20, -4.111937e-20, 1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -1.541976e-20, -2.569961e-20, -5.139921e-21, 2.006177e-36, -1.541976e-20, 
    2.055969e-20, -1.027984e-20, 2.055969e-20, 1.541976e-20, -1.027984e-20, 
    -2.055969e-20, 2.055969e-20, 1.027984e-20, 0, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 2.055969e-20, 2.055969e-20, -2.055969e-20, 1.027984e-20, 
    -2.006177e-36, -1.541976e-20, -5.139921e-21, -1.027984e-20, 1.541976e-20, 
    -1.541976e-20, -1.027984e-20, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, -3.083953e-20, 5.139921e-21, -2.569961e-20, 2.006177e-36, 
    5.139921e-21, 2.569961e-20, -5.139921e-21, 5.139921e-21, -2.569961e-20, 
    -2.055969e-20, -5.139921e-21, 4.111937e-20, -5.139921e-21, 2.055969e-20, 
    1.027984e-20, 2.055969e-20, -1.541976e-20, 1.541976e-20, 5.139921e-21, 
    5.139921e-21, 3.083953e-20, 4.625929e-20, 5.139921e-21, 4.625929e-20, 
    -1.027984e-20, 5.139921e-21, 3.083953e-20, 1.027984e-20, -1.541976e-20, 
    1.027984e-20, 5.139921e-21, 2.569961e-20, 1.027984e-20, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -2.569961e-20, 5.139921e-21, -2.055969e-20, -2.006177e-36, 3.083953e-20, 
    3.597945e-20, -3.083953e-20, 3.597945e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -1.541976e-20, -3.083953e-20, -2.055969e-20, 
    2.055969e-20, 1.027984e-20, -2.006177e-36, 2.569961e-20, 0, 1.027984e-20, 
    5.139921e-21, -2.569961e-20, -3.083953e-20, -2.055969e-20, -2.055969e-20, 
    -1.027984e-20, 1.027984e-20, 2.569961e-20, -5.139921e-21, -4.625929e-20, 
    1.027984e-20, -1.541976e-20, 0, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -2.006177e-36, -2.055969e-20, 
    -2.006177e-36, -5.139921e-21, -2.055969e-20, -1.027984e-20, 1.027984e-20, 
    -2.006177e-36, 5.139921e-21, -1.027984e-20, 1.541976e-20, 1.541976e-20, 
    -1.541976e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 0, 
    5.139921e-21, 1.541976e-20, 2.569961e-20, -2.569961e-20, -4.111937e-20, 
    -2.006177e-36, 5.139921e-21, 1.541976e-20, 2.569961e-20, -4.625929e-20, 
    -2.055969e-20, -1.027984e-20, 4.111937e-20, -2.055969e-20, -1.027984e-20, 
    1.027984e-20, 1.541976e-20, 0, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    -1.027984e-20, -3.597945e-20, 2.055969e-20, 3.597945e-20, 0, 
    -1.541976e-20, 3.597945e-20, 2.006177e-36, -2.055969e-20, -5.139921e-21, 
    2.569961e-20, 1.541976e-20, 5.139921e-21, 1.027984e-20, -2.006177e-36, 
    -2.055969e-20, -5.139921e-21, -5.139921e-21, -1.541976e-20, 2.569961e-20, 
    1.541976e-20, 2.006177e-36, -5.653913e-20, 1.541976e-20, -5.139921e-21, 
    -2.055969e-20, 2.569961e-20, 1.541976e-20, -2.055969e-20, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, -1.541976e-20, 1.541976e-20, 0, 
    -1.027984e-20, 2.055969e-20, 0, -1.027984e-20, -5.139921e-21, 0, 
    2.569961e-20, -1.541976e-20, 1.541976e-20, -2.006177e-36, -1.027984e-20, 
    1.541976e-20, -2.569961e-20, 5.139921e-21, 0, -5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 2.569961e-20, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, 2.055969e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -2.569961e-20, 1.541976e-20, 5.139921e-21, -2.055969e-20, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21,
  -1.027984e-20, 5.139921e-21, 0, -1.541976e-20, 1.541976e-20, 5.139921e-21, 
    -2.569961e-20, 2.006177e-36, 5.139921e-21, -1.027984e-20, 2.569961e-20, 
    -1.027984e-20, 1.541976e-20, 1.027984e-20, -1.541976e-20, 1.027984e-20, 
    1.027984e-20, -1.541976e-20, -5.139921e-21, -4.111937e-20, 1.027984e-20, 
    5.139921e-21, 2.055969e-20, -1.541976e-20, 2.055969e-20, 1.541976e-20, 0, 
    0, 1.027984e-20, 5.139921e-21, 5.139921e-21, 1.541976e-20, -1.541976e-20, 
    1.541976e-20, 1.541976e-20, -1.541976e-20, 3.597945e-20, 2.055969e-20, 
    -1.027984e-20, 5.139921e-21, 2.569961e-20, -5.139921e-21, -2.055969e-20, 
    2.006177e-36, -5.139921e-21, 1.027984e-20, 5.139921e-21, 2.055969e-20, 
    -5.139921e-21, -2.055969e-20, 0, -3.083953e-20, -2.569961e-20, 
    -5.139921e-21, 1.027984e-20, -1.027984e-20, -4.111937e-20, 3.083953e-20, 
    1.541976e-20, -1.027984e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, 
    1.541976e-20, -1.541976e-20, 0, 2.055969e-20, 5.139921e-21, 
    -2.569961e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 1.027984e-20, 
    1.541976e-20, -2.006177e-36, -1.027984e-20, 2.569961e-20, -1.541976e-20, 
    -2.569961e-20, -1.541976e-20, 2.055969e-20, 0, -5.139921e-21, 
    -1.541976e-20, 2.569961e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    -2.055969e-20, -2.569961e-20, -2.055969e-20, 3.083953e-20, -2.006177e-36, 
    -1.027984e-20, -2.055969e-20, 2.055969e-20, -3.083953e-20, -2.055969e-20, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, -2.006177e-36, -1.027984e-20, 2.055969e-20, 
    -2.569961e-20, 5.139921e-21, -5.139921e-21, 0, 1.027984e-20, 
    -2.055969e-20, 5.139921e-21, -1.027984e-20, -2.055969e-20, 3.597945e-20, 
    1.541976e-20, -1.027984e-20, 0, -1.027984e-20, -1.541976e-20, 
    -2.055969e-20, 2.055969e-20, 2.055969e-20, 2.569961e-20, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, -5.653913e-20, 2.055969e-20, 
    -2.569961e-20, 5.139921e-21, -1.027984e-20, 3.083953e-20, 2.055969e-20, 
    3.083953e-20, 2.569961e-20, -5.139921e-21, 1.027984e-20, 3.597945e-20, 
    -5.139921e-20, 5.139921e-21, 5.139921e-21, 2.055969e-20, -1.541976e-20, 
    2.569961e-20, -2.055969e-20, 4.625929e-20, 1.541976e-20, 3.083953e-20, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, -2.569961e-20, 1.027984e-20, 
    5.139921e-21, 2.569961e-20, -1.027984e-20, -1.541976e-20, -2.006177e-36, 
    0, 5.139921e-21, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, -4.625929e-20, -1.027984e-20, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 1.541976e-20, -2.569961e-20, 4.625929e-20, -3.083953e-20, 
    0, 2.006177e-36, 1.541976e-20, 3.083953e-20, 3.083953e-20, 1.027984e-20, 
    -2.569961e-20, -1.541976e-20, 1.027984e-20, 2.055969e-20, -1.027984e-20, 
    -2.055969e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, -2.055969e-20, 0, 2.055969e-20, -2.055969e-20, 
    -2.055969e-20, -1.541976e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, 
    -2.569961e-20, -1.541976e-20, -2.006177e-36, -1.541976e-20, 1.027984e-20, 
    -1.541976e-20, -5.139921e-21, 1.027984e-20, -2.055969e-20, 1.027984e-20, 
    -1.027984e-20, 5.139921e-21, 2.569961e-20, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 5.139921e-21, -2.055969e-20, 3.083953e-20, 
    0, -1.027984e-20, -5.139921e-21, 2.569961e-20, 2.055969e-20, 
    2.055969e-20, -5.139921e-21, -3.083953e-20, -1.541976e-20, 2.055969e-20, 
    0, 2.055969e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    -1.541976e-20, 2.569961e-20, 1.541976e-20, 2.055969e-20, 1.027984e-20, 
    -1.027984e-20, 2.569961e-20, 5.139921e-21, -2.055969e-20, 5.139921e-21, 
    -5.139921e-21, 2.055969e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    2.055969e-20, 5.139921e-21, 3.083953e-20, 2.569961e-20, -2.569961e-20, 0, 
    -5.139921e-21, 2.055969e-20, 1.541976e-20, -1.027984e-20, 3.597945e-20, 
    -2.569961e-20, 1.541976e-20, -5.139921e-21, 3.083953e-20, -3.597945e-20, 
    -2.006177e-36, 1.541976e-20, 2.055969e-20, -2.569961e-20, -2.006177e-36, 
    -5.139921e-21, 5.139921e-21, 0, -2.055969e-20, -1.027984e-20, 
    -5.139921e-21, 0, 5.139921e-21, 2.569961e-20, -2.569961e-20, 
    5.139921e-21, 2.006177e-36, -1.027984e-20, -1.027984e-20, -1.027984e-20, 
    1.541976e-20, 1.541976e-20, 1.541976e-20, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 3.597945e-20, 
    -4.111937e-20, 1.541976e-20, 3.083953e-20, 1.541976e-20, 1.027984e-20, 
    -1.027984e-20, -2.055969e-20, -1.027984e-20, -1.027984e-20, 2.055969e-20, 
    2.569961e-20, 2.055969e-20, 0, 2.055969e-20, -2.006177e-36, 
    -2.055969e-20, -1.541976e-20, 5.139921e-21, 5.139921e-21, 0, 
    -1.027984e-20, 1.541976e-20, -5.139921e-21, 0, -1.541976e-20, 
    -2.055969e-20, 3.597945e-20, 2.055969e-20, -2.055969e-20, 1.541976e-20, 
    5.139921e-21, 2.569961e-20, -5.139921e-21, 5.139921e-21, -1.541976e-20, 
    -3.597945e-20, 1.027984e-20,
  8.598827e-29, 8.598799e-29, 8.598805e-29, 8.598782e-29, 8.598795e-29, 
    8.598779e-29, 8.598822e-29, 8.598798e-29, 8.598813e-29, 8.598825e-29, 
    8.598739e-29, 8.598781e-29, 8.598694e-29, 8.598721e-29, 8.598652e-29, 
    8.598698e-29, 8.598643e-29, 8.598654e-29, 8.598622e-29, 8.598631e-29, 
    8.598591e-29, 8.598618e-29, 8.59857e-29, 8.598597e-29, 8.598593e-29, 
    8.598619e-29, 8.598772e-29, 8.598743e-29, 8.598774e-29, 8.59877e-29, 
    8.598772e-29, 8.598794e-29, 8.598805e-29, 8.598829e-29, 8.598825e-29, 
    8.598808e-29, 8.598768e-29, 8.598781e-29, 8.598748e-29, 8.598749e-29, 
    8.598711e-29, 8.598728e-29, 8.598665e-29, 8.598683e-29, 8.598631e-29, 
    8.598644e-29, 8.598631e-29, 8.598635e-29, 8.598631e-29, 8.598651e-29, 
    8.598642e-29, 8.598659e-29, 8.598725e-29, 8.598705e-29, 8.598763e-29, 
    8.598798e-29, 8.59882e-29, 8.598837e-29, 8.598834e-29, 8.59883e-29, 
    8.598807e-29, 8.598786e-29, 8.59877e-29, 8.59876e-29, 8.598749e-29, 
    8.598716e-29, 8.598699e-29, 8.598662e-29, 8.598668e-29, 8.598657e-29, 
    8.598645e-29, 8.598627e-29, 8.59863e-29, 8.598621e-29, 8.598657e-29, 
    8.598633e-29, 8.598672e-29, 8.598662e-29, 8.598746e-29, 8.598778e-29, 
    8.598792e-29, 8.598804e-29, 8.598832e-29, 8.598813e-29, 8.59882e-29, 
    8.598802e-29, 8.59879e-29, 8.598796e-29, 8.598759e-29, 8.598773e-29, 
    8.598698e-29, 8.598731e-29, 8.598646e-29, 8.598667e-29, 8.598642e-29, 
    8.598654e-29, 8.598633e-29, 8.598652e-29, 8.598618e-29, 8.598611e-29, 
    8.598616e-29, 8.598597e-29, 8.598654e-29, 8.598631e-29, 8.598796e-29, 
    8.598795e-29, 8.59879e-29, 8.59881e-29, 8.598811e-29, 8.598829e-29, 
    8.598813e-29, 8.598807e-29, 8.598789e-29, 8.598779e-29, 8.598769e-29, 
    8.598748e-29, 8.598723e-29, 8.59869e-29, 8.598665e-29, 8.598649e-29, 
    8.598659e-29, 8.59865e-29, 8.59866e-29, 8.598665e-29, 8.598613e-29, 
    8.598642e-29, 8.5986e-29, 8.598602e-29, 8.598621e-29, 8.598601e-29, 
    8.598794e-29, 8.598799e-29, 8.598819e-29, 8.598804e-29, 8.598831e-29, 
    8.598816e-29, 8.598807e-29, 8.598773e-29, 8.598766e-29, 8.598758e-29, 
    8.598745e-29, 8.598727e-29, 8.598696e-29, 8.598669e-29, 8.598645e-29, 
    8.598646e-29, 8.598646e-29, 8.59864e-29, 8.598654e-29, 8.598638e-29, 
    8.598636e-29, 8.598642e-29, 8.598602e-29, 8.598613e-29, 8.598602e-29, 
    8.598609e-29, 8.598798e-29, 8.598788e-29, 8.598793e-29, 8.598784e-29, 
    8.598791e-29, 8.598761e-29, 8.598752e-29, 8.59871e-29, 8.598728e-29, 
    8.5987e-29, 8.598725e-29, 8.59872e-29, 8.598699e-29, 8.598723e-29, 
    8.598671e-29, 8.598707e-29, 8.59864e-29, 8.598676e-29, 8.598638e-29, 
    8.598645e-29, 8.598633e-29, 8.598623e-29, 8.59861e-29, 8.598586e-29, 
    8.598592e-29, 8.598572e-29, 8.598775e-29, 8.598763e-29, 8.598763e-29, 
    8.598751e-29, 8.598742e-29, 8.598721e-29, 8.598689e-29, 8.598701e-29, 
    8.598678e-29, 8.598674e-29, 8.598708e-29, 8.598687e-29, 8.598754e-29, 
    8.598743e-29, 8.59875e-29, 8.598773e-29, 8.598698e-29, 8.598737e-29, 
    8.598665e-29, 8.598686e-29, 8.598625e-29, 8.598655e-29, 8.598595e-29, 
    8.598569e-29, 8.598545e-29, 8.598516e-29, 8.598756e-29, 8.598764e-29, 
    8.598749e-29, 8.598729e-29, 8.59871e-29, 8.598685e-29, 8.598682e-29, 
    8.598678e-29, 8.598665e-29, 8.598655e-29, 8.598676e-29, 8.598652e-29, 
    8.598741e-29, 8.598695e-29, 8.598767e-29, 8.598745e-29, 8.59873e-29, 
    8.598737e-29, 8.598702e-29, 8.598694e-29, 8.598661e-29, 8.598678e-29, 
    8.598575e-29, 8.598621e-29, 8.598495e-29, 8.59853e-29, 8.598767e-29, 
    8.598756e-29, 8.598717e-29, 8.598736e-29, 8.598683e-29, 8.59867e-29, 
    8.59866e-29, 8.598646e-29, 8.598645e-29, 8.598637e-29, 8.59865e-29, 
    8.598637e-29, 8.598685e-29, 8.598663e-29, 8.598722e-29, 8.598707e-29, 
    8.598714e-29, 8.598721e-29, 8.598699e-29, 8.598676e-29, 8.598675e-29, 
    8.598668e-29, 8.598646e-29, 8.598683e-29, 8.59857e-29, 8.59864e-29, 
    8.598744e-29, 8.598722e-29, 8.598719e-29, 8.598728e-29, 8.598672e-29, 
    8.598692e-29, 8.598637e-29, 8.598652e-29, 8.598627e-29, 8.59864e-29, 
    8.598642e-29, 8.598657e-29, 8.598666e-29, 8.598691e-29, 8.598711e-29, 
    8.598727e-29, 8.598723e-29, 8.598705e-29, 8.598674e-29, 8.598645e-29, 
    8.598651e-29, 8.59863e-29, 8.598687e-29, 8.598663e-29, 8.598672e-29, 
    8.598648e-29, 8.598701e-29, 8.598655e-29, 8.598713e-29, 8.598708e-29, 
    8.598692e-29, 8.598661e-29, 8.598654e-29, 8.598647e-29, 8.598651e-29, 
    8.598674e-29, 8.598677e-29, 8.598693e-29, 8.598697e-29, 8.598709e-29, 
    8.598719e-29, 8.59871e-29, 8.5987e-29, 8.598674e-29, 8.598649e-29, 
    8.598623e-29, 8.598616e-29, 8.598586e-29, 8.598611e-29, 8.598569e-29, 
    8.598604e-29, 8.598544e-29, 8.598653e-29, 8.598606e-29, 8.598692e-29, 
    8.598683e-29, 8.598666e-29, 8.598627e-29, 8.598648e-29, 8.598624e-29, 
    8.598677e-29, 8.598705e-29, 8.598712e-29, 8.598725e-29, 8.598712e-29, 
    8.598713e-29, 8.5987e-29, 8.598704e-29, 8.598672e-29, 8.598689e-29, 
    8.598642e-29, 8.598624e-29, 8.598574e-29, 8.598544e-29, 8.598513e-29, 
    8.598499e-29, 8.598495e-29, 8.598493e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.135276e-08, 1.140281e-08, 1.139308e-08, 1.143345e-08, 1.141105e-08, 
    1.143749e-08, 1.136291e-08, 1.140479e-08, 1.137805e-08, 1.135727e-08, 
    1.151178e-08, 1.143525e-08, 1.15913e-08, 1.154248e-08, 1.166513e-08, 
    1.158371e-08, 1.168155e-08, 1.166278e-08, 1.171927e-08, 1.170308e-08, 
    1.177533e-08, 1.172674e-08, 1.181279e-08, 1.176373e-08, 1.17714e-08, 
    1.172513e-08, 1.145065e-08, 1.150225e-08, 1.144759e-08, 1.145495e-08, 
    1.145165e-08, 1.141152e-08, 1.139129e-08, 1.134894e-08, 1.135662e-08, 
    1.138773e-08, 1.145826e-08, 1.143432e-08, 1.149466e-08, 1.14933e-08, 
    1.156048e-08, 1.153019e-08, 1.164311e-08, 1.161101e-08, 1.170376e-08, 
    1.168043e-08, 1.170266e-08, 1.169592e-08, 1.170275e-08, 1.166854e-08, 
    1.16832e-08, 1.16531e-08, 1.153586e-08, 1.157031e-08, 1.146756e-08, 
    1.140577e-08, 1.136474e-08, 1.133563e-08, 1.133974e-08, 1.134759e-08, 
    1.138791e-08, 1.142583e-08, 1.145473e-08, 1.147406e-08, 1.14931e-08, 
    1.155075e-08, 1.158127e-08, 1.16496e-08, 1.163727e-08, 1.165815e-08, 
    1.167811e-08, 1.171162e-08, 1.170611e-08, 1.172087e-08, 1.165761e-08, 
    1.169965e-08, 1.163024e-08, 1.164923e-08, 1.149827e-08, 1.144078e-08, 
    1.141634e-08, 1.139495e-08, 1.134291e-08, 1.137885e-08, 1.136468e-08, 
    1.139838e-08, 1.14198e-08, 1.140921e-08, 1.147459e-08, 1.144917e-08, 
    1.158307e-08, 1.152539e-08, 1.167579e-08, 1.16398e-08, 1.168441e-08, 
    1.166165e-08, 1.170065e-08, 1.166555e-08, 1.172636e-08, 1.173961e-08, 
    1.173056e-08, 1.176532e-08, 1.16636e-08, 1.170266e-08, 1.140891e-08, 
    1.141064e-08, 1.141869e-08, 1.138331e-08, 1.138114e-08, 1.134872e-08, 
    1.137757e-08, 1.138986e-08, 1.142104e-08, 1.143949e-08, 1.145703e-08, 
    1.149558e-08, 1.153864e-08, 1.159886e-08, 1.164213e-08, 1.167113e-08, 
    1.165335e-08, 1.166905e-08, 1.16515e-08, 1.164327e-08, 1.173464e-08, 
    1.168334e-08, 1.176032e-08, 1.175606e-08, 1.172122e-08, 1.175654e-08, 
    1.141185e-08, 1.140191e-08, 1.13674e-08, 1.139441e-08, 1.134519e-08, 
    1.137274e-08, 1.138858e-08, 1.14497e-08, 1.146313e-08, 1.147558e-08, 
    1.150017e-08, 1.153174e-08, 1.158711e-08, 1.163529e-08, 1.167928e-08, 
    1.167605e-08, 1.167719e-08, 1.168701e-08, 1.166267e-08, 1.169101e-08, 
    1.169576e-08, 1.168333e-08, 1.175549e-08, 1.173487e-08, 1.175597e-08, 
    1.174255e-08, 1.140514e-08, 1.142187e-08, 1.141283e-08, 1.142983e-08, 
    1.141785e-08, 1.14711e-08, 1.148707e-08, 1.156177e-08, 1.153112e-08, 
    1.157991e-08, 1.153607e-08, 1.154384e-08, 1.15815e-08, 1.153844e-08, 
    1.163263e-08, 1.156877e-08, 1.168739e-08, 1.162362e-08, 1.169139e-08, 
    1.167909e-08, 1.169946e-08, 1.171771e-08, 1.174067e-08, 1.178303e-08, 
    1.177322e-08, 1.180865e-08, 1.144681e-08, 1.146851e-08, 1.14666e-08, 
    1.14893e-08, 1.15061e-08, 1.15425e-08, 1.160088e-08, 1.157893e-08, 
    1.161923e-08, 1.162732e-08, 1.156609e-08, 1.160369e-08, 1.148303e-08, 
    1.150252e-08, 1.149091e-08, 1.144852e-08, 1.158398e-08, 1.151446e-08, 
    1.164284e-08, 1.160518e-08, 1.171511e-08, 1.166044e-08, 1.176782e-08, 
    1.181373e-08, 1.185694e-08, 1.190743e-08, 1.148035e-08, 1.146561e-08, 
    1.1492e-08, 1.152853e-08, 1.156242e-08, 1.160748e-08, 1.161209e-08, 
    1.162053e-08, 1.164239e-08, 1.166078e-08, 1.16232e-08, 1.166539e-08, 
    1.150704e-08, 1.159002e-08, 1.146003e-08, 1.149917e-08, 1.152637e-08, 
    1.151444e-08, 1.157642e-08, 1.159103e-08, 1.165038e-08, 1.16197e-08, 
    1.180239e-08, 1.172156e-08, 1.194588e-08, 1.188319e-08, 1.146045e-08, 
    1.14803e-08, 1.154936e-08, 1.15165e-08, 1.161049e-08, 1.163362e-08, 
    1.165243e-08, 1.167647e-08, 1.167906e-08, 1.169331e-08, 1.166997e-08, 
    1.169239e-08, 1.160757e-08, 1.164547e-08, 1.154147e-08, 1.156678e-08, 
    1.155514e-08, 1.154237e-08, 1.158179e-08, 1.162379e-08, 1.162469e-08, 
    1.163815e-08, 1.16761e-08, 1.161087e-08, 1.181282e-08, 1.168809e-08, 
    1.150194e-08, 1.154016e-08, 1.154562e-08, 1.153081e-08, 1.16313e-08, 
    1.159489e-08, 1.169296e-08, 1.166646e-08, 1.170989e-08, 1.16883e-08, 
    1.168513e-08, 1.165741e-08, 1.164016e-08, 1.159656e-08, 1.156109e-08, 
    1.153296e-08, 1.15395e-08, 1.15704e-08, 1.162636e-08, 1.16793e-08, 
    1.16677e-08, 1.170659e-08, 1.160367e-08, 1.164682e-08, 1.163014e-08, 
    1.167363e-08, 1.157834e-08, 1.165948e-08, 1.15576e-08, 1.156654e-08, 
    1.159417e-08, 1.164975e-08, 1.166205e-08, 1.167518e-08, 1.166708e-08, 
    1.162778e-08, 1.162134e-08, 1.15935e-08, 1.158581e-08, 1.156459e-08, 
    1.154703e-08, 1.156307e-08, 1.157993e-08, 1.162779e-08, 1.167093e-08, 
    1.171797e-08, 1.172948e-08, 1.178443e-08, 1.17397e-08, 1.181352e-08, 
    1.175075e-08, 1.185941e-08, 1.166419e-08, 1.174891e-08, 1.159543e-08, 
    1.161196e-08, 1.164186e-08, 1.171046e-08, 1.167343e-08, 1.171674e-08, 
    1.162109e-08, 1.157146e-08, 1.155863e-08, 1.153467e-08, 1.155917e-08, 
    1.155718e-08, 1.158063e-08, 1.157309e-08, 1.162938e-08, 1.159915e-08, 
    1.168505e-08, 1.17164e-08, 1.180493e-08, 1.185921e-08, 1.191447e-08, 
    1.193887e-08, 1.194629e-08, 1.194939e-08 ;

 SOIL1N_TO_SOIL3N =
  1.347056e-10, 1.352997e-10, 1.351842e-10, 1.356634e-10, 1.353976e-10, 
    1.357113e-10, 1.348261e-10, 1.353233e-10, 1.350059e-10, 1.347591e-10, 
    1.365932e-10, 1.356847e-10, 1.375371e-10, 1.369577e-10, 1.384134e-10, 
    1.374469e-10, 1.386083e-10, 1.383856e-10, 1.390561e-10, 1.38864e-10, 
    1.397216e-10, 1.391448e-10, 1.401663e-10, 1.395839e-10, 1.39675e-10, 
    1.391258e-10, 1.358676e-10, 1.364801e-10, 1.358313e-10, 1.359186e-10, 
    1.358794e-10, 1.35403e-10, 1.35163e-10, 1.346603e-10, 1.347515e-10, 
    1.351208e-10, 1.359579e-10, 1.356738e-10, 1.3639e-10, 1.363738e-10, 
    1.371712e-10, 1.368117e-10, 1.381521e-10, 1.377711e-10, 1.38872e-10, 
    1.385951e-10, 1.38859e-10, 1.38779e-10, 1.388601e-10, 1.38454e-10, 
    1.38628e-10, 1.382707e-10, 1.36879e-10, 1.37288e-10, 1.360683e-10, 
    1.353349e-10, 1.348479e-10, 1.345023e-10, 1.345511e-10, 1.346443e-10, 
    1.351229e-10, 1.35573e-10, 1.35916e-10, 1.361454e-10, 1.363715e-10, 
    1.370557e-10, 1.37418e-10, 1.382291e-10, 1.380827e-10, 1.383307e-10, 
    1.385676e-10, 1.389654e-10, 1.388999e-10, 1.390751e-10, 1.383242e-10, 
    1.388232e-10, 1.379994e-10, 1.382247e-10, 1.364329e-10, 1.357504e-10, 
    1.354603e-10, 1.352064e-10, 1.345887e-10, 1.350153e-10, 1.348471e-10, 
    1.352472e-10, 1.355014e-10, 1.353757e-10, 1.361517e-10, 1.3585e-10, 
    1.374395e-10, 1.367548e-10, 1.3854e-10, 1.381128e-10, 1.386424e-10, 
    1.383721e-10, 1.388352e-10, 1.384184e-10, 1.391404e-10, 1.392975e-10, 
    1.391901e-10, 1.396028e-10, 1.383953e-10, 1.38859e-10, 1.353722e-10, 
    1.353927e-10, 1.354882e-10, 1.350682e-10, 1.350425e-10, 1.346577e-10, 
    1.350001e-10, 1.35146e-10, 1.355162e-10, 1.357351e-10, 1.359433e-10, 
    1.364009e-10, 1.369121e-10, 1.376269e-10, 1.381405e-10, 1.384847e-10, 
    1.382736e-10, 1.3846e-10, 1.382517e-10, 1.38154e-10, 1.392386e-10, 
    1.386296e-10, 1.395434e-10, 1.394929e-10, 1.390793e-10, 1.394986e-10, 
    1.354071e-10, 1.352891e-10, 1.348794e-10, 1.352e-10, 1.346158e-10, 
    1.349428e-10, 1.351308e-10, 1.358563e-10, 1.360157e-10, 1.361635e-10, 
    1.364554e-10, 1.368301e-10, 1.374873e-10, 1.380593e-10, 1.385814e-10, 
    1.385431e-10, 1.385566e-10, 1.386732e-10, 1.383843e-10, 1.387207e-10, 
    1.387771e-10, 1.386295e-10, 1.394861e-10, 1.392414e-10, 1.394918e-10, 
    1.393325e-10, 1.353274e-10, 1.35526e-10, 1.354187e-10, 1.356204e-10, 
    1.354783e-10, 1.361103e-10, 1.362998e-10, 1.371866e-10, 1.368227e-10, 
    1.374019e-10, 1.368815e-10, 1.369738e-10, 1.374208e-10, 1.369097e-10, 
    1.380277e-10, 1.372697e-10, 1.386778e-10, 1.379207e-10, 1.387252e-10, 
    1.385791e-10, 1.38821e-10, 1.390376e-10, 1.393102e-10, 1.39813e-10, 
    1.396966e-10, 1.401172e-10, 1.35822e-10, 1.360795e-10, 1.360569e-10, 
    1.363264e-10, 1.365257e-10, 1.369578e-10, 1.376508e-10, 1.373902e-10, 
    1.378687e-10, 1.379647e-10, 1.372378e-10, 1.376841e-10, 1.362519e-10, 
    1.364833e-10, 1.363455e-10, 1.358423e-10, 1.374502e-10, 1.36625e-10, 
    1.38149e-10, 1.377018e-10, 1.390067e-10, 1.383578e-10, 1.396325e-10, 
    1.401774e-10, 1.406904e-10, 1.412898e-10, 1.362201e-10, 1.360451e-10, 
    1.363585e-10, 1.36792e-10, 1.371943e-10, 1.377291e-10, 1.377839e-10, 
    1.378841e-10, 1.381436e-10, 1.383618e-10, 1.379157e-10, 1.384165e-10, 
    1.365369e-10, 1.375219e-10, 1.359789e-10, 1.364435e-10, 1.367664e-10, 
    1.366248e-10, 1.373604e-10, 1.375338e-10, 1.382384e-10, 1.378742e-10, 
    1.400429e-10, 1.390834e-10, 1.417463e-10, 1.41002e-10, 1.35984e-10, 
    1.362195e-10, 1.370393e-10, 1.366492e-10, 1.377648e-10, 1.380394e-10, 
    1.382627e-10, 1.385481e-10, 1.385789e-10, 1.38748e-10, 1.384709e-10, 
    1.38737e-10, 1.377303e-10, 1.381802e-10, 1.369456e-10, 1.372461e-10, 
    1.371079e-10, 1.369562e-10, 1.374242e-10, 1.379227e-10, 1.379334e-10, 
    1.380933e-10, 1.385437e-10, 1.377694e-10, 1.401667e-10, 1.38686e-10, 
    1.364764e-10, 1.3693e-10, 1.369949e-10, 1.368191e-10, 1.380119e-10, 
    1.375797e-10, 1.387439e-10, 1.384292e-10, 1.389448e-10, 1.386886e-10, 
    1.386509e-10, 1.383219e-10, 1.38117e-10, 1.375995e-10, 1.371785e-10, 
    1.368446e-10, 1.369223e-10, 1.37289e-10, 1.379532e-10, 1.385817e-10, 
    1.38444e-10, 1.389056e-10, 1.376839e-10, 1.381962e-10, 1.379982e-10, 
    1.385144e-10, 1.373833e-10, 1.383464e-10, 1.371371e-10, 1.372431e-10, 
    1.375711e-10, 1.382309e-10, 1.383769e-10, 1.385328e-10, 1.384366e-10, 
    1.379701e-10, 1.378937e-10, 1.375632e-10, 1.374719e-10, 1.372201e-10, 
    1.370116e-10, 1.37202e-10, 1.374021e-10, 1.379703e-10, 1.384824e-10, 
    1.390407e-10, 1.391774e-10, 1.398297e-10, 1.392986e-10, 1.401749e-10, 
    1.394298e-10, 1.407197e-10, 1.384023e-10, 1.39408e-10, 1.375861e-10, 
    1.377823e-10, 1.381373e-10, 1.389516e-10, 1.38512e-10, 1.390261e-10, 
    1.378907e-10, 1.373016e-10, 1.371493e-10, 1.368649e-10, 1.371557e-10, 
    1.371321e-10, 1.374104e-10, 1.37321e-10, 1.379892e-10, 1.376302e-10, 
    1.386499e-10, 1.390221e-10, 1.400731e-10, 1.407174e-10, 1.413734e-10, 
    1.416629e-10, 1.417511e-10, 1.417879e-10 ;

 SOIL1N_vr =
  2.497637, 2.49763, 2.497631, 2.497626, 2.497629, 2.497626, 2.497635, 
    2.49763, 2.497633, 2.497636, 2.497616, 2.497626, 2.497606, 2.497612, 
    2.497596, 2.497607, 2.497594, 2.497597, 2.497589, 2.497591, 2.497582, 
    2.497588, 2.497577, 2.497584, 2.497583, 2.497589, 2.497624, 2.497617, 
    2.497624, 2.497623, 2.497624, 2.497629, 2.497632, 2.497637, 2.497636, 
    2.497632, 2.497623, 2.497626, 2.497618, 2.497618, 2.49761, 2.497614, 
    2.497599, 2.497603, 2.497591, 2.497594, 2.497591, 2.497592, 2.497591, 
    2.497596, 2.497594, 2.497598, 2.497613, 2.497608, 2.497622, 2.49763, 
    2.497635, 2.497639, 2.497638, 2.497637, 2.497632, 2.497627, 2.497623, 
    2.497621, 2.497618, 2.497611, 2.497607, 2.497598, 2.4976, 2.497597, 
    2.497595, 2.49759, 2.497591, 2.497589, 2.497597, 2.497592, 2.497601, 
    2.497598, 2.497618, 2.497625, 2.497628, 2.497631, 2.497638, 2.497633, 
    2.497635, 2.497631, 2.497628, 2.497629, 2.497621, 2.497624, 2.497607, 
    2.497614, 2.497595, 2.4976, 2.497594, 2.497597, 2.497592, 2.497596, 
    2.497589, 2.497587, 2.497588, 2.497584, 2.497597, 2.497591, 2.497629, 
    2.497629, 2.497628, 2.497633, 2.497633, 2.497637, 2.497633, 2.497632, 
    2.497628, 2.497625, 2.497623, 2.497618, 2.497613, 2.497605, 2.497599, 
    2.497596, 2.497598, 2.497596, 2.497598, 2.497599, 2.497587, 2.497594, 
    2.497584, 2.497585, 2.497589, 2.497585, 2.497629, 2.49763, 2.497635, 
    2.497631, 2.497638, 2.497634, 2.497632, 2.497624, 2.497622, 2.497621, 
    2.497617, 2.497613, 2.497606, 2.4976, 2.497595, 2.497595, 2.497595, 
    2.497594, 2.497597, 2.497593, 2.497592, 2.497594, 2.497585, 2.497587, 
    2.497585, 2.497586, 2.49763, 2.497628, 2.497629, 2.497627, 2.497628, 
    2.497621, 2.497619, 2.49761, 2.497614, 2.497607, 2.497613, 2.497612, 
    2.497607, 2.497613, 2.497601, 2.497609, 2.497593, 2.497602, 2.497593, 
    2.497595, 2.497592, 2.49759, 2.497587, 2.497581, 2.497582, 2.497578, 
    2.497624, 2.497622, 2.497622, 2.497619, 2.497617, 2.497612, 2.497605, 
    2.497607, 2.497602, 2.497601, 2.497609, 2.497604, 2.49762, 2.497617, 
    2.497619, 2.497624, 2.497607, 2.497616, 2.497599, 2.497604, 2.49759, 
    2.497597, 2.497583, 2.497577, 2.497572, 2.497566, 2.49762, 2.497622, 
    2.497619, 2.497614, 2.49761, 2.497604, 2.497603, 2.497602, 2.497599, 
    2.497597, 2.497602, 2.497596, 2.497617, 2.497606, 2.497623, 2.497618, 
    2.497614, 2.497616, 2.497608, 2.497606, 2.497598, 2.497602, 2.497579, 
    2.497589, 2.497561, 2.497569, 2.497623, 2.49762, 2.497611, 2.497615, 
    2.497603, 2.4976, 2.497598, 2.497595, 2.497595, 2.497593, 2.497596, 
    2.497593, 2.497604, 2.497599, 2.497612, 2.497609, 2.497611, 2.497612, 
    2.497607, 2.497602, 2.497602, 2.4976, 2.497595, 2.497603, 2.497577, 
    2.497593, 2.497617, 2.497612, 2.497612, 2.497614, 2.497601, 2.497605, 
    2.497593, 2.497596, 2.497591, 2.497593, 2.497594, 2.497597, 2.4976, 
    2.497605, 2.49761, 2.497613, 2.497612, 2.497608, 2.497601, 2.497595, 
    2.497596, 2.497591, 2.497604, 2.497599, 2.497601, 2.497595, 2.497607, 
    2.497597, 2.49761, 2.497609, 2.497606, 2.497598, 2.497597, 2.497595, 
    2.497596, 2.497601, 2.497602, 2.497606, 2.497607, 2.497609, 2.497612, 
    2.497609, 2.497607, 2.497601, 2.497596, 2.49759, 2.497588, 2.497581, 
    2.497587, 2.497577, 2.497585, 2.497571, 2.497597, 2.497586, 2.497605, 
    2.497603, 2.497599, 2.497591, 2.497595, 2.49759, 2.497602, 2.497608, 
    2.49761, 2.497613, 2.49761, 2.49761, 2.497607, 2.497608, 2.497601, 
    2.497605, 2.497594, 2.49759, 2.497578, 2.497571, 2.497565, 2.497561, 
    2.497561, 2.49756,
  2.49791, 2.497902, 2.497903, 2.497897, 2.4979, 2.497896, 2.497908, 
    2.497901, 2.497906, 2.497909, 2.497885, 2.497897, 2.497872, 2.49788, 
    2.49786, 2.497873, 2.497858, 2.49786, 2.497851, 2.497854, 2.497843, 
    2.49785, 2.497837, 2.497844, 2.497843, 2.497851, 2.497894, 2.497886, 
    2.497895, 2.497893, 2.497894, 2.4979, 2.497904, 2.49791, 2.497909, 
    2.497904, 2.497893, 2.497897, 2.497887, 2.497887, 2.497877, 2.497881, 
    2.497864, 2.497869, 2.497854, 2.497858, 2.497854, 2.497855, 2.497854, 
    2.497859, 2.497857, 2.497862, 2.49788, 2.497875, 2.497891, 2.497901, 
    2.497908, 2.497912, 2.497912, 2.49791, 2.497904, 2.497898, 2.497894, 
    2.49789, 2.497887, 2.497878, 2.497873, 2.497863, 2.497864, 2.497861, 
    2.497858, 2.497853, 2.497854, 2.497851, 2.497861, 2.497854, 2.497866, 
    2.497863, 2.497887, 2.497896, 2.4979, 2.497903, 2.497911, 2.497905, 
    2.497908, 2.497902, 2.497899, 2.497901, 2.49789, 2.497894, 2.497873, 
    2.497882, 2.497858, 2.497864, 2.497857, 2.497861, 2.497854, 2.49786, 
    2.49785, 2.497848, 2.49785, 2.497844, 2.49786, 2.497854, 2.497901, 
    2.4979, 2.497899, 2.497905, 2.497905, 2.49791, 2.497906, 2.497904, 
    2.497899, 2.497896, 2.497893, 2.497887, 2.49788, 2.497871, 2.497864, 
    2.497859, 2.497862, 2.497859, 2.497862, 2.497864, 2.497849, 2.497857, 
    2.497845, 2.497846, 2.497851, 2.497846, 2.4979, 2.497902, 2.497907, 
    2.497903, 2.497911, 2.497906, 2.497904, 2.497894, 2.497892, 2.49789, 
    2.497886, 2.497881, 2.497872, 2.497865, 2.497858, 2.497858, 2.497858, 
    2.497857, 2.49786, 2.497856, 2.497855, 2.497857, 2.497846, 2.497849, 
    2.497846, 2.497848, 2.497901, 2.497899, 2.4979, 2.497897, 2.497899, 
    2.497891, 2.497888, 2.497876, 2.497881, 2.497874, 2.49788, 2.497879, 
    2.497873, 2.49788, 2.497865, 2.497875, 2.497857, 2.497867, 2.497856, 
    2.497858, 2.497855, 2.497852, 2.497848, 2.497841, 2.497843, 2.497837, 
    2.497895, 2.497891, 2.497892, 2.497888, 2.497885, 2.49788, 2.49787, 
    2.497874, 2.497867, 2.497866, 2.497876, 2.49787, 2.497889, 2.497886, 
    2.497888, 2.497895, 2.497873, 2.497884, 2.497864, 2.497869, 2.497852, 
    2.497861, 2.497844, 2.497837, 2.49783, 2.497822, 2.49789, 2.497892, 
    2.497888, 2.497882, 2.497876, 2.497869, 2.497869, 2.497867, 2.497864, 
    2.497861, 2.497867, 2.49786, 2.497885, 2.497872, 2.497893, 2.497886, 
    2.497882, 2.497884, 2.497874, 2.497872, 2.497862, 2.497867, 2.497838, 
    2.497851, 2.497816, 2.497826, 2.497893, 2.49789, 2.497878, 2.497884, 
    2.497869, 2.497865, 2.497862, 2.497858, 2.497858, 2.497856, 2.497859, 
    2.497856, 2.497869, 2.497863, 2.49788, 2.497876, 2.497878, 2.49788, 
    2.497873, 2.497867, 2.497866, 2.497864, 2.497858, 2.497869, 2.497837, 
    2.497856, 2.497886, 2.49788, 2.497879, 2.497881, 2.497865, 2.497871, 
    2.497856, 2.49786, 2.497853, 2.497856, 2.497857, 2.497861, 2.497864, 
    2.497871, 2.497877, 2.497881, 2.49788, 2.497875, 2.497866, 2.497858, 
    2.49786, 2.497854, 2.49787, 2.497863, 2.497866, 2.497859, 2.497874, 
    2.497861, 2.497877, 2.497876, 2.497871, 2.497863, 2.49786, 2.497859, 
    2.49786, 2.497866, 2.497867, 2.497871, 2.497873, 2.497876, 2.497879, 
    2.497876, 2.497874, 2.497866, 2.497859, 2.497852, 2.49785, 2.497841, 
    2.497848, 2.497837, 2.497847, 2.497829, 2.49786, 2.497847, 2.497871, 
    2.497869, 2.497864, 2.497853, 2.497859, 2.497852, 2.497867, 2.497875, 
    2.497877, 2.497881, 2.497877, 2.497877, 2.497874, 2.497875, 2.497866, 
    2.49787, 2.497857, 2.497852, 2.497838, 2.497829, 2.497821, 2.497817, 
    2.497816, 2.497815,
  2.498032, 2.498024, 2.498025, 2.498018, 2.498022, 2.498017, 2.49803, 
    2.498023, 2.498028, 2.498031, 2.498004, 2.498018, 2.497991, 2.497999, 
    2.497978, 2.497992, 2.497975, 2.497978, 2.497968, 2.497971, 2.497959, 
    2.497967, 2.497952, 2.497961, 2.497959, 2.497967, 2.498015, 2.498006, 
    2.498016, 2.498014, 2.498015, 2.498022, 2.498025, 2.498033, 2.498031, 
    2.498026, 2.498014, 2.498018, 2.498007, 2.498008, 2.497996, 2.498001, 
    2.497982, 2.497987, 2.497971, 2.497975, 2.497971, 2.497972, 2.497971, 
    2.497977, 2.497975, 2.49798, 2.498, 2.497994, 2.498012, 2.498023, 
    2.49803, 2.498035, 2.498034, 2.498033, 2.498026, 2.498019, 2.498014, 
    2.498011, 2.498008, 2.497998, 2.497992, 2.49798, 2.497983, 2.497979, 
    2.497976, 2.49797, 2.497971, 2.497968, 2.497979, 2.497972, 2.497984, 
    2.497981, 2.498007, 2.498017, 2.498021, 2.498025, 2.498034, 2.498028, 
    2.49803, 2.498024, 2.49802, 2.498022, 2.498011, 2.498015, 2.497992, 
    2.498002, 2.497976, 2.497982, 2.497974, 2.497978, 2.497972, 2.497978, 
    2.497967, 2.497965, 2.497966, 2.49796, 2.497978, 2.497971, 2.498022, 
    2.498022, 2.498021, 2.498027, 2.498027, 2.498033, 2.498028, 2.498026, 
    2.49802, 2.498017, 2.498014, 2.498007, 2.498, 2.497989, 2.497982, 
    2.497977, 2.49798, 2.497977, 2.49798, 2.497982, 2.497966, 2.497975, 
    2.497961, 2.497962, 2.497968, 2.497962, 2.498022, 2.498024, 2.498029, 
    2.498025, 2.498034, 2.498029, 2.498026, 2.498015, 2.498013, 2.498011, 
    2.498006, 2.498001, 2.497991, 2.497983, 2.497975, 2.497976, 2.497976, 
    2.497974, 2.497978, 2.497973, 2.497972, 2.497975, 2.497962, 2.497966, 
    2.497962, 2.497964, 2.498023, 2.49802, 2.498022, 2.498019, 2.498021, 
    2.498012, 2.498009, 2.497996, 2.498001, 2.497993, 2.498, 2.497999, 
    2.497992, 2.498, 2.497983, 2.497994, 2.497974, 2.497985, 2.497973, 
    2.497975, 2.497972, 2.497969, 2.497965, 2.497957, 2.497959, 2.497953, 
    2.498016, 2.498012, 2.498012, 2.498008, 2.498005, 2.497999, 2.497989, 
    2.497993, 2.497986, 2.497984, 2.497995, 2.497988, 2.498009, 2.498006, 
    2.498008, 2.498015, 2.497992, 2.498004, 2.497982, 2.497988, 2.497969, 
    2.497979, 2.49796, 2.497952, 2.497945, 2.497936, 2.49801, 2.498013, 
    2.498008, 2.498002, 2.497996, 2.497988, 2.497987, 2.497986, 2.497982, 
    2.497978, 2.497985, 2.497978, 2.498005, 2.497991, 2.498013, 2.498007, 
    2.498002, 2.498004, 2.497993, 2.497991, 2.49798, 2.497986, 2.497954, 
    2.497968, 2.497929, 2.49794, 2.498013, 2.49801, 2.497998, 2.498003, 
    2.497987, 2.497983, 2.49798, 2.497976, 2.497975, 2.497973, 2.497977, 
    2.497973, 2.497988, 2.497981, 2.497999, 2.497995, 2.497997, 2.497999, 
    2.497992, 2.497985, 2.497985, 2.497983, 2.497976, 2.497987, 2.497952, 
    2.497974, 2.498006, 2.497999, 2.497998, 2.498001, 2.497984, 2.49799, 
    2.497973, 2.497977, 2.49797, 2.497974, 2.497974, 2.497979, 2.497982, 
    2.49799, 2.497996, 2.498001, 2.498, 2.497994, 2.497984, 2.497975, 
    2.497977, 2.497971, 2.497988, 2.497981, 2.497984, 2.497976, 2.497993, 
    2.497979, 2.497996, 2.497995, 2.49799, 2.49798, 2.497978, 2.497976, 
    2.497977, 2.497984, 2.497985, 2.49799, 2.497992, 2.497995, 2.497998, 
    2.497995, 2.497993, 2.497984, 2.497977, 2.497969, 2.497967, 2.497957, 
    2.497965, 2.497952, 2.497963, 2.497944, 2.497978, 2.497963, 2.49799, 
    2.497987, 2.497982, 2.49797, 2.497976, 2.497969, 2.497985, 2.497994, 
    2.497996, 2.498, 2.497996, 2.497997, 2.497993, 2.497994, 2.497984, 
    2.497989, 2.497974, 2.497969, 2.497953, 2.497944, 2.497935, 2.49793, 
    2.497929, 2.497928,
  2.498126, 2.498117, 2.498119, 2.498111, 2.498116, 2.498111, 2.498124, 
    2.498116, 2.498121, 2.498125, 2.498098, 2.498111, 2.498083, 2.498092, 
    2.49807, 2.498085, 2.498067, 2.498071, 2.498061, 2.498064, 2.498051, 
    2.49806, 2.498044, 2.498053, 2.498051, 2.49806, 2.498108, 2.498099, 
    2.498109, 2.498108, 2.498108, 2.498115, 2.498119, 2.498127, 2.498125, 
    2.49812, 2.498107, 2.498111, 2.498101, 2.498101, 2.498089, 2.498094, 
    2.498074, 2.49808, 2.498064, 2.498068, 2.498064, 2.498065, 2.498064, 
    2.49807, 2.498067, 2.498072, 2.498093, 2.498087, 2.498106, 2.498116, 
    2.498124, 2.498129, 2.498128, 2.498127, 2.49812, 2.498113, 2.498108, 
    2.498104, 2.498101, 2.498091, 2.498085, 2.498073, 2.498075, 2.498072, 
    2.498068, 2.498062, 2.498063, 2.49806, 2.498072, 2.498064, 2.498076, 
    2.498073, 2.4981, 2.49811, 2.498115, 2.498118, 2.498128, 2.498121, 
    2.498124, 2.498118, 2.498114, 2.498116, 2.498104, 2.498109, 2.498085, 
    2.498095, 2.498069, 2.498075, 2.498067, 2.498071, 2.498064, 2.49807, 
    2.49806, 2.498057, 2.498059, 2.498053, 2.498071, 2.498064, 2.498116, 
    2.498116, 2.498114, 2.49812, 2.498121, 2.498127, 2.498122, 2.498119, 
    2.498114, 2.498111, 2.498107, 2.498101, 2.498093, 2.498082, 2.498075, 
    2.498069, 2.498072, 2.49807, 2.498073, 2.498074, 2.498058, 2.498067, 
    2.498054, 2.498054, 2.49806, 2.498054, 2.498115, 2.498117, 2.498123, 
    2.498118, 2.498127, 2.498122, 2.49812, 2.498109, 2.498106, 2.498104, 
    2.4981, 2.498094, 2.498084, 2.498076, 2.498068, 2.498068, 2.498068, 
    2.498066, 2.498071, 2.498066, 2.498065, 2.498067, 2.498054, 2.498058, 
    2.498054, 2.498057, 2.498116, 2.498114, 2.498115, 2.498112, 2.498114, 
    2.498105, 2.498102, 2.498089, 2.498094, 2.498085, 2.498093, 2.498092, 
    2.498085, 2.498093, 2.498076, 2.498087, 2.498066, 2.498078, 2.498066, 
    2.498068, 2.498064, 2.498061, 2.498057, 2.498049, 2.498051, 2.498045, 
    2.498109, 2.498105, 2.498106, 2.498101, 2.498099, 2.498092, 2.498082, 
    2.498086, 2.498079, 2.498077, 2.498088, 2.498081, 2.498103, 2.498099, 
    2.498101, 2.498109, 2.498085, 2.498097, 2.498074, 2.498081, 2.498061, 
    2.498071, 2.498052, 2.498044, 2.498036, 2.498027, 2.498103, 2.498106, 
    2.498101, 2.498095, 2.498089, 2.49808, 2.49808, 2.498078, 2.498074, 
    2.498071, 2.498078, 2.49807, 2.498098, 2.498084, 2.498107, 2.4981, 
    2.498095, 2.498097, 2.498086, 2.498084, 2.498073, 2.498078, 2.498046, 
    2.49806, 2.498021, 2.498032, 2.498107, 2.498103, 2.498091, 2.498097, 
    2.49808, 2.498076, 2.498073, 2.498068, 2.498068, 2.498065, 2.49807, 
    2.498065, 2.49808, 2.498074, 2.498092, 2.498088, 2.49809, 2.498092, 
    2.498085, 2.498078, 2.498078, 2.498075, 2.498068, 2.49808, 2.498044, 
    2.498066, 2.498099, 2.498093, 2.498091, 2.498094, 2.498076, 2.498083, 
    2.498065, 2.49807, 2.498062, 2.498066, 2.498067, 2.498072, 2.498075, 
    2.498083, 2.498089, 2.498094, 2.498093, 2.498087, 2.498077, 2.498068, 
    2.49807, 2.498063, 2.498081, 2.498074, 2.498077, 2.498069, 2.498086, 
    2.498071, 2.49809, 2.498088, 2.498083, 2.498073, 2.498071, 2.498069, 
    2.49807, 2.498077, 2.498078, 2.498083, 2.498085, 2.498088, 2.498091, 
    2.498088, 2.498085, 2.498077, 2.498069, 2.498061, 2.498059, 2.498049, 
    2.498057, 2.498044, 2.498055, 2.498036, 2.49807, 2.498055, 2.498083, 
    2.49808, 2.498075, 2.498062, 2.498069, 2.498061, 2.498078, 2.498087, 
    2.498089, 2.498094, 2.498089, 2.49809, 2.498085, 2.498087, 2.498077, 
    2.498082, 2.498067, 2.498061, 2.498045, 2.498036, 2.498026, 2.498022, 
    2.49802, 2.49802,
  2.498261, 2.498253, 2.498254, 2.498248, 2.498251, 2.498247, 2.498259, 
    2.498252, 2.498256, 2.49826, 2.498235, 2.498247, 2.498222, 2.49823, 
    2.49821, 2.498223, 2.498207, 2.49821, 2.498201, 2.498204, 2.498192, 
    2.4982, 2.498186, 2.498194, 2.498193, 2.4982, 2.498245, 2.498236, 
    2.498245, 2.498244, 2.498245, 2.498251, 2.498254, 2.498261, 2.49826, 
    2.498255, 2.498244, 2.498247, 2.498238, 2.498238, 2.498227, 2.498232, 
    2.498214, 2.498219, 2.498204, 2.498208, 2.498204, 2.498205, 2.498204, 
    2.498209, 2.498207, 2.498212, 2.498231, 2.498225, 2.498242, 2.498252, 
    2.498259, 2.498263, 2.498263, 2.498261, 2.498255, 2.498249, 2.498244, 
    2.498241, 2.498238, 2.498229, 2.498224, 2.498213, 2.498214, 2.498211, 
    2.498208, 2.498202, 2.498203, 2.498201, 2.498211, 2.498204, 2.498216, 
    2.498213, 2.498237, 2.498246, 2.49825, 2.498254, 2.498262, 2.498256, 
    2.498259, 2.498253, 2.49825, 2.498251, 2.498241, 2.498245, 2.498223, 
    2.498233, 2.498208, 2.498214, 2.498207, 2.49821, 2.498204, 2.49821, 
    2.4982, 2.498198, 2.498199, 2.498194, 2.49821, 2.498204, 2.498251, 
    2.498251, 2.49825, 2.498256, 2.498256, 2.498261, 2.498257, 2.498255, 
    2.49825, 2.498247, 2.498244, 2.498238, 2.49823, 2.498221, 2.498214, 
    2.498209, 2.498212, 2.498209, 2.498212, 2.498214, 2.498199, 2.498207, 
    2.498194, 2.498195, 2.498201, 2.498195, 2.498251, 2.498253, 2.498258, 
    2.498254, 2.498262, 2.498257, 2.498255, 2.498245, 2.498243, 2.498241, 
    2.498237, 2.498232, 2.498223, 2.498215, 2.498208, 2.498208, 2.498208, 
    2.498206, 2.49821, 2.498206, 2.498205, 2.498207, 2.498195, 2.498199, 
    2.498195, 2.498197, 2.498252, 2.49825, 2.498251, 2.498248, 2.49825, 
    2.498241, 2.498239, 2.498227, 2.498232, 2.498224, 2.498231, 2.49823, 
    2.498224, 2.49823, 2.498215, 2.498226, 2.498206, 2.498217, 2.498206, 
    2.498208, 2.498204, 2.498201, 2.498198, 2.498191, 2.498192, 2.498187, 
    2.498245, 2.498242, 2.498242, 2.498239, 2.498236, 2.49823, 2.49822, 
    2.498224, 2.498217, 2.498216, 2.498226, 2.49822, 2.49824, 2.498236, 
    2.498238, 2.498245, 2.498223, 2.498235, 2.498214, 2.49822, 2.498202, 
    2.498211, 2.498193, 2.498186, 2.498179, 2.498171, 2.49824, 2.498242, 
    2.498238, 2.498232, 2.498227, 2.498219, 2.498219, 2.498217, 2.498214, 
    2.498211, 2.498217, 2.49821, 2.498236, 2.498222, 2.498243, 2.498237, 
    2.498233, 2.498235, 2.498224, 2.498222, 2.498212, 2.498217, 2.498188, 
    2.498201, 2.498164, 2.498174, 2.498243, 2.49824, 2.498229, 2.498234, 
    2.498219, 2.498215, 2.498212, 2.498208, 2.498208, 2.498205, 2.498209, 
    2.498205, 2.498219, 2.498213, 2.49823, 2.498226, 2.498228, 2.49823, 
    2.498224, 2.498217, 2.498217, 2.498214, 2.498208, 2.498219, 2.498186, 
    2.498206, 2.498236, 2.49823, 2.498229, 2.498232, 2.498215, 2.498221, 
    2.498205, 2.49821, 2.498203, 2.498206, 2.498207, 2.498211, 2.498214, 
    2.498221, 2.498227, 2.498231, 2.49823, 2.498225, 2.498216, 2.498208, 
    2.498209, 2.498203, 2.49822, 2.498213, 2.498216, 2.498209, 2.498224, 
    2.498211, 2.498227, 2.498226, 2.498221, 2.498213, 2.49821, 2.498208, 
    2.49821, 2.498216, 2.498217, 2.498222, 2.498223, 2.498226, 2.498229, 
    2.498227, 2.498224, 2.498216, 2.498209, 2.498201, 2.498199, 2.498191, 
    2.498198, 2.498186, 2.498196, 2.498178, 2.49821, 2.498196, 2.498221, 
    2.498219, 2.498214, 2.498203, 2.498209, 2.498202, 2.498217, 2.498225, 
    2.498227, 2.498231, 2.498227, 2.498228, 2.498224, 2.498225, 2.498216, 
    2.498221, 2.498207, 2.498202, 2.498187, 2.498178, 2.498169, 2.498165, 
    2.498164, 2.498164,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  5.98301e-08, 6.00939e-08, 6.004262e-08, 6.02554e-08, 6.013737e-08, 
    6.02767e-08, 5.988359e-08, 6.010438e-08, 5.996343e-08, 5.985386e-08, 
    6.066833e-08, 6.02649e-08, 6.108748e-08, 6.083015e-08, 6.147663e-08, 
    6.104744e-08, 6.156317e-08, 6.146426e-08, 6.176201e-08, 6.167671e-08, 
    6.205753e-08, 6.180138e-08, 6.225498e-08, 6.199637e-08, 6.203682e-08, 
    6.179292e-08, 6.03461e-08, 6.06181e-08, 6.032997e-08, 6.036876e-08, 
    6.035136e-08, 6.01398e-08, 6.003319e-08, 5.980995e-08, 5.985048e-08, 
    6.001445e-08, 6.038621e-08, 6.026001e-08, 6.057807e-08, 6.057089e-08, 
    6.0925e-08, 6.076534e-08, 6.136055e-08, 6.119138e-08, 6.168027e-08, 
    6.155731e-08, 6.167449e-08, 6.163896e-08, 6.167495e-08, 6.149462e-08, 
    6.157188e-08, 6.141321e-08, 6.079524e-08, 6.097684e-08, 6.043521e-08, 
    6.010954e-08, 5.989327e-08, 5.97398e-08, 5.97615e-08, 5.980285e-08, 
    6.001541e-08, 6.021527e-08, 6.036758e-08, 6.046947e-08, 6.056986e-08, 
    6.087372e-08, 6.103458e-08, 6.139475e-08, 6.132976e-08, 6.143987e-08, 
    6.154508e-08, 6.17217e-08, 6.169263e-08, 6.177045e-08, 6.143697e-08, 
    6.16586e-08, 6.129274e-08, 6.13928e-08, 6.059711e-08, 6.029406e-08, 
    6.016522e-08, 6.005248e-08, 5.977817e-08, 5.99676e-08, 5.989293e-08, 
    6.007059e-08, 6.018348e-08, 6.012765e-08, 6.047225e-08, 6.033828e-08, 
    6.104411e-08, 6.074007e-08, 6.153281e-08, 6.13431e-08, 6.157828e-08, 
    6.145827e-08, 6.166389e-08, 6.147884e-08, 6.179941e-08, 6.186922e-08, 
    6.182151e-08, 6.200477e-08, 6.146858e-08, 6.167448e-08, 6.012608e-08, 
    6.013519e-08, 6.017761e-08, 5.999112e-08, 5.997972e-08, 5.980883e-08, 
    5.996089e-08, 6.002564e-08, 6.019003e-08, 6.028726e-08, 6.037969e-08, 
    6.058293e-08, 6.080991e-08, 6.112733e-08, 6.13554e-08, 6.150827e-08, 
    6.141454e-08, 6.14973e-08, 6.140478e-08, 6.136142e-08, 6.184305e-08, 
    6.15726e-08, 6.197841e-08, 6.195595e-08, 6.17723e-08, 6.195848e-08, 
    6.014158e-08, 6.008919e-08, 5.990725e-08, 6.004963e-08, 5.979022e-08, 
    5.993542e-08, 6.001891e-08, 6.034107e-08, 6.041186e-08, 6.04775e-08, 
    6.060714e-08, 6.077351e-08, 6.106537e-08, 6.131934e-08, 6.15512e-08, 
    6.153422e-08, 6.154019e-08, 6.159198e-08, 6.146369e-08, 6.161305e-08, 
    6.163811e-08, 6.157257e-08, 6.195295e-08, 6.184428e-08, 6.195548e-08, 
    6.188472e-08, 6.010622e-08, 6.019439e-08, 6.014675e-08, 6.023634e-08, 
    6.017321e-08, 6.045389e-08, 6.053804e-08, 6.093184e-08, 6.077023e-08, 
    6.102744e-08, 6.079636e-08, 6.08373e-08, 6.103582e-08, 6.080885e-08, 
    6.130533e-08, 6.096871e-08, 6.1594e-08, 6.125781e-08, 6.161507e-08, 
    6.15502e-08, 6.16576e-08, 6.175379e-08, 6.187481e-08, 6.209811e-08, 
    6.204641e-08, 6.223316e-08, 6.032585e-08, 6.044021e-08, 6.043015e-08, 
    6.054984e-08, 6.063836e-08, 6.083022e-08, 6.113797e-08, 6.102225e-08, 
    6.123471e-08, 6.127735e-08, 6.095458e-08, 6.115275e-08, 6.051675e-08, 
    6.061949e-08, 6.055833e-08, 6.033486e-08, 6.10489e-08, 6.068244e-08, 
    6.135917e-08, 6.116063e-08, 6.174007e-08, 6.145189e-08, 6.201794e-08, 
    6.225992e-08, 6.248771e-08, 6.275387e-08, 6.050263e-08, 6.042492e-08, 
    6.056407e-08, 6.075658e-08, 6.093524e-08, 6.117273e-08, 6.119704e-08, 
    6.124154e-08, 6.135679e-08, 6.14537e-08, 6.12556e-08, 6.1478e-08, 
    6.064331e-08, 6.108071e-08, 6.039554e-08, 6.060183e-08, 6.074524e-08, 
    6.068234e-08, 6.100902e-08, 6.108602e-08, 6.13989e-08, 6.123716e-08, 
    6.220019e-08, 6.17741e-08, 6.295657e-08, 6.262609e-08, 6.039777e-08, 
    6.050237e-08, 6.086641e-08, 6.06932e-08, 6.118859e-08, 6.131054e-08, 
    6.140968e-08, 6.15364e-08, 6.155009e-08, 6.162517e-08, 6.150213e-08, 
    6.162032e-08, 6.117324e-08, 6.137303e-08, 6.082481e-08, 6.095823e-08, 
    6.089685e-08, 6.082953e-08, 6.103733e-08, 6.125871e-08, 6.126346e-08, 
    6.133444e-08, 6.153446e-08, 6.11906e-08, 6.225516e-08, 6.159767e-08, 
    6.061643e-08, 6.08179e-08, 6.084669e-08, 6.076864e-08, 6.129832e-08, 
    6.110638e-08, 6.162335e-08, 6.148363e-08, 6.171256e-08, 6.15988e-08, 
    6.158206e-08, 6.143595e-08, 6.134499e-08, 6.111519e-08, 6.092822e-08, 
    6.077996e-08, 6.081444e-08, 6.097729e-08, 6.127226e-08, 6.155133e-08, 
    6.149019e-08, 6.169516e-08, 6.115268e-08, 6.138013e-08, 6.129222e-08, 
    6.152147e-08, 6.101917e-08, 6.144686e-08, 6.090985e-08, 6.095693e-08, 
    6.110258e-08, 6.139555e-08, 6.14604e-08, 6.15296e-08, 6.14869e-08, 
    6.127975e-08, 6.124581e-08, 6.109904e-08, 6.105851e-08, 6.094668e-08, 
    6.085409e-08, 6.093868e-08, 6.102752e-08, 6.127984e-08, 6.150723e-08, 
    6.175516e-08, 6.181584e-08, 6.210551e-08, 6.186968e-08, 6.225882e-08, 
    6.192796e-08, 6.250072e-08, 6.147167e-08, 6.191825e-08, 6.110921e-08, 
    6.119637e-08, 6.1354e-08, 6.171559e-08, 6.152039e-08, 6.174868e-08, 
    6.124449e-08, 6.09829e-08, 6.091524e-08, 6.078897e-08, 6.091813e-08, 
    6.090762e-08, 6.103121e-08, 6.09915e-08, 6.128822e-08, 6.112883e-08, 
    6.158164e-08, 6.174688e-08, 6.221359e-08, 6.249969e-08, 6.279098e-08, 
    6.291957e-08, 6.295871e-08, 6.297508e-08 ;

 SOIL1_HR_S3 =
  7.100462e-10, 7.131781e-10, 7.125693e-10, 7.150954e-10, 7.136942e-10, 
    7.153482e-10, 7.106812e-10, 7.133024e-10, 7.116291e-10, 7.103282e-10, 
    7.199978e-10, 7.152081e-10, 7.249742e-10, 7.219191e-10, 7.295943e-10, 
    7.244987e-10, 7.306219e-10, 7.294475e-10, 7.329826e-10, 7.319699e-10, 
    7.364914e-10, 7.334501e-10, 7.388357e-10, 7.357652e-10, 7.362455e-10, 
    7.333497e-10, 7.161721e-10, 7.194014e-10, 7.159808e-10, 7.164412e-10, 
    7.162346e-10, 7.13723e-10, 7.124573e-10, 7.098069e-10, 7.102881e-10, 
    7.122348e-10, 7.166483e-10, 7.151502e-10, 7.189263e-10, 7.18841e-10, 
    7.230451e-10, 7.211495e-10, 7.282162e-10, 7.262076e-10, 7.320121e-10, 
    7.305523e-10, 7.319435e-10, 7.315217e-10, 7.31949e-10, 7.29808e-10, 
    7.307253e-10, 7.288414e-10, 7.215045e-10, 7.236606e-10, 7.172301e-10, 
    7.133637e-10, 7.107961e-10, 7.089741e-10, 7.092317e-10, 7.097227e-10, 
    7.122462e-10, 7.14619e-10, 7.164273e-10, 7.176368e-10, 7.188287e-10, 
    7.224362e-10, 7.24346e-10, 7.286223e-10, 7.278507e-10, 7.29158e-10, 
    7.304071e-10, 7.325041e-10, 7.321589e-10, 7.330828e-10, 7.291236e-10, 
    7.317548e-10, 7.274111e-10, 7.285991e-10, 7.191522e-10, 7.155544e-10, 
    7.140247e-10, 7.126863e-10, 7.094297e-10, 7.116786e-10, 7.10792e-10, 
    7.129013e-10, 7.142416e-10, 7.135787e-10, 7.176699e-10, 7.160793e-10, 
    7.244592e-10, 7.208495e-10, 7.302614e-10, 7.28009e-10, 7.308013e-10, 
    7.293765e-10, 7.318177e-10, 7.296206e-10, 7.334268e-10, 7.342555e-10, 
    7.336892e-10, 7.358649e-10, 7.294988e-10, 7.319435e-10, 7.135601e-10, 
    7.136682e-10, 7.141719e-10, 7.119579e-10, 7.118224e-10, 7.097937e-10, 
    7.115989e-10, 7.123676e-10, 7.143193e-10, 7.154736e-10, 7.16571e-10, 
    7.189839e-10, 7.216787e-10, 7.254473e-10, 7.28155e-10, 7.299701e-10, 
    7.288572e-10, 7.298397e-10, 7.287413e-10, 7.282265e-10, 7.339449e-10, 
    7.307339e-10, 7.35552e-10, 7.352854e-10, 7.331048e-10, 7.353154e-10, 
    7.137441e-10, 7.131221e-10, 7.109621e-10, 7.126524e-10, 7.095728e-10, 
    7.112965e-10, 7.122877e-10, 7.161124e-10, 7.169529e-10, 7.177322e-10, 
    7.192713e-10, 7.212465e-10, 7.247117e-10, 7.277269e-10, 7.304797e-10, 
    7.302781e-10, 7.303491e-10, 7.30964e-10, 7.294407e-10, 7.312141e-10, 
    7.315116e-10, 7.307335e-10, 7.352496e-10, 7.339594e-10, 7.352797e-10, 
    7.344396e-10, 7.133243e-10, 7.143711e-10, 7.138054e-10, 7.148691e-10, 
    7.141197e-10, 7.174518e-10, 7.184509e-10, 7.231263e-10, 7.212076e-10, 
    7.242614e-10, 7.215178e-10, 7.220039e-10, 7.243608e-10, 7.216661e-10, 
    7.275606e-10, 7.23564e-10, 7.309879e-10, 7.269965e-10, 7.31238e-10, 
    7.304679e-10, 7.317431e-10, 7.328851e-10, 7.34322e-10, 7.369732e-10, 
    7.363593e-10, 7.385766e-10, 7.159317e-10, 7.172895e-10, 7.1717e-10, 
    7.18591e-10, 7.196419e-10, 7.219199e-10, 7.255736e-10, 7.241996e-10, 
    7.267221e-10, 7.272285e-10, 7.233963e-10, 7.257491e-10, 7.181982e-10, 
    7.19418e-10, 7.186918e-10, 7.160387e-10, 7.245161e-10, 7.201653e-10, 
    7.281998e-10, 7.258426e-10, 7.327223e-10, 7.293007e-10, 7.360214e-10, 
    7.388944e-10, 7.415989e-10, 7.447592e-10, 7.180306e-10, 7.17108e-10, 
    7.1876e-10, 7.210456e-10, 7.231666e-10, 7.259863e-10, 7.262749e-10, 
    7.268032e-10, 7.281716e-10, 7.293222e-10, 7.269701e-10, 7.296106e-10, 
    7.197007e-10, 7.248938e-10, 7.167591e-10, 7.192084e-10, 7.209109e-10, 
    7.201642e-10, 7.240427e-10, 7.249568e-10, 7.286716e-10, 7.267513e-10, 
    7.381852e-10, 7.331262e-10, 7.471659e-10, 7.43242e-10, 7.167856e-10, 
    7.180274e-10, 7.223495e-10, 7.20293e-10, 7.261747e-10, 7.276225e-10, 
    7.287995e-10, 7.303041e-10, 7.304666e-10, 7.31358e-10, 7.298972e-10, 
    7.313004e-10, 7.259924e-10, 7.283644e-10, 7.218556e-10, 7.234396e-10, 
    7.227109e-10, 7.219116e-10, 7.243787e-10, 7.270071e-10, 7.270634e-10, 
    7.279062e-10, 7.30281e-10, 7.261985e-10, 7.388379e-10, 7.310315e-10, 
    7.193816e-10, 7.217735e-10, 7.221153e-10, 7.211887e-10, 7.274773e-10, 
    7.251986e-10, 7.313363e-10, 7.296775e-10, 7.323955e-10, 7.310449e-10, 
    7.308462e-10, 7.291115e-10, 7.280315e-10, 7.253031e-10, 7.230833e-10, 
    7.213232e-10, 7.217324e-10, 7.236659e-10, 7.271679e-10, 7.304812e-10, 
    7.297554e-10, 7.32189e-10, 7.257482e-10, 7.284487e-10, 7.274049e-10, 
    7.301267e-10, 7.241631e-10, 7.292409e-10, 7.228652e-10, 7.234242e-10, 
    7.251534e-10, 7.286318e-10, 7.294017e-10, 7.302233e-10, 7.297163e-10, 
    7.272569e-10, 7.26854e-10, 7.251114e-10, 7.246302e-10, 7.233025e-10, 
    7.222032e-10, 7.232075e-10, 7.242623e-10, 7.27258e-10, 7.299577e-10, 
    7.329013e-10, 7.336218e-10, 7.37061e-10, 7.342611e-10, 7.388813e-10, 
    7.34953e-10, 7.417535e-10, 7.295355e-10, 7.348377e-10, 7.252322e-10, 
    7.262669e-10, 7.281385e-10, 7.324315e-10, 7.30114e-10, 7.328244e-10, 
    7.268382e-10, 7.237325e-10, 7.229292e-10, 7.214301e-10, 7.229635e-10, 
    7.228387e-10, 7.243061e-10, 7.238345e-10, 7.273575e-10, 7.254651e-10, 
    7.308411e-10, 7.32803e-10, 7.383442e-10, 7.417413e-10, 7.451998e-10, 
    7.467267e-10, 7.471914e-10, 7.473857e-10 ;

 SOIL2C =
  5.783957, 5.783963, 5.783962, 5.783967, 5.783964, 5.783967, 5.783958, 
    5.783963, 5.78396, 5.783957, 5.783976, 5.783967, 5.783985, 5.783979, 
    5.783994, 5.783985, 5.783996, 5.783994, 5.784001, 5.783999, 5.784008, 
    5.784002, 5.784012, 5.784006, 5.784007, 5.784001, 5.783968, 5.783975, 
    5.783968, 5.783969, 5.783968, 5.783964, 5.783961, 5.783956, 5.783957, 
    5.783961, 5.783969, 5.783967, 5.783974, 5.783974, 5.783982, 5.783978, 
    5.783992, 5.783988, 5.783999, 5.783996, 5.783999, 5.783998, 5.783999, 
    5.783995, 5.783997, 5.783993, 5.783979, 5.783983, 5.78397, 5.783963, 
    5.783958, 5.783955, 5.783955, 5.783956, 5.783961, 5.783966, 5.783969, 
    5.783971, 5.783974, 5.78398, 5.783984, 5.783992, 5.783991, 5.783993, 
    5.783996, 5.784, 5.783999, 5.784001, 5.783993, 5.783998, 5.78399, 
    5.783992, 5.783974, 5.783967, 5.783964, 5.783962, 5.783956, 5.78396, 
    5.783958, 5.783962, 5.783965, 5.783964, 5.783971, 5.783968, 5.783984, 
    5.783978, 5.783996, 5.783991, 5.783997, 5.783994, 5.783998, 5.783994, 
    5.784002, 5.784003, 5.784002, 5.784006, 5.783994, 5.783999, 5.783964, 
    5.783964, 5.783965, 5.78396, 5.78396, 5.783956, 5.78396, 5.783961, 
    5.783965, 5.783967, 5.783969, 5.783974, 5.783979, 5.783986, 5.783991, 
    5.783995, 5.783993, 5.783995, 5.783993, 5.783992, 5.784003, 5.783997, 
    5.784006, 5.784005, 5.784001, 5.784005, 5.783964, 5.783963, 5.783958, 
    5.783962, 5.783956, 5.783959, 5.783961, 5.783968, 5.78397, 5.783971, 
    5.783975, 5.783978, 5.783985, 5.783991, 5.783996, 5.783996, 5.783996, 
    5.783997, 5.783994, 5.783998, 5.783998, 5.783997, 5.784005, 5.784003, 
    5.784005, 5.784004, 5.783963, 5.783965, 5.783964, 5.783966, 5.783965, 
    5.783971, 5.783973, 5.783982, 5.783978, 5.783984, 5.783979, 5.78398, 
    5.783984, 5.783979, 5.78399, 5.783983, 5.783997, 5.783989, 5.783998, 
    5.783996, 5.783998, 5.784, 5.784003, 5.784009, 5.784007, 5.784011, 
    5.783968, 5.783971, 5.78397, 5.783973, 5.783975, 5.783979, 5.783987, 
    5.783984, 5.783989, 5.78399, 5.783982, 5.783987, 5.783972, 5.783975, 
    5.783973, 5.783968, 5.783985, 5.783976, 5.783991, 5.783987, 5.784, 
    5.783994, 5.784007, 5.784012, 5.784017, 5.784023, 5.783972, 5.78397, 
    5.783973, 5.783978, 5.783982, 5.783988, 5.783988, 5.783989, 5.783991, 
    5.783994, 5.783989, 5.783994, 5.783975, 5.783985, 5.783969, 5.783974, 
    5.783978, 5.783976, 5.783984, 5.783985, 5.783992, 5.783989, 5.784011, 
    5.784001, 5.784028, 5.78402, 5.78397, 5.783972, 5.78398, 5.783977, 
    5.783988, 5.78399, 5.783993, 5.783996, 5.783996, 5.783998, 5.783995, 
    5.783998, 5.783988, 5.783992, 5.783979, 5.783982, 5.783981, 5.783979, 
    5.783984, 5.783989, 5.783989, 5.783991, 5.783996, 5.783988, 5.784012, 
    5.783997, 5.783975, 5.783979, 5.78398, 5.783978, 5.78399, 5.783986, 
    5.783998, 5.783994, 5.783999, 5.783997, 5.783997, 5.783993, 5.783991, 
    5.783986, 5.783982, 5.783978, 5.783979, 5.783983, 5.783989, 5.783996, 
    5.783995, 5.783999, 5.783987, 5.783992, 5.78399, 5.783995, 5.783984, 
    5.783994, 5.783981, 5.783982, 5.783986, 5.783992, 5.783994, 5.783996, 
    5.783995, 5.78399, 5.783989, 5.783986, 5.783985, 5.783982, 5.78398, 
    5.783982, 5.783984, 5.78399, 5.783995, 5.784, 5.784002, 5.784009, 
    5.784003, 5.784012, 5.784005, 5.784018, 5.783994, 5.784004, 5.783986, 
    5.783988, 5.783991, 5.784, 5.783995, 5.784, 5.783989, 5.783983, 5.783981, 
    5.783978, 5.783981, 5.783981, 5.783984, 5.783983, 5.78399, 5.783986, 
    5.783997, 5.784, 5.784011, 5.784018, 5.784024, 5.784027, 5.784028, 
    5.784029 ;

 SOIL2C_TO_SOIL1C =
  1.058451e-09, 1.063122e-09, 1.062214e-09, 1.065981e-09, 1.063891e-09, 
    1.066358e-09, 1.059398e-09, 1.063307e-09, 1.060812e-09, 1.058872e-09, 
    1.073291e-09, 1.066149e-09, 1.080712e-09, 1.076156e-09, 1.087601e-09, 
    1.080003e-09, 1.089134e-09, 1.087383e-09, 1.092654e-09, 1.091144e-09, 
    1.097886e-09, 1.093351e-09, 1.101382e-09, 1.096803e-09, 1.097519e-09, 
    1.093201e-09, 1.067586e-09, 1.072402e-09, 1.067301e-09, 1.067988e-09, 
    1.06768e-09, 1.063934e-09, 1.062047e-09, 1.058095e-09, 1.058812e-09, 
    1.061715e-09, 1.068297e-09, 1.066062e-09, 1.071693e-09, 1.071566e-09, 
    1.077835e-09, 1.075009e-09, 1.085546e-09, 1.082551e-09, 1.091207e-09, 
    1.08903e-09, 1.091104e-09, 1.090475e-09, 1.091113e-09, 1.08792e-09, 
    1.089288e-09, 1.086479e-09, 1.075538e-09, 1.078753e-09, 1.069164e-09, 
    1.063398e-09, 1.05957e-09, 1.056853e-09, 1.057237e-09, 1.057969e-09, 
    1.061732e-09, 1.06527e-09, 1.067967e-09, 1.069771e-09, 1.071548e-09, 
    1.076927e-09, 1.079775e-09, 1.086152e-09, 1.085001e-09, 1.086951e-09, 
    1.088813e-09, 1.09194e-09, 1.091426e-09, 1.092803e-09, 1.086899e-09, 
    1.090823e-09, 1.084346e-09, 1.086117e-09, 1.07203e-09, 1.066665e-09, 
    1.064384e-09, 1.062388e-09, 1.057532e-09, 1.060886e-09, 1.059564e-09, 
    1.062709e-09, 1.064708e-09, 1.063719e-09, 1.06982e-09, 1.067448e-09, 
    1.079944e-09, 1.074561e-09, 1.088596e-09, 1.085238e-09, 1.089401e-09, 
    1.087277e-09, 1.090917e-09, 1.087641e-09, 1.093316e-09, 1.094552e-09, 
    1.093707e-09, 1.096952e-09, 1.087459e-09, 1.091104e-09, 1.063691e-09, 
    1.063853e-09, 1.064604e-09, 1.061302e-09, 1.0611e-09, 1.058075e-09, 
    1.060767e-09, 1.061913e-09, 1.064823e-09, 1.066545e-09, 1.068181e-09, 
    1.071779e-09, 1.075798e-09, 1.081418e-09, 1.085455e-09, 1.088162e-09, 
    1.086502e-09, 1.087967e-09, 1.086329e-09, 1.085562e-09, 1.094089e-09, 
    1.089301e-09, 1.096485e-09, 1.096088e-09, 1.092836e-09, 1.096132e-09, 
    1.063966e-09, 1.063038e-09, 1.059817e-09, 1.062338e-09, 1.057745e-09, 
    1.060316e-09, 1.061794e-09, 1.067497e-09, 1.068751e-09, 1.069913e-09, 
    1.072208e-09, 1.075153e-09, 1.080321e-09, 1.084817e-09, 1.088922e-09, 
    1.088621e-09, 1.088727e-09, 1.089644e-09, 1.087372e-09, 1.090017e-09, 
    1.09046e-09, 1.0893e-09, 1.096034e-09, 1.09411e-09, 1.096079e-09, 
    1.094827e-09, 1.06334e-09, 1.064901e-09, 1.064057e-09, 1.065643e-09, 
    1.064526e-09, 1.069495e-09, 1.070985e-09, 1.077957e-09, 1.075095e-09, 
    1.079649e-09, 1.075558e-09, 1.076283e-09, 1.079797e-09, 1.075779e-09, 
    1.084569e-09, 1.078609e-09, 1.089679e-09, 1.083728e-09, 1.090052e-09, 
    1.088904e-09, 1.090806e-09, 1.092509e-09, 1.094651e-09, 1.098604e-09, 
    1.097689e-09, 1.100995e-09, 1.067228e-09, 1.069253e-09, 1.069074e-09, 
    1.071193e-09, 1.072761e-09, 1.076157e-09, 1.081606e-09, 1.079557e-09, 
    1.083319e-09, 1.084074e-09, 1.078359e-09, 1.081867e-09, 1.070608e-09, 
    1.072427e-09, 1.071344e-09, 1.067388e-09, 1.080029e-09, 1.073541e-09, 
    1.085522e-09, 1.082007e-09, 1.092266e-09, 1.087164e-09, 1.097185e-09, 
    1.101469e-09, 1.105502e-09, 1.110214e-09, 1.070358e-09, 1.068982e-09, 
    1.071445e-09, 1.074854e-09, 1.078017e-09, 1.082221e-09, 1.082652e-09, 
    1.083439e-09, 1.08548e-09, 1.087196e-09, 1.083688e-09, 1.087626e-09, 
    1.072848e-09, 1.080592e-09, 1.068462e-09, 1.072114e-09, 1.074653e-09, 
    1.073539e-09, 1.079323e-09, 1.080686e-09, 1.086225e-09, 1.083362e-09, 
    1.100412e-09, 1.092868e-09, 1.113803e-09, 1.107952e-09, 1.068501e-09, 
    1.070353e-09, 1.076798e-09, 1.073732e-09, 1.082502e-09, 1.084661e-09, 
    1.086416e-09, 1.08866e-09, 1.088902e-09, 1.090231e-09, 1.088053e-09, 
    1.090145e-09, 1.08223e-09, 1.085767e-09, 1.076062e-09, 1.078424e-09, 
    1.077337e-09, 1.076145e-09, 1.079824e-09, 1.083743e-09, 1.083827e-09, 
    1.085084e-09, 1.088625e-09, 1.082538e-09, 1.101385e-09, 1.089745e-09, 
    1.072372e-09, 1.075939e-09, 1.076449e-09, 1.075067e-09, 1.084445e-09, 
    1.081047e-09, 1.090199e-09, 1.087725e-09, 1.091778e-09, 1.089764e-09, 
    1.089468e-09, 1.086881e-09, 1.085271e-09, 1.081202e-09, 1.077892e-09, 
    1.075268e-09, 1.075878e-09, 1.078761e-09, 1.083983e-09, 1.088924e-09, 
    1.087842e-09, 1.09147e-09, 1.081866e-09, 1.085893e-09, 1.084337e-09, 
    1.088395e-09, 1.079503e-09, 1.087075e-09, 1.077567e-09, 1.078401e-09, 
    1.080979e-09, 1.086166e-09, 1.087314e-09, 1.088539e-09, 1.087783e-09, 
    1.084116e-09, 1.083515e-09, 1.080917e-09, 1.080199e-09, 1.078219e-09, 
    1.07658e-09, 1.078078e-09, 1.07965e-09, 1.084118e-09, 1.088143e-09, 
    1.092533e-09, 1.093607e-09, 1.098735e-09, 1.09456e-09, 1.10145e-09, 
    1.095592e-09, 1.105732e-09, 1.087514e-09, 1.09542e-09, 1.081097e-09, 
    1.08264e-09, 1.085431e-09, 1.091832e-09, 1.088376e-09, 1.092418e-09, 
    1.083492e-09, 1.07886e-09, 1.077663e-09, 1.075427e-09, 1.077714e-09, 
    1.077528e-09, 1.079716e-09, 1.079013e-09, 1.084266e-09, 1.081444e-09, 
    1.089461e-09, 1.092386e-09, 1.100649e-09, 1.105714e-09, 1.110871e-09, 
    1.113148e-09, 1.113841e-09, 1.114131e-09 ;

 SOIL2C_TO_SOIL3C =
  7.560366e-11, 7.593726e-11, 7.587241e-11, 7.614148e-11, 7.599223e-11, 
    7.616841e-11, 7.56713e-11, 7.59505e-11, 7.577227e-11, 7.563371e-11, 
    7.666366e-11, 7.615349e-11, 7.719372e-11, 7.68683e-11, 7.768582e-11, 
    7.714307e-11, 7.779526e-11, 7.767018e-11, 7.804671e-11, 7.793884e-11, 
    7.842043e-11, 7.809649e-11, 7.867012e-11, 7.834308e-11, 7.839423e-11, 
    7.808581e-11, 7.625617e-11, 7.660014e-11, 7.623579e-11, 7.628484e-11, 
    7.626283e-11, 7.599531e-11, 7.586048e-11, 7.557818e-11, 7.562943e-11, 
    7.583678e-11, 7.630689e-11, 7.614732e-11, 7.654953e-11, 7.654045e-11, 
    7.698824e-11, 7.678633e-11, 7.753903e-11, 7.73251e-11, 7.794334e-11, 
    7.778785e-11, 7.793603e-11, 7.78911e-11, 7.793662e-11, 7.770858e-11, 
    7.780628e-11, 7.760563e-11, 7.682414e-11, 7.70538e-11, 7.636886e-11, 
    7.595703e-11, 7.568354e-11, 7.548947e-11, 7.551691e-11, 7.55692e-11, 
    7.5838e-11, 7.609074e-11, 7.628335e-11, 7.641219e-11, 7.653914e-11, 
    7.692338e-11, 7.712681e-11, 7.758228e-11, 7.75001e-11, 7.763934e-11, 
    7.777239e-11, 7.799574e-11, 7.795898e-11, 7.805738e-11, 7.763568e-11, 
    7.791594e-11, 7.745328e-11, 7.757982e-11, 7.657359e-11, 7.619037e-11, 
    7.602744e-11, 7.588487e-11, 7.5538e-11, 7.577754e-11, 7.568311e-11, 
    7.590778e-11, 7.605053e-11, 7.597994e-11, 7.641571e-11, 7.624629e-11, 
    7.713886e-11, 7.675439e-11, 7.775686e-11, 7.751697e-11, 7.781437e-11, 
    7.766261e-11, 7.792263e-11, 7.768862e-11, 7.809401e-11, 7.818228e-11, 
    7.812196e-11, 7.83537e-11, 7.767564e-11, 7.793603e-11, 7.597795e-11, 
    7.598946e-11, 7.604312e-11, 7.580728e-11, 7.579287e-11, 7.557677e-11, 
    7.576905e-11, 7.585094e-11, 7.605882e-11, 7.618177e-11, 7.629866e-11, 
    7.655566e-11, 7.68427e-11, 7.724411e-11, 7.753252e-11, 7.772585e-11, 
    7.76073e-11, 7.771196e-11, 7.759497e-11, 7.754013e-11, 7.81492e-11, 
    7.780719e-11, 7.832037e-11, 7.829198e-11, 7.805972e-11, 7.829518e-11, 
    7.599756e-11, 7.593129e-11, 7.570122e-11, 7.588127e-11, 7.555324e-11, 
    7.573685e-11, 7.584242e-11, 7.624981e-11, 7.633934e-11, 7.642234e-11, 
    7.658628e-11, 7.679667e-11, 7.716576e-11, 7.748692e-11, 7.778013e-11, 
    7.775864e-11, 7.776621e-11, 7.78317e-11, 7.766946e-11, 7.785834e-11, 
    7.789003e-11, 7.780716e-11, 7.828817e-11, 7.815074e-11, 7.829137e-11, 
    7.82019e-11, 7.595283e-11, 7.606433e-11, 7.600408e-11, 7.611738e-11, 
    7.603756e-11, 7.639248e-11, 7.64989e-11, 7.699689e-11, 7.679252e-11, 
    7.711779e-11, 7.682557e-11, 7.687734e-11, 7.712838e-11, 7.684137e-11, 
    7.74692e-11, 7.704352e-11, 7.783425e-11, 7.740911e-11, 7.786089e-11, 
    7.777886e-11, 7.791468e-11, 7.803632e-11, 7.818936e-11, 7.847174e-11, 
    7.840636e-11, 7.864253e-11, 7.623056e-11, 7.637518e-11, 7.636246e-11, 
    7.651382e-11, 7.662575e-11, 7.686839e-11, 7.725756e-11, 7.711122e-11, 
    7.737989e-11, 7.743383e-11, 7.702565e-11, 7.727625e-11, 7.647198e-11, 
    7.660191e-11, 7.652456e-11, 7.624196e-11, 7.714492e-11, 7.66815e-11, 
    7.753728e-11, 7.728621e-11, 7.801897e-11, 7.765454e-11, 7.837036e-11, 
    7.867636e-11, 7.896443e-11, 7.930102e-11, 7.645412e-11, 7.635585e-11, 
    7.653182e-11, 7.677527e-11, 7.700118e-11, 7.730153e-11, 7.733226e-11, 
    7.738853e-11, 7.753428e-11, 7.765683e-11, 7.740631e-11, 7.768755e-11, 
    7.663202e-11, 7.718515e-11, 7.631869e-11, 7.657958e-11, 7.676092e-11, 
    7.668138e-11, 7.70945e-11, 7.719186e-11, 7.758753e-11, 7.7383e-11, 
    7.860083e-11, 7.8062e-11, 7.955735e-11, 7.913942e-11, 7.632152e-11, 
    7.645379e-11, 7.691416e-11, 7.669511e-11, 7.732158e-11, 7.747579e-11, 
    7.760116e-11, 7.776142e-11, 7.777872e-11, 7.787367e-11, 7.771808e-11, 
    7.786753e-11, 7.730216e-11, 7.755481e-11, 7.686154e-11, 7.703026e-11, 
    7.695265e-11, 7.686751e-11, 7.713029e-11, 7.741024e-11, 7.741625e-11, 
    7.750602e-11, 7.775895e-11, 7.732412e-11, 7.867034e-11, 7.78389e-11, 
    7.659803e-11, 7.68528e-11, 7.688921e-11, 7.679051e-11, 7.746033e-11, 
    7.721762e-11, 7.787136e-11, 7.769468e-11, 7.798417e-11, 7.784032e-11, 
    7.781915e-11, 7.763439e-11, 7.751936e-11, 7.722874e-11, 7.699231e-11, 
    7.680483e-11, 7.684842e-11, 7.705436e-11, 7.742738e-11, 7.778028e-11, 
    7.770298e-11, 7.796218e-11, 7.727616e-11, 7.75638e-11, 7.745262e-11, 
    7.774253e-11, 7.710733e-11, 7.764818e-11, 7.696908e-11, 7.702862e-11, 
    7.721281e-11, 7.75833e-11, 7.76653e-11, 7.775282e-11, 7.769881e-11, 
    7.743685e-11, 7.739394e-11, 7.720833e-11, 7.715708e-11, 7.701566e-11, 
    7.689857e-11, 7.700555e-11, 7.711789e-11, 7.743697e-11, 7.772452e-11, 
    7.803805e-11, 7.811479e-11, 7.848109e-11, 7.818288e-11, 7.867498e-11, 
    7.825657e-11, 7.898089e-11, 7.767955e-11, 7.824429e-11, 7.722119e-11, 
    7.733141e-11, 7.753075e-11, 7.7988e-11, 7.774117e-11, 7.802985e-11, 
    7.739226e-11, 7.706146e-11, 7.69759e-11, 7.681623e-11, 7.697955e-11, 
    7.696627e-11, 7.712255e-11, 7.707233e-11, 7.744756e-11, 7.7246e-11, 
    7.781861e-11, 7.802758e-11, 7.861777e-11, 7.897959e-11, 7.934794e-11, 
    7.951056e-11, 7.956006e-11, 7.958075e-11 ;

 SOIL2C_vr =
  20.00591, 20.00593, 20.00593, 20.00594, 20.00593, 20.00594, 20.00592, 
    20.00593, 20.00592, 20.00591, 20.00596, 20.00594, 20.00599, 20.00597, 
    20.00601, 20.00599, 20.00602, 20.00601, 20.00603, 20.00603, 20.00605, 
    20.00603, 20.00606, 20.00604, 20.00605, 20.00603, 20.00594, 20.00596, 
    20.00594, 20.00595, 20.00595, 20.00593, 20.00592, 20.00591, 20.00591, 
    20.00592, 20.00595, 20.00594, 20.00596, 20.00596, 20.00598, 20.00597, 
    20.00601, 20.00599, 20.00603, 20.00602, 20.00603, 20.00602, 20.00603, 
    20.00601, 20.00602, 20.00601, 20.00597, 20.00598, 20.00595, 20.00593, 
    20.00592, 20.00591, 20.00591, 20.00591, 20.00592, 20.00594, 20.00595, 
    20.00595, 20.00596, 20.00598, 20.00599, 20.00601, 20.006, 20.00601, 
    20.00602, 20.00603, 20.00603, 20.00603, 20.00601, 20.00602, 20.006, 
    20.00601, 20.00596, 20.00594, 20.00593, 20.00593, 20.00591, 20.00592, 
    20.00592, 20.00593, 20.00593, 20.00593, 20.00595, 20.00594, 20.00599, 
    20.00597, 20.00602, 20.006, 20.00602, 20.00601, 20.00602, 20.00601, 
    20.00603, 20.00604, 20.00603, 20.00604, 20.00601, 20.00603, 20.00593, 
    20.00593, 20.00593, 20.00592, 20.00592, 20.00591, 20.00592, 20.00592, 
    20.00593, 20.00594, 20.00595, 20.00596, 20.00597, 20.00599, 20.00601, 
    20.00601, 20.00601, 20.00601, 20.00601, 20.00601, 20.00603, 20.00602, 
    20.00604, 20.00604, 20.00603, 20.00604, 20.00593, 20.00593, 20.00592, 
    20.00593, 20.00591, 20.00592, 20.00592, 20.00594, 20.00595, 20.00595, 
    20.00596, 20.00597, 20.00599, 20.006, 20.00602, 20.00602, 20.00602, 
    20.00602, 20.00601, 20.00602, 20.00602, 20.00602, 20.00604, 20.00603, 
    20.00604, 20.00604, 20.00593, 20.00593, 20.00593, 20.00594, 20.00593, 
    20.00595, 20.00595, 20.00598, 20.00597, 20.00599, 20.00597, 20.00597, 
    20.00599, 20.00597, 20.006, 20.00598, 20.00602, 20.006, 20.00602, 
    20.00602, 20.00602, 20.00603, 20.00604, 20.00605, 20.00605, 20.00606, 
    20.00594, 20.00595, 20.00595, 20.00596, 20.00596, 20.00597, 20.00599, 
    20.00599, 20.006, 20.006, 20.00598, 20.00599, 20.00595, 20.00596, 
    20.00596, 20.00594, 20.00599, 20.00596, 20.00601, 20.00599, 20.00603, 
    20.00601, 20.00605, 20.00606, 20.00607, 20.00609, 20.00595, 20.00595, 
    20.00596, 20.00597, 20.00598, 20.00599, 20.006, 20.006, 20.00601, 
    20.00601, 20.006, 20.00601, 20.00596, 20.00599, 20.00595, 20.00596, 
    20.00597, 20.00596, 20.00599, 20.00599, 20.00601, 20.006, 20.00606, 
    20.00603, 20.0061, 20.00608, 20.00595, 20.00595, 20.00598, 20.00596, 
    20.00599, 20.006, 20.00601, 20.00602, 20.00602, 20.00602, 20.00601, 
    20.00602, 20.00599, 20.00601, 20.00597, 20.00598, 20.00598, 20.00597, 
    20.00599, 20.006, 20.006, 20.006, 20.00602, 20.00599, 20.00606, 20.00602, 
    20.00596, 20.00597, 20.00597, 20.00597, 20.006, 20.00599, 20.00602, 
    20.00601, 20.00603, 20.00602, 20.00602, 20.00601, 20.006, 20.00599, 
    20.00598, 20.00597, 20.00597, 20.00598, 20.006, 20.00602, 20.00601, 
    20.00603, 20.00599, 20.00601, 20.006, 20.00602, 20.00599, 20.00601, 
    20.00598, 20.00598, 20.00599, 20.00601, 20.00601, 20.00602, 20.00601, 
    20.006, 20.006, 20.00599, 20.00599, 20.00598, 20.00598, 20.00598, 
    20.00599, 20.006, 20.00601, 20.00603, 20.00603, 20.00605, 20.00604, 
    20.00606, 20.00604, 20.00607, 20.00601, 20.00604, 20.00599, 20.006, 
    20.00601, 20.00603, 20.00602, 20.00603, 20.006, 20.00598, 20.00598, 
    20.00597, 20.00598, 20.00598, 20.00599, 20.00598, 20.006, 20.00599, 
    20.00602, 20.00603, 20.00606, 20.00607, 20.00609, 20.0061, 20.0061, 
    20.0061,
  20.00534, 20.00536, 20.00536, 20.00538, 20.00537, 20.00538, 20.00535, 
    20.00537, 20.00535, 20.00535, 20.00541, 20.00538, 20.00544, 20.00542, 
    20.00547, 20.00544, 20.00548, 20.00547, 20.00549, 20.00549, 20.00552, 
    20.0055, 20.00553, 20.00551, 20.00551, 20.0055, 20.00538, 20.0054, 
    20.00538, 20.00538, 20.00538, 20.00537, 20.00536, 20.00534, 20.00534, 
    20.00536, 20.00539, 20.00538, 20.0054, 20.0054, 20.00543, 20.00541, 
    20.00546, 20.00545, 20.00549, 20.00548, 20.00549, 20.00548, 20.00549, 
    20.00547, 20.00548, 20.00547, 20.00542, 20.00543, 20.00539, 20.00537, 
    20.00535, 20.00534, 20.00534, 20.00534, 20.00536, 20.00537, 20.00538, 
    20.00539, 20.0054, 20.00542, 20.00544, 20.00546, 20.00546, 20.00547, 
    20.00548, 20.00549, 20.00549, 20.00549, 20.00547, 20.00548, 20.00546, 
    20.00546, 20.0054, 20.00538, 20.00537, 20.00536, 20.00534, 20.00535, 
    20.00535, 20.00536, 20.00537, 20.00537, 20.00539, 20.00538, 20.00544, 
    20.00541, 20.00547, 20.00546, 20.00548, 20.00547, 20.00549, 20.00547, 
    20.0055, 20.0055, 20.0055, 20.00551, 20.00547, 20.00549, 20.00537, 
    20.00537, 20.00537, 20.00536, 20.00536, 20.00534, 20.00535, 20.00536, 
    20.00537, 20.00538, 20.00539, 20.0054, 20.00542, 20.00544, 20.00546, 
    20.00547, 20.00547, 20.00547, 20.00546, 20.00546, 20.0055, 20.00548, 
    20.00551, 20.00551, 20.00549, 20.00551, 20.00537, 20.00536, 20.00535, 
    20.00536, 20.00534, 20.00535, 20.00536, 20.00538, 20.00539, 20.00539, 
    20.0054, 20.00542, 20.00544, 20.00546, 20.00548, 20.00547, 20.00548, 
    20.00548, 20.00547, 20.00548, 20.00548, 20.00548, 20.00551, 20.0055, 
    20.00551, 20.0055, 20.00537, 20.00537, 20.00537, 20.00537, 20.00537, 
    20.00539, 20.0054, 20.00543, 20.00542, 20.00544, 20.00542, 20.00542, 
    20.00544, 20.00542, 20.00546, 20.00543, 20.00548, 20.00545, 20.00548, 
    20.00548, 20.00548, 20.00549, 20.0055, 20.00552, 20.00551, 20.00553, 
    20.00538, 20.00539, 20.00539, 20.0054, 20.00541, 20.00542, 20.00545, 
    20.00544, 20.00545, 20.00546, 20.00543, 20.00545, 20.0054, 20.00541, 
    20.0054, 20.00538, 20.00544, 20.00541, 20.00546, 20.00545, 20.00549, 
    20.00547, 20.00551, 20.00553, 20.00555, 20.00557, 20.0054, 20.00539, 
    20.0054, 20.00541, 20.00543, 20.00545, 20.00545, 20.00545, 20.00546, 
    20.00547, 20.00545, 20.00547, 20.00541, 20.00544, 20.00539, 20.0054, 
    20.00541, 20.00541, 20.00543, 20.00544, 20.00546, 20.00545, 20.00553, 
    20.00549, 20.00558, 20.00556, 20.00539, 20.0054, 20.00542, 20.00541, 
    20.00545, 20.00546, 20.00546, 20.00548, 20.00548, 20.00548, 20.00547, 
    20.00548, 20.00545, 20.00546, 20.00542, 20.00543, 20.00543, 20.00542, 
    20.00544, 20.00545, 20.00546, 20.00546, 20.00547, 20.00545, 20.00553, 
    20.00548, 20.0054, 20.00542, 20.00542, 20.00542, 20.00546, 20.00544, 
    20.00548, 20.00547, 20.00549, 20.00548, 20.00548, 20.00547, 20.00546, 
    20.00544, 20.00543, 20.00542, 20.00542, 20.00543, 20.00546, 20.00548, 
    20.00547, 20.00549, 20.00545, 20.00546, 20.00546, 20.00547, 20.00544, 
    20.00547, 20.00543, 20.00543, 20.00544, 20.00546, 20.00547, 20.00547, 
    20.00547, 20.00546, 20.00545, 20.00544, 20.00544, 20.00543, 20.00542, 
    20.00543, 20.00544, 20.00546, 20.00547, 20.00549, 20.0055, 20.00552, 
    20.0055, 20.00553, 20.0055, 20.00555, 20.00547, 20.0055, 20.00544, 
    20.00545, 20.00546, 20.00549, 20.00547, 20.00549, 20.00545, 20.00543, 
    20.00543, 20.00542, 20.00543, 20.00543, 20.00544, 20.00543, 20.00546, 
    20.00544, 20.00548, 20.00549, 20.00553, 20.00555, 20.00557, 20.00558, 
    20.00558, 20.00558,
  20.00503, 20.00505, 20.00505, 20.00507, 20.00506, 20.00507, 20.00504, 
    20.00505, 20.00504, 20.00503, 20.0051, 20.00507, 20.00514, 20.00512, 
    20.00517, 20.00513, 20.00518, 20.00517, 20.00519, 20.00519, 20.00522, 
    20.0052, 20.00524, 20.00521, 20.00522, 20.0052, 20.00507, 20.0051, 
    20.00507, 20.00508, 20.00508, 20.00506, 20.00505, 20.00503, 20.00503, 
    20.00505, 20.00508, 20.00507, 20.00509, 20.00509, 20.00512, 20.00511, 
    20.00516, 20.00515, 20.00519, 20.00518, 20.00519, 20.00518, 20.00519, 
    20.00517, 20.00518, 20.00517, 20.00511, 20.00513, 20.00508, 20.00505, 
    20.00504, 20.00502, 20.00503, 20.00503, 20.00505, 20.00506, 20.00508, 
    20.00508, 20.00509, 20.00512, 20.00513, 20.00516, 20.00516, 20.00517, 
    20.00517, 20.00519, 20.00519, 20.00519, 20.00517, 20.00518, 20.00515, 
    20.00516, 20.0051, 20.00507, 20.00506, 20.00505, 20.00503, 20.00504, 
    20.00504, 20.00505, 20.00506, 20.00506, 20.00508, 20.00507, 20.00513, 
    20.00511, 20.00517, 20.00516, 20.00518, 20.00517, 20.00519, 20.00517, 
    20.0052, 20.0052, 20.0052, 20.00521, 20.00517, 20.00519, 20.00506, 
    20.00506, 20.00506, 20.00504, 20.00504, 20.00503, 20.00504, 20.00505, 
    20.00506, 20.00507, 20.00508, 20.00509, 20.00511, 20.00514, 20.00516, 
    20.00517, 20.00517, 20.00517, 20.00516, 20.00516, 20.0052, 20.00518, 
    20.00521, 20.00521, 20.00519, 20.00521, 20.00506, 20.00505, 20.00504, 
    20.00505, 20.00503, 20.00504, 20.00505, 20.00507, 20.00508, 20.00508, 
    20.0051, 20.00511, 20.00513, 20.00516, 20.00518, 20.00517, 20.00517, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00518, 20.00521, 20.0052, 
    20.00521, 20.0052, 20.00505, 20.00506, 20.00506, 20.00507, 20.00506, 
    20.00508, 20.00509, 20.00512, 20.00511, 20.00513, 20.00511, 20.00512, 
    20.00513, 20.00511, 20.00516, 20.00513, 20.00518, 20.00515, 20.00518, 
    20.00518, 20.00518, 20.00519, 20.0052, 20.00522, 20.00522, 20.00523, 
    20.00507, 20.00508, 20.00508, 20.00509, 20.0051, 20.00512, 20.00514, 
    20.00513, 20.00515, 20.00515, 20.00513, 20.00514, 20.00509, 20.0051, 
    20.00509, 20.00507, 20.00513, 20.0051, 20.00516, 20.00514, 20.00519, 
    20.00517, 20.00521, 20.00524, 20.00525, 20.00528, 20.00509, 20.00508, 
    20.00509, 20.00511, 20.00512, 20.00514, 20.00515, 20.00515, 20.00516, 
    20.00517, 20.00515, 20.00517, 20.0051, 20.00514, 20.00508, 20.0051, 
    20.00511, 20.0051, 20.00513, 20.00514, 20.00516, 20.00515, 20.00523, 
    20.0052, 20.00529, 20.00527, 20.00508, 20.00509, 20.00512, 20.0051, 
    20.00515, 20.00516, 20.00516, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00518, 20.00514, 20.00516, 20.00512, 20.00513, 20.00512, 20.00512, 
    20.00513, 20.00515, 20.00515, 20.00516, 20.00517, 20.00515, 20.00524, 
    20.00518, 20.0051, 20.00511, 20.00512, 20.00511, 20.00516, 20.00514, 
    20.00518, 20.00517, 20.00519, 20.00518, 20.00518, 20.00517, 20.00516, 
    20.00514, 20.00512, 20.00511, 20.00511, 20.00513, 20.00515, 20.00518, 
    20.00517, 20.00519, 20.00514, 20.00516, 20.00515, 20.00517, 20.00513, 
    20.00517, 20.00512, 20.00513, 20.00514, 20.00516, 20.00517, 20.00517, 
    20.00517, 20.00515, 20.00515, 20.00514, 20.00513, 20.00513, 20.00512, 
    20.00513, 20.00513, 20.00515, 20.00517, 20.00519, 20.0052, 20.00522, 
    20.0052, 20.00524, 20.00521, 20.00526, 20.00517, 20.00521, 20.00514, 
    20.00515, 20.00516, 20.00519, 20.00517, 20.00519, 20.00515, 20.00513, 
    20.00512, 20.00511, 20.00512, 20.00512, 20.00513, 20.00513, 20.00515, 
    20.00514, 20.00518, 20.00519, 20.00523, 20.00526, 20.00528, 20.00529, 
    20.00529, 20.00529,
  20.00479, 20.00481, 20.00481, 20.00483, 20.00482, 20.00483, 20.0048, 
    20.00481, 20.0048, 20.00479, 20.00486, 20.00483, 20.0049, 20.00488, 
    20.00493, 20.0049, 20.00494, 20.00493, 20.00496, 20.00495, 20.00498, 
    20.00496, 20.005, 20.00498, 20.00498, 20.00496, 20.00484, 20.00486, 
    20.00484, 20.00484, 20.00484, 20.00482, 20.00481, 20.00479, 20.00479, 
    20.00481, 20.00484, 20.00483, 20.00486, 20.00485, 20.00488, 20.00487, 
    20.00492, 20.00491, 20.00495, 20.00494, 20.00495, 20.00495, 20.00495, 
    20.00493, 20.00494, 20.00493, 20.00488, 20.00489, 20.00484, 20.00482, 
    20.0048, 20.00478, 20.00479, 20.00479, 20.00481, 20.00482, 20.00484, 
    20.00485, 20.00485, 20.00488, 20.00489, 20.00493, 20.00492, 20.00493, 
    20.00494, 20.00495, 20.00495, 20.00496, 20.00493, 20.00495, 20.00492, 
    20.00493, 20.00486, 20.00483, 20.00482, 20.00481, 20.00479, 20.0048, 
    20.0048, 20.00481, 20.00482, 20.00482, 20.00485, 20.00484, 20.0049, 
    20.00487, 20.00494, 20.00492, 20.00494, 20.00493, 20.00495, 20.00493, 
    20.00496, 20.00497, 20.00496, 20.00498, 20.00493, 20.00495, 20.00482, 
    20.00482, 20.00482, 20.0048, 20.0048, 20.00479, 20.0048, 20.00481, 
    20.00482, 20.00483, 20.00484, 20.00486, 20.00488, 20.0049, 20.00492, 
    20.00494, 20.00493, 20.00493, 20.00493, 20.00492, 20.00496, 20.00494, 
    20.00498, 20.00497, 20.00496, 20.00497, 20.00482, 20.00481, 20.0048, 
    20.00481, 20.00479, 20.0048, 20.00481, 20.00484, 20.00484, 20.00485, 
    20.00486, 20.00487, 20.0049, 20.00492, 20.00494, 20.00494, 20.00494, 
    20.00494, 20.00493, 20.00494, 20.00495, 20.00494, 20.00497, 20.00496, 
    20.00497, 20.00497, 20.00481, 20.00482, 20.00482, 20.00483, 20.00482, 
    20.00484, 20.00485, 20.00489, 20.00487, 20.00489, 20.00488, 20.00488, 
    20.00489, 20.00488, 20.00492, 20.00489, 20.00494, 20.00491, 20.00495, 
    20.00494, 20.00495, 20.00496, 20.00497, 20.00499, 20.00498, 20.005, 
    20.00483, 20.00484, 20.00484, 20.00485, 20.00486, 20.00488, 20.0049, 
    20.00489, 20.00491, 20.00492, 20.00489, 20.00491, 20.00485, 20.00486, 
    20.00485, 20.00484, 20.0049, 20.00486, 20.00492, 20.00491, 20.00496, 
    20.00493, 20.00498, 20.005, 20.00502, 20.00504, 20.00485, 20.00484, 
    20.00485, 20.00487, 20.00489, 20.00491, 20.00491, 20.00491, 20.00492, 
    20.00493, 20.00491, 20.00493, 20.00486, 20.0049, 20.00484, 20.00486, 
    20.00487, 20.00486, 20.00489, 20.0049, 20.00493, 20.00491, 20.005, 
    20.00496, 20.00506, 20.00503, 20.00484, 20.00485, 20.00488, 20.00487, 
    20.00491, 20.00492, 20.00493, 20.00494, 20.00494, 20.00495, 20.00493, 
    20.00495, 20.00491, 20.00492, 20.00488, 20.00489, 20.00488, 20.00488, 
    20.00489, 20.00491, 20.00492, 20.00492, 20.00494, 20.00491, 20.005, 
    20.00494, 20.00486, 20.00488, 20.00488, 20.00487, 20.00492, 20.0049, 
    20.00495, 20.00493, 20.00495, 20.00494, 20.00494, 20.00493, 20.00492, 
    20.0049, 20.00489, 20.00487, 20.00488, 20.00489, 20.00492, 20.00494, 
    20.00493, 20.00495, 20.00491, 20.00492, 20.00492, 20.00494, 20.00489, 
    20.00493, 20.00488, 20.00489, 20.0049, 20.00493, 20.00493, 20.00494, 
    20.00493, 20.00492, 20.00491, 20.0049, 20.0049, 20.00489, 20.00488, 
    20.00489, 20.00489, 20.00492, 20.00494, 20.00496, 20.00496, 20.00499, 
    20.00497, 20.005, 20.00497, 20.00502, 20.00493, 20.00497, 20.0049, 
    20.00491, 20.00492, 20.00495, 20.00494, 20.00496, 20.00491, 20.00489, 
    20.00488, 20.00487, 20.00488, 20.00488, 20.00489, 20.00489, 20.00492, 
    20.0049, 20.00494, 20.00496, 20.005, 20.00502, 20.00505, 20.00506, 
    20.00506, 20.00506,
  20.00426, 20.00427, 20.00427, 20.00429, 20.00428, 20.00429, 20.00426, 
    20.00428, 20.00426, 20.00426, 20.00432, 20.00429, 20.00435, 20.00433, 
    20.00438, 20.00435, 20.00438, 20.00438, 20.0044, 20.00439, 20.00442, 
    20.0044, 20.00444, 20.00442, 20.00442, 20.0044, 20.00429, 20.00431, 
    20.00429, 20.0043, 20.00429, 20.00428, 20.00427, 20.00425, 20.00426, 
    20.00427, 20.0043, 20.00429, 20.00431, 20.00431, 20.00434, 20.00433, 
    20.00437, 20.00436, 20.00439, 20.00438, 20.00439, 20.00439, 20.00439, 
    20.00438, 20.00439, 20.00437, 20.00433, 20.00434, 20.0043, 20.00428, 
    20.00426, 20.00425, 20.00425, 20.00425, 20.00427, 20.00428, 20.0043, 
    20.0043, 20.00431, 20.00433, 20.00434, 20.00437, 20.00437, 20.00438, 
    20.00438, 20.0044, 20.00439, 20.0044, 20.00438, 20.00439, 20.00437, 
    20.00437, 20.00431, 20.00429, 20.00428, 20.00427, 20.00425, 20.00426, 
    20.00426, 20.00427, 20.00428, 20.00428, 20.0043, 20.00429, 20.00435, 
    20.00432, 20.00438, 20.00437, 20.00439, 20.00438, 20.00439, 20.00438, 
    20.0044, 20.00441, 20.00441, 20.00442, 20.00438, 20.00439, 20.00428, 
    20.00428, 20.00428, 20.00427, 20.00427, 20.00425, 20.00426, 20.00427, 
    20.00428, 20.00429, 20.0043, 20.00431, 20.00433, 20.00435, 20.00437, 
    20.00438, 20.00437, 20.00438, 20.00437, 20.00437, 20.00441, 20.00439, 
    20.00442, 20.00442, 20.0044, 20.00442, 20.00428, 20.00427, 20.00426, 
    20.00427, 20.00425, 20.00426, 20.00427, 20.00429, 20.0043, 20.0043, 
    20.00431, 20.00433, 20.00435, 20.00437, 20.00438, 20.00438, 20.00438, 
    20.00439, 20.00438, 20.00439, 20.00439, 20.00439, 20.00442, 20.00441, 
    20.00442, 20.00441, 20.00428, 20.00428, 20.00428, 20.00429, 20.00428, 
    20.0043, 20.00431, 20.00434, 20.00433, 20.00434, 20.00433, 20.00433, 
    20.00434, 20.00433, 20.00437, 20.00434, 20.00439, 20.00436, 20.00439, 
    20.00438, 20.00439, 20.0044, 20.00441, 20.00443, 20.00442, 20.00444, 
    20.00429, 20.0043, 20.0043, 20.00431, 20.00432, 20.00433, 20.00435, 
    20.00434, 20.00436, 20.00436, 20.00434, 20.00435, 20.00431, 20.00431, 
    20.00431, 20.00429, 20.00435, 20.00432, 20.00437, 20.00435, 20.0044, 
    20.00438, 20.00442, 20.00444, 20.00446, 20.00447, 20.0043, 20.0043, 
    20.00431, 20.00432, 20.00434, 20.00436, 20.00436, 20.00436, 20.00437, 
    20.00438, 20.00436, 20.00438, 20.00432, 20.00435, 20.0043, 20.00431, 
    20.00432, 20.00432, 20.00434, 20.00435, 20.00437, 20.00436, 20.00443, 
    20.0044, 20.00449, 20.00447, 20.0043, 20.0043, 20.00433, 20.00432, 
    20.00436, 20.00437, 20.00437, 20.00438, 20.00438, 20.00439, 20.00438, 
    20.00439, 20.00436, 20.00437, 20.00433, 20.00434, 20.00434, 20.00433, 
    20.00435, 20.00436, 20.00436, 20.00437, 20.00438, 20.00436, 20.00444, 
    20.00439, 20.00431, 20.00433, 20.00433, 20.00433, 20.00437, 20.00435, 
    20.00439, 20.00438, 20.0044, 20.00439, 20.00439, 20.00438, 20.00437, 
    20.00435, 20.00434, 20.00433, 20.00433, 20.00434, 20.00436, 20.00438, 
    20.00438, 20.0044, 20.00435, 20.00437, 20.00437, 20.00438, 20.00434, 
    20.00438, 20.00434, 20.00434, 20.00435, 20.00437, 20.00438, 20.00438, 
    20.00438, 20.00436, 20.00436, 20.00435, 20.00435, 20.00434, 20.00433, 
    20.00434, 20.00434, 20.00436, 20.00438, 20.0044, 20.0044, 20.00443, 
    20.00441, 20.00444, 20.00441, 20.00446, 20.00438, 20.00441, 20.00435, 
    20.00436, 20.00437, 20.0044, 20.00438, 20.0044, 20.00436, 20.00434, 
    20.00434, 20.00433, 20.00434, 20.00434, 20.00434, 20.00434, 20.00436, 
    20.00435, 20.00439, 20.0044, 20.00443, 20.00446, 20.00448, 20.00449, 
    20.00449, 20.00449,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258142, 0.5258148, 0.5258147, 0.5258151, 0.5258149, 0.5258152, 
    0.5258144, 0.5258148, 0.5258145, 0.5258143, 0.525816, 0.5258151, 
    0.5258169, 0.5258163, 0.5258176, 0.5258168, 0.5258178, 0.5258176, 
    0.5258182, 0.525818, 0.5258189, 0.5258183, 0.5258192, 0.5258187, 
    0.5258188, 0.5258183, 0.5258153, 0.5258159, 0.5258153, 0.5258154, 
    0.5258153, 0.5258149, 0.5258147, 0.5258142, 0.5258143, 0.5258147, 
    0.5258154, 0.5258151, 0.5258158, 0.5258158, 0.5258165, 0.5258162, 
    0.5258174, 0.5258171, 0.5258181, 0.5258178, 0.525818, 0.525818, 0.525818, 
    0.5258177, 0.5258179, 0.5258175, 0.5258163, 0.5258166, 0.5258155, 
    0.5258148, 0.5258144, 0.5258141, 0.5258141, 0.5258142, 0.5258147, 
    0.5258151, 0.5258154, 0.5258155, 0.5258158, 0.5258164, 0.5258167, 
    0.5258175, 0.5258173, 0.5258176, 0.5258178, 0.5258182, 0.5258181, 
    0.5258183, 0.5258176, 0.525818, 0.5258173, 0.5258175, 0.5258158, 
    0.5258152, 0.525815, 0.5258147, 0.5258141, 0.5258145, 0.5258144, 
    0.5258148, 0.525815, 0.5258149, 0.5258156, 0.5258153, 0.5258167, 
    0.5258161, 0.5258178, 0.5258174, 0.5258179, 0.5258176, 0.525818, 
    0.5258176, 0.5258183, 0.5258185, 0.5258183, 0.5258188, 0.5258176, 
    0.525818, 0.5258148, 0.5258149, 0.525815, 0.5258146, 0.5258145, 
    0.5258142, 0.5258145, 0.5258147, 0.525815, 0.5258152, 0.5258154, 
    0.5258158, 0.5258163, 0.5258169, 0.5258174, 0.5258178, 0.5258175, 
    0.5258177, 0.5258175, 0.5258174, 0.5258184, 0.5258179, 0.5258187, 
    0.5258186, 0.5258183, 0.5258186, 0.5258149, 0.5258148, 0.5258144, 
    0.5258147, 0.5258142, 0.5258145, 0.5258147, 0.5258153, 0.5258154, 
    0.5258156, 0.5258158, 0.5258162, 0.5258168, 0.5258173, 0.5258178, 
    0.5258178, 0.5258178, 0.5258179, 0.5258176, 0.5258179, 0.525818, 
    0.5258179, 0.5258186, 0.5258184, 0.5258186, 0.5258185, 0.5258148, 
    0.525815, 0.5258149, 0.5258151, 0.525815, 0.5258155, 0.5258157, 
    0.5258165, 0.5258162, 0.5258167, 0.5258163, 0.5258163, 0.5258167, 
    0.5258163, 0.5258173, 0.5258166, 0.5258179, 0.5258172, 0.5258179, 
    0.5258178, 0.525818, 0.5258182, 0.5258185, 0.5258189, 0.5258188, 
    0.5258192, 0.5258152, 0.5258155, 0.5258155, 0.5258157, 0.5258159, 
    0.5258163, 0.525817, 0.5258167, 0.5258172, 0.5258172, 0.5258166, 
    0.525817, 0.5258157, 0.5258159, 0.5258157, 0.5258153, 0.5258168, 
    0.525816, 0.5258174, 0.525817, 0.5258182, 0.5258176, 0.5258188, 
    0.5258193, 0.5258198, 0.5258203, 0.5258157, 0.5258155, 0.5258158, 
    0.5258161, 0.5258166, 0.525817, 0.5258171, 0.5258172, 0.5258174, 
    0.5258176, 0.5258172, 0.5258176, 0.5258159, 0.5258169, 0.5258154, 
    0.5258158, 0.5258161, 0.525816, 0.5258167, 0.5258169, 0.5258175, 
    0.5258172, 0.5258192, 0.5258183, 0.5258207, 0.52582, 0.5258154, 
    0.5258157, 0.5258164, 0.525816, 0.525817, 0.5258173, 0.5258175, 
    0.5258178, 0.5258178, 0.525818, 0.5258177, 0.5258179, 0.525817, 
    0.5258175, 0.5258163, 0.5258166, 0.5258164, 0.5258163, 0.5258167, 
    0.5258172, 0.5258172, 0.5258173, 0.5258178, 0.525817, 0.5258192, 
    0.5258179, 0.5258159, 0.5258163, 0.5258164, 0.5258162, 0.5258173, 
    0.5258169, 0.525818, 0.5258177, 0.5258182, 0.5258179, 0.5258179, 
    0.5258176, 0.5258174, 0.5258169, 0.5258165, 0.5258162, 0.5258163, 
    0.5258166, 0.5258172, 0.5258178, 0.5258177, 0.5258181, 0.525817, 
    0.5258175, 0.5258173, 0.5258178, 0.5258167, 0.5258176, 0.5258165, 
    0.5258166, 0.5258169, 0.5258175, 0.5258176, 0.5258178, 0.5258177, 
    0.5258173, 0.5258172, 0.5258169, 0.5258168, 0.5258166, 0.5258164, 
    0.5258166, 0.5258167, 0.5258173, 0.5258177, 0.5258182, 0.5258183, 
    0.5258189, 0.5258185, 0.5258193, 0.5258186, 0.5258198, 0.5258176, 
    0.5258186, 0.5258169, 0.5258171, 0.5258174, 0.5258182, 0.5258178, 
    0.5258182, 0.5258172, 0.5258166, 0.5258165, 0.5258163, 0.5258165, 
    0.5258165, 0.5258167, 0.5258167, 0.5258173, 0.5258169, 0.5258179, 
    0.5258182, 0.5258192, 0.5258198, 0.5258204, 0.5258207, 0.5258207, 
    0.5258208 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  1.28498e-20, -2.569961e-21, 0, -1.027984e-20, -7.709882e-21, 2.569961e-21, 
    -1.541976e-20, 1.28498e-20, 0, -7.709882e-21, -1.003089e-36, 
    -2.569961e-21, -1.541976e-20, -1.003089e-36, 1.28498e-20, 1.28498e-20, 
    1.003089e-36, 2.055969e-20, -1.798972e-20, 0, -5.139921e-21, 
    7.709882e-21, -7.709882e-21, -1.003089e-36, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, 2.312965e-20, -2.569961e-21, 2.569961e-21, 0, 2.569961e-21, 
    2.312965e-20, -7.709882e-21, -1.541976e-20, -1.541976e-20, -7.709882e-21, 
    7.709882e-21, -5.139921e-21, -5.139921e-21, 7.709882e-21, -2.569961e-21, 
    1.28498e-20, 1.027984e-20, -1.027984e-20, -1.003089e-36, -1.003089e-36, 
    -5.139921e-21, -1.798972e-20, -1.28498e-20, 1.027984e-20, 1.027984e-20, 
    7.709882e-21, -1.027984e-20, -7.709882e-21, -2.055969e-20, -2.569961e-21, 
    -2.569961e-21, 1.541976e-20, -7.709882e-21, -7.709882e-21, -5.139921e-21, 
    1.28498e-20, 2.569961e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -1.003089e-36, 7.709882e-21, -1.027984e-20, -1.003089e-36, -1.28498e-20, 
    1.798972e-20, -1.027984e-20, -1.003089e-36, -2.569961e-21, -7.709882e-21, 
    1.28498e-20, -7.709882e-21, 1.28498e-20, 7.709882e-21, 2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, 1.003089e-36, -1.027984e-20, 
    -7.709882e-21, -1.28498e-20, -1.28498e-20, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 
    0, 1.28498e-20, -1.027984e-20, 5.139921e-21, -5.139921e-21, 2.055969e-20, 
    -1.027984e-20, -2.569961e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    7.709882e-21, 1.027984e-20, -1.541976e-20, -2.569961e-21, -1.027984e-20, 
    1.541976e-20, -1.027984e-20, 7.709882e-21, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, -1.027984e-20, -7.709882e-21, 2.569961e-21, 7.709882e-21, 
    1.003089e-36, 0, 7.709882e-21, 1.027984e-20, 1.003089e-36, 0, 
    1.003089e-36, 5.139921e-21, -5.139921e-21, 0, 1.027984e-20, 5.139921e-21, 
    1.798972e-20, 1.027984e-20, 7.709882e-21, 1.027984e-20, 1.28498e-20, 
    -5.139921e-21, 1.28498e-20, 1.28498e-20, -1.027984e-20, 1.027984e-20, 
    -5.139921e-21, -7.709882e-21, -5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 0, -2.569961e-21, 0, 2.055969e-20, 2.055969e-20, 
    1.027984e-20, 1.027984e-20, 1.027984e-20, -1.28498e-20, 5.139921e-21, 
    -1.28498e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 7.709882e-21, 
    2.569961e-21, -2.569961e-21, 1.541976e-20, 5.139921e-21, 1.28498e-20, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 0, 
    -7.709882e-21, -5.139921e-21, -5.015443e-37, 2.569961e-21, 5.139921e-21, 
    7.709882e-21, -1.28498e-20, 0, -5.139921e-21, 2.569961e-21, 1.798972e-20, 
    5.139921e-21, -1.027984e-20, -2.569961e-21, 7.709882e-21, 7.709882e-21, 
    2.826957e-20, 1.541976e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, 1.003089e-36, 1.541976e-20, 0, -2.569961e-21, 
    1.798972e-20, 5.139921e-21, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    -1.28498e-20, -1.541976e-20, 2.569961e-21, -1.003089e-36, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 1.027984e-20, 0, -1.28498e-20, 0, 0, 
    2.055969e-20, 2.569961e-21, 1.027984e-20, 2.055969e-20, 1.798972e-20, 
    2.569961e-21, 2.569961e-21, -1.541976e-20, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, -1.541976e-20, 1.28498e-20, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, 7.709882e-21, 1.027984e-20, 2.569961e-21, 1.027984e-20, 
    2.569961e-21, 0, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 7.709882e-21, -5.139921e-21, 1.027984e-20, -1.541976e-20, 
    -7.709882e-21, 5.139921e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, -1.28498e-20, 0, -1.003089e-36, -2.569961e-21, 
    7.709882e-21, 1.027984e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, 
    -7.709882e-21, 1.003089e-36, -1.003089e-36, -1.027984e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, 1.003089e-36, 
    -2.569961e-21, 2.569961e-21, -5.015443e-37, -1.027984e-20, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, 2.569961e-21, -1.027984e-20, -7.709882e-21, 
    -2.569961e-21, 1.003089e-36, 1.003089e-36, 2.055969e-20, -1.027984e-20, 
    -5.139921e-21, -7.709882e-21, -1.541976e-20, -1.003089e-36, 1.28498e-20, 
    -5.139921e-21, 7.709882e-21, -7.709882e-21, -1.541976e-20, 5.139921e-21, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, 1.027984e-20, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 5.139921e-21, -1.28498e-20, -5.139921e-21, 
    -1.027984e-20, 1.28498e-20, -2.569961e-21, 0, -1.003089e-36, 
    1.003089e-36, 1.541976e-20, 7.709882e-21, -5.139921e-21, -2.569961e-21, 
    2.569961e-21, 5.139921e-21, -1.28498e-20, -5.139921e-21, -7.709882e-21,
  -5.139921e-21, -5.139921e-21, 5.139921e-21, 1.541976e-20, 7.709882e-21, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, -1.003089e-36, 1.027984e-20, 
    7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, 0, 
    -7.709882e-21, -2.569961e-21, -1.027984e-20, 0, 2.569961e-21, 
    -5.139921e-21, 1.28498e-20, 2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 1.28498e-20, -2.569961e-21, -1.027984e-20, 0, 
    5.139921e-21, 7.709882e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 1.28498e-20, 1.027984e-20, -1.027984e-20, 
    -2.569961e-21, 1.28498e-20, -7.709882e-21, 5.139921e-21, -1.28498e-20, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, 1.003089e-36, 7.709882e-21, 
    -1.027984e-20, -1.28498e-20, 2.569961e-21, 5.139921e-21, -1.003089e-36, 
    -1.027984e-20, 2.569961e-21, -5.139921e-21, 5.139921e-21, -1.798972e-20, 
    -2.055969e-20, 1.027984e-20, -5.139921e-21, -2.569961e-21, -1.027984e-20, 
    0, -2.569961e-21, 5.139921e-21, 1.28498e-20, 5.139921e-21, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 1.027984e-20, -1.027984e-20, 7.709882e-21, 
    2.569961e-21, 0, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    1.541976e-20, -2.569961e-21, 0, 1.027984e-20, -1.003089e-36, 
    2.569961e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, -5.139921e-21, 
    1.003089e-36, -2.569961e-21, 2.569961e-21, 5.139921e-21, 1.027984e-20, 
    -2.569961e-21, 1.541976e-20, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    -1.28498e-20, 1.798972e-20, 2.569961e-21, 1.28498e-20, 1.003089e-36, 
    7.709882e-21, 1.003089e-36, -7.709882e-21, -5.139921e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, 1.003089e-36, 5.139921e-21, 2.569961e-21, 
    1.003089e-36, 2.569961e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    1.541976e-20, 0, 1.28498e-20, 0, 2.569961e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, 0, -2.569961e-21, 
    -1.027984e-20, 1.027984e-20, -2.569961e-21, -7.709882e-21, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 0, 2.569961e-21, 0, 2.569961e-21, 0, 
    -2.569961e-21, 7.709882e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, 0, -7.709882e-21, 
    -1.541976e-20, 2.569961e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, 2.569961e-21, -1.798972e-20, 
    7.709882e-21, 0, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 1.28498e-20, 5.139921e-21, 
    5.139921e-21, 0, 1.003089e-36, 2.569961e-21, -2.569961e-21, 1.003089e-36, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, 
    1.027984e-20, 2.569961e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 
    2.569961e-21, -1.027984e-20, 0, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, -2.569961e-21, 1.027984e-20, 2.569961e-21, 1.027984e-20, 
    -2.569961e-21, -5.139921e-21, 0, 5.139921e-21, 0, -5.139921e-21, 
    -1.28498e-20, 5.139921e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, 0, 2.312965e-20, 1.28498e-20, 7.709882e-21, 
    -1.541976e-20, -7.709882e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 0, 1.003089e-36, 5.139921e-21, 0, 0, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, 0, -7.709882e-21, 
    7.709882e-21, 1.003089e-36, -2.569961e-21, -7.709882e-21, 5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 1.003089e-36, -1.027984e-20, 1.027984e-20, 
    2.569961e-21, 5.139921e-21, 1.027984e-20, -2.569961e-21, 0, 
    -7.709882e-21, 0, 1.28498e-20, -7.709882e-21, -1.541976e-20, 
    5.139921e-21, 0, 1.003089e-36, 1.541976e-20, -7.709882e-21, 1.003089e-36, 
    2.569961e-21, -7.709882e-21, 0, 1.027984e-20, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, -7.709882e-21, 0, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 7.709882e-21, 5.139921e-21, -1.28498e-20, 
    2.569961e-21, 0, -7.709882e-21, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, 1.027984e-20, -5.139921e-21, -2.569961e-21, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, -7.709882e-21, 
    0, -7.709882e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 
    1.027984e-20, 2.569961e-21, 1.28498e-20, 1.027984e-20, -5.139921e-21, 
    2.569961e-21, 5.139921e-21,
  -5.139921e-21, -5.139921e-21, -1.027984e-20, -7.709882e-21, 5.139921e-21, 
    -2.569961e-21, -1.28498e-20, -1.28498e-20, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, -1.027984e-20, -7.709882e-21, -2.569961e-21, 0, 
    1.027984e-20, -1.027984e-20, 2.569961e-21, 5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -1.798972e-20, -1.027984e-20, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -1.003089e-36, 0, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, 7.709882e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, 
    7.709882e-21, -7.709882e-21, -7.709882e-21, 1.003089e-36, 7.709882e-21, 
    -1.003089e-36, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, 2.569961e-21, 0, 2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -5.139921e-21, 1.541976e-20, -7.709882e-21, 
    2.569961e-21, -1.003089e-36, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, -7.709882e-21, 1.541976e-20, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, 0, 7.709882e-21, 2.569961e-21, -1.027984e-20, 
    7.709882e-21, -7.709882e-21, -5.139921e-21, -7.709882e-21, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -7.709882e-21, -1.027984e-20, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, 1.003089e-36, 1.28498e-20, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 
    5.139921e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, 0, 
    5.139921e-21, 1.28498e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    5.139921e-21, 1.28498e-20, -1.027984e-20, -2.569961e-21, 1.027984e-20, 0, 
    2.569961e-21, 7.709882e-21, 0, 7.709882e-21, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, 1.28498e-20, 5.139921e-21, 5.139921e-21, 2.569961e-21, 0, 
    5.139921e-21, -7.709882e-21, -7.709882e-21, 2.569961e-21, 1.541976e-20, 
    -2.569961e-21, -2.569961e-21, -1.027984e-20, -7.709882e-21, 0, 
    1.28498e-20, 7.709882e-21, -2.569961e-21, 7.709882e-21, 5.139921e-21, 
    -2.569961e-21, 0, 1.027984e-20, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, 1.027984e-20, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, -2.055969e-20, -1.798972e-20, 1.003089e-36, 
    0, 5.139921e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, 
    -1.28498e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, 1.541976e-20, 
    0, 0, -1.027984e-20, 0, -1.027984e-20, -1.003089e-36, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, -1.027984e-20, -1.798972e-20, 
    1.027984e-20, 7.709882e-21, -1.541976e-20, 0, 5.139921e-21, 0, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 2.569961e-21, -7.709882e-21, 
    -7.709882e-21, 1.541976e-20, -1.003089e-36, 5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 1.28498e-20, 2.569961e-21, -1.798972e-20, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 1.28498e-20, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 0, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, 7.709882e-21, 1.027984e-20, 
    5.139921e-21, -1.003089e-36, -2.569961e-21, 5.139921e-21, -1.003089e-36, 
    2.569961e-21, -1.28498e-20, -1.28498e-20, 1.798972e-20, -2.569961e-21, 
    -1.28498e-20, -1.003089e-36, 0, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, 1.003089e-36, -1.28498e-20, 
    1.28498e-20, -1.28498e-20, 0, 2.569961e-21, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, -1.798972e-20, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.28498e-20, -2.569961e-21, -1.027984e-20, 1.28498e-20, 0, 
    2.569961e-21, 2.569961e-21, -2.569961e-21, -1.798972e-20, 2.569961e-21, 
    1.541976e-20, 2.055969e-20, -2.569961e-21, 1.027984e-20, 1.003089e-36, 
    -1.28498e-20, -7.709882e-21, -1.541976e-20, -2.569961e-21, -1.027984e-20, 
    0, 7.709882e-21, 1.027984e-20, 5.139921e-21, 1.28498e-20, -1.003089e-36, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, 7.709882e-21, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 2.055969e-20, 7.709882e-21, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, 1.003089e-36, -1.28498e-20, -5.139921e-21, -7.709882e-21, 
    -1.28498e-20, 5.139921e-21, 0, -2.569961e-21, -1.28498e-20, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, -1.003089e-36, -2.569961e-21, 
    1.027984e-20, -2.569961e-21, -1.027984e-20, 0, -1.027984e-20, 
    1.541976e-20, 1.28498e-20, -5.139921e-21, 1.28498e-20, 1.28498e-20, 
    -7.709882e-21, 1.541976e-20, -1.28498e-20, -2.569961e-21, -1.027984e-20, 
    2.569961e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, 0, 
    7.709882e-21, 0, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -7.709882e-21, -1.003089e-36, 0, 1.027984e-20, -2.569961e-21, 
    7.709882e-21, 2.569961e-21,
  7.709882e-21, 2.569961e-21, -2.569961e-20, 1.541976e-20, 0, 1.027984e-20, 
    2.569961e-21, 5.139921e-21, -1.28498e-20, 2.055969e-20, 5.139921e-21, 
    -1.541976e-20, -2.569961e-21, -1.28498e-20, -7.709882e-21, 2.569961e-21, 
    2.055969e-20, -2.569961e-21, -2.569961e-21, 1.003089e-36, 5.139921e-21, 
    -2.569961e-21, 0, -1.027984e-20, 2.569961e-21, 1.027984e-20, 0, 
    -1.027984e-20, -5.139921e-21, 2.569961e-21, 5.139921e-21, 1.003089e-36, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    1.027984e-20, 7.709882e-21, -1.027984e-20, -1.28498e-20, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 7.709882e-21, -1.003089e-36, 7.709882e-21, 
    7.709882e-21, 2.569961e-21, 1.027984e-20, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, -1.541976e-20, 1.003089e-36, 1.28498e-20, -1.027984e-20, 
    5.139921e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 0, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, -2.569961e-21, 
    1.003089e-36, -5.139921e-21, 0, 7.709882e-21, -1.027984e-20, 
    -1.541976e-20, -1.027984e-20, -1.027984e-20, -2.569961e-21, 1.003089e-36, 
    -7.709882e-21, 1.28498e-20, 1.027984e-20, 1.027984e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -2.055969e-20, -7.709882e-21, 
    -1.541976e-20, -1.003089e-36, -5.139921e-21, -2.569961e-21, 7.709882e-21, 
    -5.139921e-21, 1.28498e-20, 7.709882e-21, 2.569961e-21, 2.055969e-20, 
    7.709882e-21, 1.027984e-20, -2.055969e-20, 2.569961e-21, -7.709882e-21, 
    7.709882e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 1.027984e-20, 
    2.569961e-21, 2.569961e-21, 1.541976e-20, 7.709882e-21, -2.569961e-21, 
    -1.541976e-20, 2.569961e-21, -1.28498e-20, 2.569961e-21, -7.709882e-21, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, 0, -5.139921e-21, 
    -1.28498e-20, -1.541976e-20, -1.003089e-36, -5.139921e-21, -1.28498e-20, 
    -7.709882e-21, 2.569961e-21, -1.027984e-20, -1.027984e-20, -7.709882e-21, 
    5.139921e-21, -1.003089e-36, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 0, -1.28498e-20, -7.709882e-21, 
    -2.569961e-21, -1.541976e-20, 1.28498e-20, -7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 0, 2.569961e-21, 2.055969e-20, -1.541976e-20, 
    -7.709882e-21, 7.709882e-21, -1.798972e-20, -1.541976e-20, 1.027984e-20, 
    -1.28498e-20, 1.003089e-36, -7.709882e-21, -7.709882e-21, -2.569961e-21, 
    5.139921e-21, -1.28498e-20, 1.027984e-20, -7.709882e-21, -1.798972e-20, 
    -5.139921e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    1.027984e-20, -5.139921e-21, -1.28498e-20, 7.709882e-21, 1.027984e-20, 
    1.28498e-20, -1.28498e-20, -2.569961e-21, -1.798972e-20, -7.709882e-21, 
    1.28498e-20, -1.28498e-20, -1.003089e-36, -2.569961e-21, 1.027984e-20, 
    1.027984e-20, 0, 7.709882e-21, -2.569961e-21, 2.569961e-21, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, -2.569961e-20, -7.709882e-21, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, -7.709882e-21, 
    1.027984e-20, -7.709882e-21, 7.709882e-21, -5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 0, -7.709882e-21, -5.139921e-21, -1.027984e-20, 
    1.798972e-20, -5.139921e-21, 7.709882e-21, -1.003089e-36, -1.798972e-20, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, -7.709882e-21, 1.28498e-20, 
    1.003089e-36, 1.798972e-20, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, 5.139921e-21, -1.541976e-20, -1.541976e-20, -2.569961e-21, 
    7.709882e-21, 7.709882e-21, 7.709882e-21, -1.003089e-36, -7.709882e-21, 
    0, 5.139921e-21, 1.541976e-20, 1.027984e-20, -7.709882e-21, 1.541976e-20, 
    1.003089e-36, -5.139921e-21, -5.139921e-21, -1.541976e-20, 2.569961e-21, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, -5.139921e-21, 1.28498e-20, 
    -1.28498e-20, -1.003089e-36, 7.709882e-21, -5.139921e-21, 1.541976e-20, 
    -1.027984e-20, 2.569961e-21, 1.28498e-20, 7.709882e-21, 2.569961e-21, 
    5.139921e-21, 1.027984e-20, -2.569961e-21, 2.569961e-21, -1.003089e-36, 
    1.541976e-20, -2.055969e-20, -5.139921e-21, -7.709882e-21, 5.139921e-21, 
    1.027984e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, -1.027984e-20, 
    0, 7.709882e-21, 5.139921e-21, 3.083953e-20, 0, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, -2.312965e-20, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 7.709882e-21, 1.027984e-20, 1.541976e-20, 
    7.709882e-21, -2.055969e-20, -2.312965e-20, 5.139921e-21, 2.569961e-21, 
    1.027984e-20, -1.027984e-20, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    1.027984e-20, -1.541976e-20, 7.709882e-21, -5.139921e-21, 2.569961e-20, 
    0, -1.027984e-20, 1.027984e-20, -1.541976e-20, -7.709882e-21, 
    -1.541976e-20, 5.139921e-21, 2.569961e-21, -7.709882e-21, 1.027984e-20, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, 7.709882e-21, -7.709882e-21, 5.139921e-21, -1.28498e-20, 
    0, 2.569961e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 2.569961e-20, 
    -7.709882e-21, 5.139921e-21,
  -5.139921e-21, -1.027984e-20, 1.541976e-20, -2.569961e-21, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, 7.709882e-21, 1.28498e-20, 
    -1.003089e-36, 1.027984e-20, -1.027984e-20, -5.139921e-21, 1.541976e-20, 
    -2.055969e-20, 5.139921e-21, 5.139921e-21, 5.015443e-37, -2.569961e-21, 
    -5.139921e-21, 1.027984e-20, 1.798972e-20, -1.027984e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 1.003089e-36, 1.28498e-20, 2.055969e-20, 
    -2.569961e-21, -1.003089e-36, 1.28498e-20, 5.139921e-21, -5.139921e-21, 
    -1.003089e-36, 1.541976e-20, -1.541976e-20, 0, 1.541976e-20, 
    -5.139921e-21, -1.003089e-36, 2.569961e-21, 1.798972e-20, 7.709882e-21, 
    -2.569961e-21, 1.003089e-36, 1.28498e-20, 1.003089e-36, 5.139921e-21, 
    -1.003089e-36, 1.28498e-20, 2.055969e-20, 2.826957e-20, -2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 1.027984e-20, 5.139921e-21, -2.312965e-20, 
    -1.027984e-20, 1.28498e-20, 5.139921e-21, 0, -1.541976e-20, 
    -7.709882e-21, 1.798972e-20, 5.139921e-21, -1.027984e-20, 2.569961e-21, 
    2.569961e-21, 1.798972e-20, 7.709882e-21, 2.569961e-21, -1.541976e-20, 
    7.709882e-21, -1.027984e-20, 7.709882e-21, -2.055969e-20, 1.28498e-20, 
    -3.009266e-36, 7.709882e-21, 5.139921e-21, -1.027984e-20, 7.709882e-21, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -1.798972e-20, 2.826957e-20, 1.003089e-36, 2.569961e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-20, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -1.541976e-20, 1.027984e-20, 1.28498e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.003089e-36, 5.139921e-21, -5.139921e-21, 
    1.798972e-20, 1.027984e-20, -5.139921e-21, 7.709882e-21, -5.139921e-21, 
    1.28498e-20, 5.139921e-21, 7.709882e-21, 0, 1.28498e-20, -1.027984e-20, 
    -1.541976e-20, -2.569961e-21, 5.139921e-21, -1.28498e-20, 1.027984e-20, 
    7.709882e-21, 1.027984e-20, 7.709882e-21, 5.139921e-21, 7.709882e-21, 
    2.569961e-21, 1.027984e-20, 5.139921e-21, -1.027984e-20, -1.003089e-36, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -7.709882e-21, 7.709882e-21, -1.027984e-20, 1.28498e-20, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, -2.569961e-21, 1.541976e-20, 
    1.798972e-20, -5.139921e-21, 7.709882e-21, 5.139921e-21, 5.139921e-21, 
    7.709882e-21, -1.027984e-20, -1.28498e-20, 7.709882e-21, -1.027984e-20, 
    -2.569961e-21, -5.139921e-21, 3.083953e-20, 7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 1.28498e-20, -7.709882e-21, -1.027984e-20, 7.709882e-21, 
    0, 1.027984e-20, -5.139921e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.798972e-20, 0, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, 1.28498e-20, -2.569961e-21, 2.569961e-21, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, -1.798972e-20, 1.541976e-20, 
    1.541976e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 2.312965e-20, 
    7.709882e-21, -1.798972e-20, -1.28498e-20, 7.709882e-21, 5.139921e-21, 
    1.541976e-20, -1.28498e-20, -1.027984e-20, 2.826957e-20, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, 1.28498e-20, 1.003089e-36, 7.709882e-21, -1.027984e-20, 
    1.798972e-20, -2.569961e-21, 7.709882e-21, 1.28498e-20, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, -5.139921e-21, 
    -1.027984e-20, -1.28498e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, 1.28498e-20, -1.027984e-20, -1.28498e-20, 
    -2.569961e-21, 7.709882e-21, 1.798972e-20, -1.027984e-20, 1.28498e-20, 
    7.709882e-21, -7.709882e-21, 2.569961e-21, 1.28498e-20, 2.826957e-20, 
    1.027984e-20, 2.569961e-21, 5.139921e-21, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 5.139921e-21, 1.28498e-20, -2.569961e-21, 1.28498e-20, 
    1.003089e-36, 1.027984e-20, -2.569961e-21, -3.009266e-36, 1.798972e-20, 
    -1.28498e-20, 7.709882e-21, 1.798972e-20, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-20, 2.569961e-21, 0, -2.569961e-21, 1.28498e-20, 
    -7.709882e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, 
    -1.28498e-20, -7.709882e-21, 2.055969e-20, -2.569961e-21, -1.027984e-20, 
    7.709882e-21, -2.569961e-21, 1.541976e-20, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, -1.798972e-20, 1.003089e-36, -1.28498e-20, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, -1.798972e-20, 1.027984e-20, 2.569961e-21, 
    1.003089e-36, 7.709882e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, 
    2.055969e-20, 2.569961e-21, -5.139921e-21, 5.139921e-21, 1.798972e-20, 
    1.003089e-36, 7.709882e-21, 2.569961e-21, 2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 1.798972e-20, -5.139921e-21, 7.709882e-21, 7.709882e-21, 
    -1.027984e-20, -1.541976e-20, 2.569961e-21, -7.709882e-21, -5.139921e-21, 
    1.798972e-20, -2.569961e-21, -1.541976e-20, -2.569961e-21, -2.569961e-21, 
    0, 1.003089e-36, -2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -1.027984e-20, -1.027984e-20,
  6.259378e-29, 6.259384e-29, 6.259382e-29, 6.259388e-29, 6.259385e-29, 
    6.259388e-29, 6.259379e-29, 6.259384e-29, 6.259381e-29, 6.259378e-29, 
    6.259398e-29, 6.259388e-29, 6.259407e-29, 6.259401e-29, 6.259417e-29, 
    6.259407e-29, 6.259419e-29, 6.259416e-29, 6.259423e-29, 6.259421e-29, 
    6.25943e-29, 6.259424e-29, 6.259435e-29, 6.259429e-29, 6.25943e-29, 
    6.259424e-29, 6.25939e-29, 6.259396e-29, 6.25939e-29, 6.25939e-29, 
    6.25939e-29, 6.259385e-29, 6.259382e-29, 6.259377e-29, 6.259378e-29, 
    6.259382e-29, 6.259391e-29, 6.259388e-29, 6.259395e-29, 6.259395e-29, 
    6.259404e-29, 6.2594e-29, 6.259414e-29, 6.25941e-29, 6.259422e-29, 
    6.259419e-29, 6.259421e-29, 6.25942e-29, 6.259421e-29, 6.259417e-29, 
    6.259419e-29, 6.259415e-29, 6.259401e-29, 6.259405e-29, 6.259392e-29, 
    6.259384e-29, 6.259379e-29, 6.259376e-29, 6.259376e-29, 6.259377e-29, 
    6.259382e-29, 6.259387e-29, 6.25939e-29, 6.259393e-29, 6.259395e-29, 
    6.259402e-29, 6.259406e-29, 6.259414e-29, 6.259413e-29, 6.259416e-29, 
    6.259418e-29, 6.259422e-29, 6.259422e-29, 6.259423e-29, 6.259416e-29, 
    6.259421e-29, 6.259412e-29, 6.259414e-29, 6.259396e-29, 6.259388e-29, 
    6.259385e-29, 6.259383e-29, 6.259376e-29, 6.259381e-29, 6.259379e-29, 
    6.259384e-29, 6.259386e-29, 6.259385e-29, 6.259393e-29, 6.25939e-29, 
    6.259407e-29, 6.259399e-29, 6.259418e-29, 6.259413e-29, 6.259419e-29, 
    6.259416e-29, 6.259421e-29, 6.259417e-29, 6.259424e-29, 6.259426e-29, 
    6.259425e-29, 6.259429e-29, 6.259416e-29, 6.259421e-29, 6.259385e-29, 
    6.259385e-29, 6.259386e-29, 6.259381e-29, 6.259381e-29, 6.259377e-29, 
    6.259381e-29, 6.259382e-29, 6.259386e-29, 6.259388e-29, 6.259391e-29, 
    6.259396e-29, 6.259401e-29, 6.259408e-29, 6.259414e-29, 6.259417e-29, 
    6.259415e-29, 6.259417e-29, 6.259415e-29, 6.259414e-29, 6.259425e-29, 
    6.259419e-29, 6.259428e-29, 6.259428e-29, 6.259423e-29, 6.259428e-29, 
    6.259385e-29, 6.259384e-29, 6.259379e-29, 6.259383e-29, 6.259377e-29, 
    6.25938e-29, 6.259382e-29, 6.25939e-29, 6.259391e-29, 6.259393e-29, 
    6.259396e-29, 6.2594e-29, 6.259407e-29, 6.259413e-29, 6.259419e-29, 
    6.259418e-29, 6.259418e-29, 6.259419e-29, 6.259416e-29, 6.25942e-29, 
    6.25942e-29, 6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259428e-29, 
    6.259426e-29, 6.259384e-29, 6.259386e-29, 6.259385e-29, 6.259387e-29, 
    6.259386e-29, 6.259393e-29, 6.259394e-29, 6.259404e-29, 6.2594e-29, 
    6.259406e-29, 6.259401e-29, 6.259402e-29, 6.259406e-29, 6.259401e-29, 
    6.259413e-29, 6.259405e-29, 6.259419e-29, 6.259411e-29, 6.25942e-29, 
    6.259419e-29, 6.259421e-29, 6.259423e-29, 6.259426e-29, 6.259431e-29, 
    6.25943e-29, 6.259434e-29, 6.25939e-29, 6.259392e-29, 6.259392e-29, 
    6.259394e-29, 6.259397e-29, 6.259401e-29, 6.259408e-29, 6.259406e-29, 
    6.259411e-29, 6.259412e-29, 6.259404e-29, 6.259409e-29, 6.259394e-29, 
    6.259396e-29, 6.259395e-29, 6.25939e-29, 6.259407e-29, 6.259398e-29, 
    6.259414e-29, 6.259409e-29, 6.259423e-29, 6.259416e-29, 6.259429e-29, 
    6.259435e-29, 6.25944e-29, 6.259447e-29, 6.259393e-29, 6.259391e-29, 
    6.259395e-29, 6.259399e-29, 6.259404e-29, 6.25941e-29, 6.25941e-29, 
    6.259411e-29, 6.259414e-29, 6.259416e-29, 6.259411e-29, 6.259417e-29, 
    6.259397e-29, 6.259407e-29, 6.259391e-29, 6.259396e-29, 6.259399e-29, 
    6.259398e-29, 6.259405e-29, 6.259407e-29, 6.259415e-29, 6.259411e-29, 
    6.259434e-29, 6.259423e-29, 6.259452e-29, 6.259444e-29, 6.259391e-29, 
    6.259393e-29, 6.259402e-29, 6.259398e-29, 6.25941e-29, 6.259413e-29, 
    6.259415e-29, 6.259418e-29, 6.259419e-29, 6.25942e-29, 6.259417e-29, 
    6.25942e-29, 6.25941e-29, 6.259414e-29, 6.259401e-29, 6.259404e-29, 
    6.259403e-29, 6.259401e-29, 6.259406e-29, 6.259411e-29, 6.259411e-29, 
    6.259413e-29, 6.259418e-29, 6.25941e-29, 6.259435e-29, 6.259419e-29, 
    6.259396e-29, 6.259401e-29, 6.259402e-29, 6.2594e-29, 6.259413e-29, 
    6.259408e-29, 6.25942e-29, 6.259417e-29, 6.259422e-29, 6.259419e-29, 
    6.259419e-29, 6.259416e-29, 6.259413e-29, 6.259408e-29, 6.259404e-29, 
    6.2594e-29, 6.259401e-29, 6.259405e-29, 6.259412e-29, 6.259419e-29, 
    6.259417e-29, 6.259422e-29, 6.259409e-29, 6.259414e-29, 6.259412e-29, 
    6.259417e-29, 6.259406e-29, 6.259416e-29, 6.259403e-29, 6.259404e-29, 
    6.259408e-29, 6.259414e-29, 6.259416e-29, 6.259418e-29, 6.259417e-29, 
    6.259412e-29, 6.259411e-29, 6.259408e-29, 6.259407e-29, 6.259404e-29, 
    6.259402e-29, 6.259404e-29, 6.259406e-29, 6.259412e-29, 6.259417e-29, 
    6.259423e-29, 6.259425e-29, 6.259431e-29, 6.259426e-29, 6.259435e-29, 
    6.259427e-29, 6.259441e-29, 6.259416e-29, 6.259427e-29, 6.259408e-29, 
    6.25941e-29, 6.259414e-29, 6.259422e-29, 6.259417e-29, 6.259423e-29, 
    6.259411e-29, 6.259405e-29, 6.259404e-29, 6.259401e-29, 6.259404e-29, 
    6.259403e-29, 6.259406e-29, 6.259405e-29, 6.259412e-29, 6.259408e-29, 
    6.259419e-29, 6.259423e-29, 6.259434e-29, 6.259441e-29, 6.259447e-29, 
    6.25945e-29, 6.259452e-29, 6.259452e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.138285e-10, 2.14772e-10, 2.145886e-10, 2.153497e-10, 2.149275e-10, 
    2.154258e-10, 2.140198e-10, 2.148095e-10, 2.143054e-10, 2.139135e-10, 
    2.168265e-10, 2.153836e-10, 2.183257e-10, 2.174053e-10, 2.197175e-10, 
    2.181824e-10, 2.20027e-10, 2.196732e-10, 2.207382e-10, 2.204331e-10, 
    2.217952e-10, 2.20879e-10, 2.225014e-10, 2.215764e-10, 2.217211e-10, 
    2.208487e-10, 2.15674e-10, 2.166469e-10, 2.156164e-10, 2.157551e-10, 
    2.156929e-10, 2.149362e-10, 2.145549e-10, 2.137565e-10, 2.139014e-10, 
    2.144879e-10, 2.158175e-10, 2.153662e-10, 2.165037e-10, 2.16478e-10, 
    2.177445e-10, 2.171735e-10, 2.193023e-10, 2.186972e-10, 2.204458e-10, 
    2.20006e-10, 2.204252e-10, 2.202981e-10, 2.204268e-10, 2.197818e-10, 
    2.200582e-10, 2.194907e-10, 2.172804e-10, 2.179299e-10, 2.159928e-10, 
    2.14828e-10, 2.140545e-10, 2.135056e-10, 2.135832e-10, 2.137311e-10, 
    2.144913e-10, 2.152061e-10, 2.157509e-10, 2.161153e-10, 2.164743e-10, 
    2.175611e-10, 2.181364e-10, 2.194246e-10, 2.191922e-10, 2.19586e-10, 
    2.199623e-10, 2.20594e-10, 2.2049e-10, 2.207683e-10, 2.195756e-10, 
    2.203683e-10, 2.190598e-10, 2.194177e-10, 2.165718e-10, 2.154879e-10, 
    2.150271e-10, 2.146239e-10, 2.136428e-10, 2.143203e-10, 2.140532e-10, 
    2.146887e-10, 2.150924e-10, 2.148927e-10, 2.161252e-10, 2.156461e-10, 
    2.181705e-10, 2.170831e-10, 2.199184e-10, 2.192399e-10, 2.20081e-10, 
    2.196518e-10, 2.203873e-10, 2.197254e-10, 2.208719e-10, 2.211216e-10, 
    2.20951e-10, 2.216064e-10, 2.196887e-10, 2.204251e-10, 2.148871e-10, 
    2.149197e-10, 2.150714e-10, 2.144045e-10, 2.143637e-10, 2.137525e-10, 
    2.142963e-10, 2.145279e-10, 2.151158e-10, 2.154636e-10, 2.157942e-10, 
    2.165211e-10, 2.173329e-10, 2.184682e-10, 2.192839e-10, 2.198307e-10, 
    2.194954e-10, 2.197914e-10, 2.194605e-10, 2.193054e-10, 2.21028e-10, 
    2.200607e-10, 2.215122e-10, 2.214318e-10, 2.20775e-10, 2.214409e-10, 
    2.149426e-10, 2.147552e-10, 2.141045e-10, 2.146137e-10, 2.136859e-10, 
    2.142052e-10, 2.145038e-10, 2.15656e-10, 2.159092e-10, 2.16144e-10, 
    2.166076e-10, 2.172027e-10, 2.182466e-10, 2.191549e-10, 2.199842e-10, 
    2.199234e-10, 2.199448e-10, 2.201301e-10, 2.196712e-10, 2.202054e-10, 
    2.20295e-10, 2.200606e-10, 2.214211e-10, 2.210324e-10, 2.214301e-10, 
    2.211771e-10, 2.148161e-10, 2.151314e-10, 2.14961e-10, 2.152815e-10, 
    2.150557e-10, 2.160595e-10, 2.163605e-10, 2.17769e-10, 2.17191e-10, 
    2.181109e-10, 2.172844e-10, 2.174309e-10, 2.181409e-10, 2.173291e-10, 
    2.191048e-10, 2.179009e-10, 2.201373e-10, 2.189349e-10, 2.202126e-10, 
    2.199806e-10, 2.203648e-10, 2.207088e-10, 2.211416e-10, 2.219403e-10, 
    2.217554e-10, 2.224233e-10, 2.156016e-10, 2.160106e-10, 2.159746e-10, 
    2.164027e-10, 2.167193e-10, 2.174056e-10, 2.185062e-10, 2.180923e-10, 
    2.188522e-10, 2.190048e-10, 2.178503e-10, 2.185591e-10, 2.162844e-10, 
    2.166518e-10, 2.164331e-10, 2.156338e-10, 2.181877e-10, 2.16877e-10, 
    2.192974e-10, 2.185873e-10, 2.206597e-10, 2.19629e-10, 2.216535e-10, 
    2.22519e-10, 2.233337e-10, 2.242857e-10, 2.162339e-10, 2.15956e-10, 
    2.164536e-10, 2.171422e-10, 2.177811e-10, 2.186306e-10, 2.187175e-10, 
    2.188766e-10, 2.192889e-10, 2.196355e-10, 2.189269e-10, 2.197224e-10, 
    2.16737e-10, 2.183014e-10, 2.158509e-10, 2.165887e-10, 2.171016e-10, 
    2.168766e-10, 2.18045e-10, 2.183204e-10, 2.194395e-10, 2.18861e-10, 
    2.223054e-10, 2.207814e-10, 2.250107e-10, 2.238287e-10, 2.158588e-10, 
    2.162329e-10, 2.17535e-10, 2.169155e-10, 2.186873e-10, 2.191234e-10, 
    2.19478e-10, 2.199313e-10, 2.199802e-10, 2.202488e-10, 2.198087e-10, 
    2.202314e-10, 2.186324e-10, 2.193469e-10, 2.173862e-10, 2.178634e-10, 
    2.176439e-10, 2.174031e-10, 2.181463e-10, 2.189381e-10, 2.18955e-10, 
    2.192089e-10, 2.199243e-10, 2.186945e-10, 2.22502e-10, 2.201504e-10, 
    2.166409e-10, 2.173614e-10, 2.174644e-10, 2.171853e-10, 2.190797e-10, 
    2.183933e-10, 2.202422e-10, 2.197425e-10, 2.205613e-10, 2.201544e-10, 
    2.200946e-10, 2.19572e-10, 2.192467e-10, 2.184247e-10, 2.17756e-10, 
    2.172258e-10, 2.173491e-10, 2.179315e-10, 2.189865e-10, 2.199846e-10, 
    2.19766e-10, 2.204991e-10, 2.185588e-10, 2.193724e-10, 2.190579e-10, 
    2.198779e-10, 2.180813e-10, 2.19611e-10, 2.176903e-10, 2.178587e-10, 
    2.183796e-10, 2.194275e-10, 2.196594e-10, 2.19907e-10, 2.197542e-10, 
    2.190133e-10, 2.188919e-10, 2.18367e-10, 2.18222e-10, 2.178221e-10, 
    2.174909e-10, 2.177935e-10, 2.181112e-10, 2.190136e-10, 2.198269e-10, 
    2.207137e-10, 2.209307e-10, 2.219667e-10, 2.211233e-10, 2.225151e-10, 
    2.213317e-10, 2.233803e-10, 2.196997e-10, 2.21297e-10, 2.184034e-10, 
    2.187151e-10, 2.192789e-10, 2.205721e-10, 2.19874e-10, 2.206905e-10, 
    2.188872e-10, 2.179516e-10, 2.177096e-10, 2.17258e-10, 2.177199e-10, 
    2.176824e-10, 2.181244e-10, 2.179823e-10, 2.190436e-10, 2.184735e-10, 
    2.200931e-10, 2.206841e-10, 2.223533e-10, 2.233766e-10, 2.244184e-10, 
    2.248784e-10, 2.250184e-10, 2.250769e-10 ;

 SOIL2N_TO_SOIL3N =
  1.527347e-11, 1.534086e-11, 1.532776e-11, 1.538212e-11, 1.535197e-11, 
    1.538756e-11, 1.528713e-11, 1.534354e-11, 1.530753e-11, 1.527954e-11, 
    1.548761e-11, 1.538454e-11, 1.559469e-11, 1.552895e-11, 1.56941e-11, 
    1.558446e-11, 1.571621e-11, 1.569095e-11, 1.576701e-11, 1.574522e-11, 
    1.584251e-11, 1.577707e-11, 1.589295e-11, 1.582688e-11, 1.583722e-11, 
    1.577491e-11, 1.540529e-11, 1.547478e-11, 1.540117e-11, 1.541108e-11, 
    1.540663e-11, 1.535259e-11, 1.532535e-11, 1.526832e-11, 1.527867e-11, 
    1.532056e-11, 1.541553e-11, 1.53833e-11, 1.546455e-11, 1.546272e-11, 
    1.555318e-11, 1.551239e-11, 1.566445e-11, 1.562123e-11, 1.574613e-11, 
    1.571472e-11, 1.574465e-11, 1.573558e-11, 1.574477e-11, 1.56987e-11, 
    1.571844e-11, 1.567791e-11, 1.552003e-11, 1.556642e-11, 1.542805e-11, 
    1.534486e-11, 1.52896e-11, 1.52504e-11, 1.525594e-11, 1.526651e-11, 
    1.532081e-11, 1.537187e-11, 1.541078e-11, 1.54368e-11, 1.546245e-11, 
    1.554008e-11, 1.558117e-11, 1.567319e-11, 1.565659e-11, 1.568472e-11, 
    1.571159e-11, 1.575672e-11, 1.574929e-11, 1.576917e-11, 1.568397e-11, 
    1.574059e-11, 1.564713e-11, 1.567269e-11, 1.546941e-11, 1.539199e-11, 
    1.535908e-11, 1.533028e-11, 1.52602e-11, 1.530859e-11, 1.528952e-11, 
    1.533491e-11, 1.536374e-11, 1.534948e-11, 1.543752e-11, 1.540329e-11, 
    1.558361e-11, 1.550594e-11, 1.570846e-11, 1.565999e-11, 1.572007e-11, 
    1.568942e-11, 1.574195e-11, 1.569467e-11, 1.577657e-11, 1.57944e-11, 
    1.578221e-11, 1.582903e-11, 1.569205e-11, 1.574465e-11, 1.534908e-11, 
    1.535141e-11, 1.536225e-11, 1.53146e-11, 1.531169e-11, 1.526803e-11, 
    1.530688e-11, 1.532342e-11, 1.536542e-11, 1.539026e-11, 1.541387e-11, 
    1.546579e-11, 1.552378e-11, 1.560487e-11, 1.566314e-11, 1.570219e-11, 
    1.567824e-11, 1.569939e-11, 1.567575e-11, 1.566467e-11, 1.578772e-11, 
    1.571862e-11, 1.58223e-11, 1.581656e-11, 1.576964e-11, 1.581721e-11, 
    1.535304e-11, 1.533965e-11, 1.529318e-11, 1.532955e-11, 1.526328e-11, 
    1.530037e-11, 1.53217e-11, 1.5404e-11, 1.542209e-11, 1.543886e-11, 
    1.547197e-11, 1.551448e-11, 1.558904e-11, 1.565392e-11, 1.571316e-11, 
    1.570882e-11, 1.571034e-11, 1.572358e-11, 1.56908e-11, 1.572896e-11, 
    1.573536e-11, 1.571862e-11, 1.581579e-11, 1.578803e-11, 1.581644e-11, 
    1.579836e-11, 1.534401e-11, 1.536653e-11, 1.535436e-11, 1.537725e-11, 
    1.536112e-11, 1.543283e-11, 1.545432e-11, 1.555493e-11, 1.551364e-11, 
    1.557935e-11, 1.552032e-11, 1.553078e-11, 1.558149e-11, 1.552351e-11, 
    1.565034e-11, 1.556435e-11, 1.572409e-11, 1.56382e-11, 1.572947e-11, 
    1.57129e-11, 1.574034e-11, 1.576491e-11, 1.579583e-11, 1.585288e-11, 
    1.583967e-11, 1.588738e-11, 1.540011e-11, 1.542933e-11, 1.542676e-11, 
    1.545734e-11, 1.547995e-11, 1.552897e-11, 1.560759e-11, 1.557802e-11, 
    1.56323e-11, 1.56432e-11, 1.556074e-11, 1.561136e-11, 1.544889e-11, 
    1.547513e-11, 1.545951e-11, 1.540242e-11, 1.558483e-11, 1.549121e-11, 
    1.56641e-11, 1.561338e-11, 1.576141e-11, 1.568779e-11, 1.58324e-11, 
    1.589421e-11, 1.595241e-11, 1.602041e-11, 1.544528e-11, 1.542542e-11, 
    1.546097e-11, 1.551015e-11, 1.555579e-11, 1.561647e-11, 1.562268e-11, 
    1.563405e-11, 1.566349e-11, 1.568825e-11, 1.563764e-11, 1.569445e-11, 
    1.548122e-11, 1.559296e-11, 1.541792e-11, 1.547062e-11, 1.550726e-11, 
    1.549119e-11, 1.557465e-11, 1.559432e-11, 1.567425e-11, 1.563293e-11, 
    1.587896e-11, 1.57701e-11, 1.607219e-11, 1.598776e-11, 1.541849e-11, 
    1.544521e-11, 1.553821e-11, 1.549396e-11, 1.562052e-11, 1.565167e-11, 
    1.5677e-11, 1.570938e-11, 1.571287e-11, 1.573205e-11, 1.570062e-11, 
    1.573081e-11, 1.56166e-11, 1.566764e-11, 1.552758e-11, 1.556167e-11, 
    1.554599e-11, 1.552879e-11, 1.558188e-11, 1.563843e-11, 1.563965e-11, 
    1.565778e-11, 1.570888e-11, 1.562103e-11, 1.5893e-11, 1.572503e-11, 
    1.547435e-11, 1.552582e-11, 1.553317e-11, 1.551323e-11, 1.564855e-11, 
    1.559952e-11, 1.573159e-11, 1.569589e-11, 1.575438e-11, 1.572532e-11, 
    1.572104e-11, 1.568371e-11, 1.566048e-11, 1.560177e-11, 1.5554e-11, 
    1.551613e-11, 1.552493e-11, 1.556654e-11, 1.564189e-11, 1.571319e-11, 
    1.569757e-11, 1.574993e-11, 1.561135e-11, 1.566946e-11, 1.564699e-11, 
    1.570556e-11, 1.557724e-11, 1.56865e-11, 1.554931e-11, 1.556134e-11, 
    1.559855e-11, 1.567339e-11, 1.568996e-11, 1.570764e-11, 1.569673e-11, 
    1.564381e-11, 1.563514e-11, 1.559764e-11, 1.558729e-11, 1.555872e-11, 
    1.553506e-11, 1.555668e-11, 1.557937e-11, 1.564383e-11, 1.570192e-11, 
    1.576526e-11, 1.578077e-11, 1.585477e-11, 1.579452e-11, 1.589393e-11, 
    1.580941e-11, 1.595573e-11, 1.569284e-11, 1.580693e-11, 1.560024e-11, 
    1.562251e-11, 1.566278e-11, 1.575515e-11, 1.570529e-11, 1.576361e-11, 
    1.56348e-11, 1.556797e-11, 1.555069e-11, 1.551843e-11, 1.555142e-11, 
    1.554874e-11, 1.558031e-11, 1.557017e-11, 1.564597e-11, 1.560525e-11, 
    1.572093e-11, 1.576315e-11, 1.588238e-11, 1.595547e-11, 1.602989e-11, 
    1.606274e-11, 1.607274e-11, 1.607692e-11 ;

 SOIL2N_vr =
  1.818719, 1.818721, 1.81872, 1.818722, 1.818721, 1.818722, 1.81872, 
    1.818721, 1.81872, 1.818719, 1.818724, 1.818722, 1.818726, 1.818725, 
    1.818728, 1.818726, 1.818729, 1.818728, 1.81873, 1.81873, 1.818732, 
    1.81873, 1.818733, 1.818731, 1.818732, 1.81873, 1.818722, 1.818724, 
    1.818722, 1.818722, 1.818722, 1.818721, 1.81872, 1.818719, 1.818719, 
    1.81872, 1.818722, 1.818722, 1.818723, 1.818723, 1.818725, 1.818725, 
    1.818728, 1.818727, 1.81873, 1.818729, 1.81873, 1.818729, 1.81873, 
    1.818729, 1.818729, 1.818728, 1.818725, 1.818726, 1.818723, 1.818721, 
    1.81872, 1.818719, 1.818719, 1.818719, 1.81872, 1.818721, 1.818722, 
    1.818723, 1.818723, 1.818725, 1.818726, 1.818728, 1.818728, 1.818728, 
    1.818729, 1.81873, 1.81873, 1.81873, 1.818728, 1.818729, 1.818727, 
    1.818728, 1.818724, 1.818722, 1.818721, 1.818721, 1.818719, 1.81872, 
    1.81872, 1.818721, 1.818721, 1.818721, 1.818723, 1.818722, 1.818726, 
    1.818724, 1.818729, 1.818728, 1.818729, 1.818728, 1.81873, 1.818728, 
    1.81873, 1.818731, 1.81873, 1.818731, 1.818728, 1.81873, 1.818721, 
    1.818721, 1.818721, 1.81872, 1.81872, 1.818719, 1.81872, 1.81872, 
    1.818721, 1.818722, 1.818722, 1.818723, 1.818725, 1.818727, 1.818728, 
    1.818729, 1.818728, 1.818729, 1.818728, 1.818728, 1.81873, 1.818729, 
    1.818731, 1.818731, 1.81873, 1.818731, 1.818721, 1.818721, 1.81872, 
    1.818721, 1.818719, 1.81872, 1.81872, 1.818722, 1.818722, 1.818723, 
    1.818724, 1.818725, 1.818726, 1.818728, 1.818729, 1.818729, 1.818729, 
    1.818729, 1.818728, 1.818729, 1.818729, 1.818729, 1.818731, 1.81873, 
    1.818731, 1.818731, 1.818721, 1.818721, 1.818721, 1.818722, 1.818721, 
    1.818723, 1.818723, 1.818725, 1.818725, 1.818726, 1.818725, 1.818725, 
    1.818726, 1.818725, 1.818727, 1.818726, 1.818729, 1.818727, 1.818729, 
    1.818729, 1.818729, 1.81873, 1.818731, 1.818732, 1.818732, 1.818733, 
    1.818722, 1.818723, 1.818723, 1.818723, 1.818724, 1.818725, 1.818727, 
    1.818726, 1.818727, 1.818727, 1.818726, 1.818727, 1.818723, 1.818724, 
    1.818723, 1.818722, 1.818726, 1.818724, 1.818728, 1.818727, 1.81873, 
    1.818728, 1.818731, 1.818733, 1.818734, 1.818735, 1.818723, 1.818723, 
    1.818723, 1.818725, 1.818725, 1.818727, 1.818727, 1.818727, 1.818728, 
    1.818728, 1.818727, 1.818728, 1.818724, 1.818726, 1.818722, 1.818724, 
    1.818724, 1.818724, 1.818726, 1.818726, 1.818728, 1.818727, 1.818732, 
    1.81873, 1.818737, 1.818735, 1.818722, 1.818723, 1.818725, 1.818724, 
    1.818727, 1.818727, 1.818728, 1.818729, 1.818729, 1.818729, 1.818729, 
    1.818729, 1.818727, 1.818728, 1.818725, 1.818726, 1.818725, 1.818725, 
    1.818726, 1.818727, 1.818727, 1.818728, 1.818729, 1.818727, 1.818733, 
    1.818729, 1.818724, 1.818725, 1.818725, 1.818725, 1.818727, 1.818726, 
    1.818729, 1.818728, 1.81873, 1.818729, 1.818729, 1.818728, 1.818728, 
    1.818726, 1.818725, 1.818725, 1.818725, 1.818726, 1.818727, 1.818729, 
    1.818729, 1.81873, 1.818727, 1.818728, 1.818727, 1.818729, 1.818726, 
    1.818728, 1.818725, 1.818726, 1.818726, 1.818728, 1.818728, 1.818729, 
    1.818728, 1.818727, 1.818727, 1.818726, 1.818726, 1.818725, 1.818725, 
    1.818725, 1.818726, 1.818727, 1.818729, 1.81873, 1.81873, 1.818732, 
    1.818731, 1.818733, 1.818731, 1.818734, 1.818728, 1.818731, 1.818726, 
    1.818727, 1.818728, 1.81873, 1.818729, 1.81873, 1.818727, 1.818726, 
    1.818725, 1.818725, 1.818725, 1.818725, 1.818726, 1.818726, 1.818727, 
    1.818727, 1.818729, 1.81873, 1.818733, 1.818734, 1.818736, 1.818736, 
    1.818737, 1.818737,
  1.818668, 1.818669, 1.818669, 1.818671, 1.81867, 1.818671, 1.818668, 
    1.81867, 1.818668, 1.818668, 1.818673, 1.818671, 1.818676, 1.818675, 
    1.818679, 1.818676, 1.81868, 1.818679, 1.818681, 1.818681, 1.818683, 
    1.818681, 1.818685, 1.818683, 1.818683, 1.818681, 1.818671, 1.818673, 
    1.818671, 1.818671, 1.818671, 1.81867, 1.818669, 1.818667, 1.818668, 
    1.818669, 1.818671, 1.818671, 1.818673, 1.818673, 1.818675, 1.818674, 
    1.818678, 1.818677, 1.818681, 1.81868, 1.818681, 1.81868, 1.818681, 
    1.818679, 1.81868, 1.818679, 1.818674, 1.818676, 1.818672, 1.81867, 
    1.818668, 1.818667, 1.818667, 1.818667, 1.818669, 1.81867, 1.818671, 
    1.818672, 1.818673, 1.818675, 1.818676, 1.818679, 1.818678, 1.818679, 
    1.81868, 1.818681, 1.818681, 1.818681, 1.818679, 1.81868, 1.818678, 
    1.818678, 1.818673, 1.818671, 1.81867, 1.818669, 1.818667, 1.818669, 
    1.818668, 1.818669, 1.81867, 1.81867, 1.818672, 1.818671, 1.818676, 
    1.818674, 1.81868, 1.818678, 1.81868, 1.818679, 1.81868, 1.818679, 
    1.818681, 1.818682, 1.818682, 1.818683, 1.818679, 1.818681, 1.81867, 
    1.81867, 1.81867, 1.818669, 1.818669, 1.818667, 1.818668, 1.818669, 
    1.81867, 1.818671, 1.818671, 1.818673, 1.818674, 1.818677, 1.818678, 
    1.818679, 1.818679, 1.818679, 1.818679, 1.818678, 1.818682, 1.81868, 
    1.818683, 1.818682, 1.818681, 1.818683, 1.81867, 1.818669, 1.818668, 
    1.818669, 1.818667, 1.818668, 1.818669, 1.818671, 1.818672, 1.818672, 
    1.818673, 1.818674, 1.818676, 1.818678, 1.81868, 1.81868, 1.81868, 
    1.81868, 1.818679, 1.81868, 1.81868, 1.81868, 1.818682, 1.818682, 
    1.818682, 1.818682, 1.81867, 1.81867, 1.81867, 1.818671, 1.81867, 
    1.818672, 1.818673, 1.818675, 1.818674, 1.818676, 1.818674, 1.818675, 
    1.818676, 1.818674, 1.818678, 1.818676, 1.81868, 1.818678, 1.81868, 
    1.81868, 1.81868, 1.818681, 1.818682, 1.818684, 1.818683, 1.818684, 
    1.818671, 1.818672, 1.818672, 1.818673, 1.818673, 1.818675, 1.818677, 
    1.818676, 1.818677, 1.818678, 1.818676, 1.818677, 1.818672, 1.818673, 
    1.818673, 1.818671, 1.818676, 1.818674, 1.818678, 1.818677, 1.818681, 
    1.818679, 1.818683, 1.818685, 1.818686, 1.818688, 1.818672, 1.818672, 
    1.818673, 1.818674, 1.818675, 1.818677, 1.818677, 1.818678, 1.818678, 
    1.818679, 1.818678, 1.818679, 1.818673, 1.818676, 1.818672, 1.818673, 
    1.818674, 1.818674, 1.818676, 1.818676, 1.818679, 1.818677, 1.818684, 
    1.818681, 1.818689, 1.818687, 1.818672, 1.818672, 1.818675, 1.818674, 
    1.818677, 1.818678, 1.818679, 1.81868, 1.81868, 1.81868, 1.818679, 
    1.81868, 1.818677, 1.818678, 1.818675, 1.818676, 1.818675, 1.818675, 
    1.818676, 1.818678, 1.818678, 1.818678, 1.81868, 1.818677, 1.818685, 
    1.81868, 1.818673, 1.818675, 1.818675, 1.818674, 1.818678, 1.818677, 
    1.81868, 1.818679, 1.818681, 1.81868, 1.81868, 1.818679, 1.818678, 
    1.818677, 1.818675, 1.818674, 1.818675, 1.818676, 1.818678, 1.81868, 
    1.818679, 1.818681, 1.818677, 1.818678, 1.818678, 1.818679, 1.818676, 
    1.818679, 1.818675, 1.818676, 1.818676, 1.818679, 1.818679, 1.81868, 
    1.818679, 1.818678, 1.818678, 1.818676, 1.818676, 1.818675, 1.818675, 
    1.818675, 1.818676, 1.818678, 1.818679, 1.818681, 1.818681, 1.818684, 
    1.818682, 1.818685, 1.818682, 1.818686, 1.818679, 1.818682, 1.818677, 
    1.818677, 1.818678, 1.818681, 1.818679, 1.818681, 1.818678, 1.818676, 
    1.818675, 1.818674, 1.818675, 1.818675, 1.818676, 1.818676, 1.818678, 
    1.818677, 1.81868, 1.818681, 1.818684, 1.818686, 1.818688, 1.818689, 
    1.818689, 1.81869,
  1.818639, 1.818641, 1.818641, 1.818642, 1.818642, 1.818643, 1.81864, 
    1.818641, 1.81864, 1.818639, 1.818646, 1.818642, 1.818649, 1.818647, 
    1.818652, 1.818648, 1.818653, 1.818652, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.818656, 1.818656, 1.818654, 1.818643, 1.818645, 
    1.818643, 1.818643, 1.818643, 1.818642, 1.818641, 1.818639, 1.818639, 
    1.818641, 1.818643, 1.818642, 1.818645, 1.818645, 1.818648, 1.818646, 
    1.818651, 1.81865, 1.818653, 1.818652, 1.818653, 1.818653, 1.818653, 
    1.818652, 1.818653, 1.818651, 1.818647, 1.818648, 1.818644, 1.818641, 
    1.81864, 1.818638, 1.818639, 1.818639, 1.818641, 1.818642, 1.818643, 
    1.818644, 1.818645, 1.818647, 1.818648, 1.818651, 1.818651, 1.818652, 
    1.818652, 1.818654, 1.818653, 1.818654, 1.818651, 1.818653, 1.81865, 
    1.818651, 1.818645, 1.818643, 1.818642, 1.818641, 1.818639, 1.81864, 
    1.81864, 1.818641, 1.818642, 1.818641, 1.818644, 1.818643, 1.818648, 
    1.818646, 1.818652, 1.818651, 1.818653, 1.818652, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818654, 1.818656, 1.818652, 1.818653, 1.818641, 
    1.818642, 1.818642, 1.81864, 1.81864, 1.818639, 1.81864, 1.818641, 
    1.818642, 1.818643, 1.818643, 1.818645, 1.818647, 1.818649, 1.818651, 
    1.818652, 1.818651, 1.818652, 1.818651, 1.818651, 1.818655, 1.818653, 
    1.818656, 1.818655, 1.818654, 1.818655, 1.818642, 1.818641, 1.81864, 
    1.818641, 1.818639, 1.81864, 1.818641, 1.818643, 1.818644, 1.818644, 
    1.818645, 1.818646, 1.818649, 1.818651, 1.818652, 1.818652, 1.818652, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818653, 1.818655, 1.818655, 
    1.818655, 1.818655, 1.818641, 1.818642, 1.818642, 1.818642, 1.818642, 
    1.818644, 1.818645, 1.818648, 1.818646, 1.818648, 1.818647, 1.818647, 
    1.818648, 1.818647, 1.81865, 1.818648, 1.818653, 1.81865, 1.818653, 
    1.818652, 1.818653, 1.818654, 1.818655, 1.818657, 1.818656, 1.818658, 
    1.818643, 1.818644, 1.818644, 1.818645, 1.818645, 1.818647, 1.818649, 
    1.818648, 1.81865, 1.81865, 1.818648, 1.818649, 1.818644, 1.818645, 
    1.818645, 1.818643, 1.818648, 1.818646, 1.818651, 1.818649, 1.818654, 
    1.818652, 1.818656, 1.818658, 1.81866, 1.818662, 1.818644, 1.818644, 
    1.818645, 1.818646, 1.818648, 1.818649, 1.81865, 1.81865, 1.818651, 
    1.818652, 1.81865, 1.818652, 1.818645, 1.818649, 1.818643, 1.818645, 
    1.818646, 1.818646, 1.818648, 1.818649, 1.818651, 1.81865, 1.818657, 
    1.818654, 1.818663, 1.818661, 1.818644, 1.818644, 1.818647, 1.818646, 
    1.81865, 1.81865, 1.818651, 1.818652, 1.818652, 1.818653, 1.818652, 
    1.818653, 1.818649, 1.818651, 1.818647, 1.818648, 1.818647, 1.818647, 
    1.818648, 1.81865, 1.81865, 1.818651, 1.818652, 1.81865, 1.818658, 
    1.818653, 1.818645, 1.818647, 1.818647, 1.818646, 1.81865, 1.818649, 
    1.818653, 1.818652, 1.818654, 1.818653, 1.818653, 1.818651, 1.818651, 
    1.818649, 1.818648, 1.818646, 1.818647, 1.818648, 1.81865, 1.818652, 
    1.818652, 1.818653, 1.818649, 1.818651, 1.81865, 1.818652, 1.818648, 
    1.818652, 1.818648, 1.818648, 1.818649, 1.818651, 1.818652, 1.818652, 
    1.818652, 1.81865, 1.81865, 1.818649, 1.818649, 1.818648, 1.818647, 
    1.818648, 1.818648, 1.81865, 1.818652, 1.818654, 1.818654, 1.818657, 
    1.818655, 1.818658, 1.818655, 1.81866, 1.818652, 1.818655, 1.818649, 
    1.81865, 1.818651, 1.818654, 1.818652, 1.818654, 1.81865, 1.818648, 
    1.818648, 1.818647, 1.818648, 1.818647, 1.818648, 1.818648, 1.81865, 
    1.818649, 1.818653, 1.818654, 1.818657, 1.81866, 1.818662, 1.818663, 
    1.818663, 1.818663,
  1.818617, 1.818619, 1.818619, 1.818621, 1.81862, 1.818621, 1.818618, 
    1.818619, 1.818618, 1.818618, 1.818624, 1.818621, 1.818627, 1.818625, 
    1.81863, 1.818627, 1.818631, 1.81863, 1.818632, 1.818632, 1.818635, 
    1.818633, 1.818636, 1.818634, 1.818635, 1.818633, 1.818621, 1.818624, 
    1.818621, 1.818622, 1.818622, 1.81862, 1.818619, 1.818617, 1.818618, 
    1.818619, 1.818622, 1.818621, 1.818623, 1.818623, 1.818626, 1.818625, 
    1.818629, 1.818628, 1.818632, 1.818631, 1.818632, 1.818632, 1.818632, 
    1.81863, 1.818631, 1.81863, 1.818625, 1.818626, 1.818622, 1.81862, 
    1.818618, 1.818617, 1.818617, 1.818617, 1.818619, 1.81862, 1.818622, 
    1.818622, 1.818623, 1.818626, 1.818627, 1.81863, 1.818629, 1.81863, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.81863, 1.818632, 1.818629, 
    1.81863, 1.818623, 1.818621, 1.81862, 1.818619, 1.818617, 1.818618, 
    1.818618, 1.818619, 1.81862, 1.81862, 1.818622, 1.818621, 1.818627, 
    1.818624, 1.818631, 1.818629, 1.818631, 1.81863, 1.818632, 1.81863, 
    1.818633, 1.818633, 1.818633, 1.818634, 1.81863, 1.818632, 1.81862, 
    1.81862, 1.81862, 1.818619, 1.818619, 1.818617, 1.818618, 1.818619, 
    1.81862, 1.818621, 1.818622, 1.818623, 1.818625, 1.818628, 1.818629, 
    1.818631, 1.81863, 1.81863, 1.81863, 1.818629, 1.818633, 1.818631, 
    1.818634, 1.818634, 1.818633, 1.818634, 1.81862, 1.818619, 1.818618, 
    1.818619, 1.818617, 1.818618, 1.818619, 1.818621, 1.818622, 1.818622, 
    1.818623, 1.818625, 1.818627, 1.818629, 1.818631, 1.818631, 1.818631, 
    1.818631, 1.81863, 1.818631, 1.818632, 1.818631, 1.818634, 1.818633, 
    1.818634, 1.818633, 1.818619, 1.81862, 1.81862, 1.818621, 1.81862, 
    1.818622, 1.818623, 1.818626, 1.818625, 1.818627, 1.818625, 1.818625, 
    1.818627, 1.818625, 1.818629, 1.818626, 1.818631, 1.818629, 1.818631, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.818635, 1.818635, 1.818636, 
    1.818621, 1.818622, 1.818622, 1.818623, 1.818624, 1.818625, 1.818628, 
    1.818627, 1.818628, 1.818629, 1.818626, 1.818628, 1.818623, 1.818624, 
    1.818623, 1.818621, 1.818627, 1.818624, 1.818629, 1.818628, 1.818632, 
    1.81863, 1.818635, 1.818636, 1.818638, 1.81864, 1.818623, 1.818622, 
    1.818623, 1.818625, 1.818626, 1.818628, 1.818628, 1.818628, 1.818629, 
    1.81863, 1.818629, 1.81863, 1.818624, 1.818627, 1.818622, 1.818623, 
    1.818624, 1.818624, 1.818627, 1.818627, 1.81863, 1.818628, 1.818636, 
    1.818633, 1.818642, 1.818639, 1.818622, 1.818623, 1.818625, 1.818624, 
    1.818628, 1.818629, 1.81863, 1.818631, 1.818631, 1.818631, 1.81863, 
    1.818631, 1.818628, 1.81863, 1.818625, 1.818626, 1.818626, 1.818625, 
    1.818627, 1.818629, 1.818629, 1.818629, 1.818631, 1.818628, 1.818636, 
    1.818631, 1.818624, 1.818625, 1.818625, 1.818625, 1.818629, 1.818627, 
    1.818631, 1.81863, 1.818632, 1.818631, 1.818631, 1.81863, 1.818629, 
    1.818627, 1.818626, 1.818625, 1.818625, 1.818626, 1.818629, 1.818631, 
    1.81863, 1.818632, 1.818628, 1.81863, 1.818629, 1.818631, 1.818627, 
    1.81863, 1.818626, 1.818626, 1.818627, 1.81863, 1.81863, 1.818631, 
    1.81863, 1.818629, 1.818628, 1.818627, 1.818627, 1.818626, 1.818625, 
    1.818626, 1.818627, 1.818629, 1.81863, 1.818632, 1.818633, 1.818635, 
    1.818633, 1.818636, 1.818634, 1.818638, 1.81863, 1.818634, 1.818627, 
    1.818628, 1.818629, 1.818632, 1.818631, 1.818632, 1.818628, 1.818626, 
    1.818626, 1.818625, 1.818626, 1.818626, 1.818627, 1.818627, 1.818629, 
    1.818628, 1.818631, 1.818632, 1.818636, 1.818638, 1.818641, 1.818642, 
    1.818642, 1.818642,
  1.818569, 1.81857, 1.81857, 1.818572, 1.818571, 1.818572, 1.818569, 
    1.81857, 1.81857, 1.818569, 1.818574, 1.818572, 1.818577, 1.818576, 
    1.81858, 1.818577, 1.818581, 1.81858, 1.818582, 1.818581, 1.818584, 
    1.818582, 1.818585, 1.818583, 1.818584, 1.818582, 1.818572, 1.818574, 
    1.818572, 1.818572, 1.818572, 1.818571, 1.81857, 1.818568, 1.818569, 
    1.81857, 1.818572, 1.818572, 1.818574, 1.818574, 1.818576, 1.818575, 
    1.818579, 1.818578, 1.818581, 1.818581, 1.818581, 1.818581, 1.818581, 
    1.81858, 1.818581, 1.818579, 1.818575, 1.818576, 1.818573, 1.81857, 
    1.818569, 1.818568, 1.818568, 1.818568, 1.81857, 1.818571, 1.818572, 
    1.818573, 1.818574, 1.818576, 1.818577, 1.818579, 1.818579, 1.81858, 
    1.81858, 1.818582, 1.818581, 1.818582, 1.81858, 1.818581, 1.818579, 
    1.818579, 1.818574, 1.818572, 1.818571, 1.81857, 1.818568, 1.81857, 
    1.818569, 1.81857, 1.818571, 1.818571, 1.818573, 1.818572, 1.818577, 
    1.818575, 1.81858, 1.818579, 1.818581, 1.81858, 1.818581, 1.81858, 
    1.818582, 1.818583, 1.818582, 1.818583, 1.81858, 1.818581, 1.818571, 
    1.818571, 1.818571, 1.81857, 1.81857, 1.818568, 1.81857, 1.81857, 
    1.818571, 1.818572, 1.818572, 1.818574, 1.818575, 1.818578, 1.818579, 
    1.81858, 1.818579, 1.81858, 1.818579, 1.818579, 1.818582, 1.818581, 
    1.818583, 1.818583, 1.818582, 1.818583, 1.818571, 1.81857, 1.818569, 
    1.81857, 1.818568, 1.818569, 1.81857, 1.818572, 1.818573, 1.818573, 
    1.818574, 1.818575, 1.818577, 1.818579, 1.81858, 1.81858, 1.81858, 
    1.818581, 1.81858, 1.818581, 1.818581, 1.818581, 1.818583, 1.818582, 
    1.818583, 1.818583, 1.81857, 1.818571, 1.818571, 1.818571, 1.818571, 
    1.818573, 1.818573, 1.818576, 1.818575, 1.818577, 1.818575, 1.818576, 
    1.818577, 1.818575, 1.818579, 1.818576, 1.818581, 1.818578, 1.818581, 
    1.81858, 1.818581, 1.818582, 1.818583, 1.818584, 1.818584, 1.818585, 
    1.818572, 1.818573, 1.818573, 1.818574, 1.818574, 1.818576, 1.818578, 
    1.818577, 1.818578, 1.818579, 1.818576, 1.818578, 1.818573, 1.818574, 
    1.818574, 1.818572, 1.818577, 1.818574, 1.818579, 1.818578, 1.818582, 
    1.81858, 1.818584, 1.818585, 1.818587, 1.818589, 1.818573, 1.818573, 
    1.818574, 1.818575, 1.818576, 1.818578, 1.818578, 1.818578, 1.818579, 
    1.81858, 1.818578, 1.81858, 1.818574, 1.818577, 1.818573, 1.818574, 
    1.818575, 1.818574, 1.818577, 1.818577, 1.818579, 1.818578, 1.818585, 
    1.818582, 1.81859, 1.818588, 1.818573, 1.818573, 1.818576, 1.818575, 
    1.818578, 1.818579, 1.818579, 1.81858, 1.81858, 1.818581, 1.81858, 
    1.818581, 1.818578, 1.818579, 1.818576, 1.818576, 1.818576, 1.818576, 
    1.818577, 1.818578, 1.818578, 1.818579, 1.81858, 1.818578, 1.818585, 
    1.818581, 1.818574, 1.818575, 1.818576, 1.818575, 1.818579, 1.818577, 
    1.818581, 1.81858, 1.818582, 1.818581, 1.818581, 1.81858, 1.818579, 
    1.818577, 1.818576, 1.818575, 1.818575, 1.818576, 1.818578, 1.81858, 
    1.81858, 1.818581, 1.818578, 1.818579, 1.818579, 1.81858, 1.818577, 
    1.81858, 1.818576, 1.818576, 1.818577, 1.818579, 1.81858, 1.81858, 
    1.81858, 1.818579, 1.818578, 1.818577, 1.818577, 1.818576, 1.818576, 
    1.818576, 1.818577, 1.818579, 1.81858, 1.818582, 1.818582, 1.818584, 
    1.818583, 1.818585, 1.818583, 1.818587, 1.81858, 1.818583, 1.818577, 
    1.818578, 1.818579, 1.818582, 1.81858, 1.818582, 1.818578, 1.818577, 
    1.818576, 1.818575, 1.818576, 1.818576, 1.818577, 1.818577, 1.818579, 
    1.818578, 1.818581, 1.818582, 1.818585, 1.818587, 1.818589, 1.81859, 
    1.81859, 1.81859,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.293663e-09, 1.299371e-09, 1.298261e-09, 1.302865e-09, 1.300312e-09, 
    1.303326e-09, 1.29482e-09, 1.299597e-09, 1.296548e-09, 1.294177e-09, 
    1.3118e-09, 1.303071e-09, 1.32087e-09, 1.315302e-09, 1.329291e-09, 
    1.320004e-09, 1.331163e-09, 1.329023e-09, 1.335466e-09, 1.33362e-09, 
    1.341861e-09, 1.336318e-09, 1.346133e-09, 1.340537e-09, 1.341412e-09, 
    1.336135e-09, 1.304828e-09, 1.310714e-09, 1.304479e-09, 1.305318e-09, 
    1.304942e-09, 1.300364e-09, 1.298057e-09, 1.293227e-09, 1.294104e-09, 
    1.297652e-09, 1.305696e-09, 1.302965e-09, 1.309847e-09, 1.309692e-09, 
    1.317354e-09, 1.3139e-09, 1.326779e-09, 1.323118e-09, 1.333697e-09, 
    1.331037e-09, 1.333572e-09, 1.332803e-09, 1.333582e-09, 1.32968e-09, 
    1.331352e-09, 1.327919e-09, 1.314546e-09, 1.318476e-09, 1.306756e-09, 
    1.299709e-09, 1.29503e-09, 1.291709e-09, 1.292178e-09, 1.293073e-09, 
    1.297672e-09, 1.301997e-09, 1.305293e-09, 1.307497e-09, 1.30967e-09, 
    1.316245e-09, 1.319725e-09, 1.327519e-09, 1.326113e-09, 1.328495e-09, 
    1.330772e-09, 1.334594e-09, 1.333965e-09, 1.335649e-09, 1.328433e-09, 
    1.333228e-09, 1.325312e-09, 1.327477e-09, 1.310259e-09, 1.303702e-09, 
    1.300914e-09, 1.298475e-09, 1.292539e-09, 1.296638e-09, 1.295022e-09, 
    1.298866e-09, 1.301309e-09, 1.300101e-09, 1.307558e-09, 1.304659e-09, 
    1.319932e-09, 1.313353e-09, 1.330506e-09, 1.326401e-09, 1.33149e-09, 
    1.328894e-09, 1.333343e-09, 1.329339e-09, 1.336275e-09, 1.337786e-09, 
    1.336753e-09, 1.340719e-09, 1.329117e-09, 1.333572e-09, 1.300067e-09, 
    1.300264e-09, 1.301182e-09, 1.297147e-09, 1.2969e-09, 1.293203e-09, 
    1.296493e-09, 1.297894e-09, 1.301451e-09, 1.303555e-09, 1.305555e-09, 
    1.309952e-09, 1.314864e-09, 1.321733e-09, 1.326668e-09, 1.329976e-09, 
    1.327947e-09, 1.329738e-09, 1.327736e-09, 1.326798e-09, 1.33722e-09, 
    1.331367e-09, 1.340149e-09, 1.339663e-09, 1.335689e-09, 1.339717e-09, 
    1.300403e-09, 1.299269e-09, 1.295332e-09, 1.298413e-09, 1.2928e-09, 
    1.295942e-09, 1.297748e-09, 1.304719e-09, 1.306251e-09, 1.307671e-09, 
    1.310476e-09, 1.314076e-09, 1.320392e-09, 1.325887e-09, 1.330904e-09, 
    1.330537e-09, 1.330666e-09, 1.331787e-09, 1.329011e-09, 1.332243e-09, 
    1.332785e-09, 1.331367e-09, 1.339598e-09, 1.337246e-09, 1.339652e-09, 
    1.338121e-09, 1.299637e-09, 1.301545e-09, 1.300514e-09, 1.302453e-09, 
    1.301087e-09, 1.30716e-09, 1.308981e-09, 1.317502e-09, 1.314005e-09, 
    1.319571e-09, 1.314571e-09, 1.315457e-09, 1.319752e-09, 1.314841e-09, 
    1.325584e-09, 1.3183e-09, 1.33183e-09, 1.324556e-09, 1.332286e-09, 
    1.330883e-09, 1.333207e-09, 1.335288e-09, 1.337907e-09, 1.342739e-09, 
    1.34162e-09, 1.345661e-09, 1.30439e-09, 1.306864e-09, 1.306647e-09, 
    1.309236e-09, 1.311152e-09, 1.315304e-09, 1.321963e-09, 1.319459e-09, 
    1.324056e-09, 1.324979e-09, 1.317994e-09, 1.322283e-09, 1.308521e-09, 
    1.310744e-09, 1.30942e-09, 1.304585e-09, 1.320035e-09, 1.312106e-09, 
    1.326749e-09, 1.322453e-09, 1.334991e-09, 1.328755e-09, 1.341004e-09, 
    1.34624e-09, 1.351169e-09, 1.356928e-09, 1.308215e-09, 1.306534e-09, 
    1.309544e-09, 1.31371e-09, 1.317576e-09, 1.322715e-09, 1.323241e-09, 
    1.324204e-09, 1.326698e-09, 1.328795e-09, 1.324508e-09, 1.32932e-09, 
    1.311259e-09, 1.320724e-09, 1.305898e-09, 1.310362e-09, 1.313465e-09, 
    1.312104e-09, 1.319172e-09, 1.320839e-09, 1.327609e-09, 1.324109e-09, 
    1.344947e-09, 1.335728e-09, 1.361315e-09, 1.354163e-09, 1.305946e-09, 
    1.308209e-09, 1.316087e-09, 1.312339e-09, 1.323058e-09, 1.325697e-09, 
    1.327842e-09, 1.330584e-09, 1.33088e-09, 1.332505e-09, 1.329843e-09, 
    1.3324e-09, 1.322726e-09, 1.327049e-09, 1.315186e-09, 1.318073e-09, 
    1.316745e-09, 1.315288e-09, 1.319785e-09, 1.324575e-09, 1.324678e-09, 
    1.326214e-09, 1.330542e-09, 1.323102e-09, 1.346137e-09, 1.33191e-09, 
    1.310677e-09, 1.315037e-09, 1.31566e-09, 1.313971e-09, 1.325432e-09, 
    1.321279e-09, 1.332465e-09, 1.329442e-09, 1.334396e-09, 1.331934e-09, 
    1.331572e-09, 1.328411e-09, 1.326442e-09, 1.32147e-09, 1.317424e-09, 
    1.314216e-09, 1.314962e-09, 1.318486e-09, 1.324868e-09, 1.330907e-09, 
    1.329584e-09, 1.334019e-09, 1.322281e-09, 1.327203e-09, 1.3253e-09, 
    1.330261e-09, 1.319392e-09, 1.328647e-09, 1.317026e-09, 1.318045e-09, 
    1.321197e-09, 1.327536e-09, 1.32894e-09, 1.330437e-09, 1.329513e-09, 
    1.325031e-09, 1.324296e-09, 1.32112e-09, 1.320243e-09, 1.317824e-09, 
    1.31582e-09, 1.31765e-09, 1.319573e-09, 1.325033e-09, 1.329953e-09, 
    1.335318e-09, 1.336631e-09, 1.342899e-09, 1.337796e-09, 1.346216e-09, 
    1.339057e-09, 1.351451e-09, 1.329183e-09, 1.338847e-09, 1.32134e-09, 
    1.323226e-09, 1.326637e-09, 1.334461e-09, 1.330238e-09, 1.335178e-09, 
    1.324268e-09, 1.318607e-09, 1.317143e-09, 1.314411e-09, 1.317206e-09, 
    1.316978e-09, 1.319652e-09, 1.318793e-09, 1.325214e-09, 1.321765e-09, 
    1.331563e-09, 1.335139e-09, 1.345237e-09, 1.351429e-09, 1.357731e-09, 
    1.360514e-09, 1.361361e-09, 1.361715e-09 ;

 SOIL2_HR_S3 =
  9.240448e-11, 9.281221e-11, 9.273295e-11, 9.306182e-11, 9.287939e-11, 
    9.309473e-11, 9.248715e-11, 9.282839e-11, 9.261055e-11, 9.244119e-11, 
    9.370003e-11, 9.307649e-11, 9.434788e-11, 9.395015e-11, 9.494933e-11, 
    9.428597e-11, 9.50831e-11, 9.493022e-11, 9.539042e-11, 9.525858e-11, 
    9.584719e-11, 9.545127e-11, 9.615236e-11, 9.575266e-11, 9.581517e-11, 
    9.543821e-11, 9.320199e-11, 9.362239e-11, 9.317708e-11, 9.323702e-11, 
    9.321013e-11, 9.288315e-11, 9.271837e-11, 9.237333e-11, 9.243597e-11, 
    9.26894e-11, 9.326398e-11, 9.306895e-11, 9.356053e-11, 9.354943e-11, 
    9.409674e-11, 9.384996e-11, 9.476993e-11, 9.450845e-11, 9.526408e-11, 
    9.507404e-11, 9.525515e-11, 9.520024e-11, 9.525587e-11, 9.497715e-11, 
    9.509656e-11, 9.485132e-11, 9.389618e-11, 9.417687e-11, 9.333972e-11, 
    9.283638e-11, 9.250211e-11, 9.22649e-11, 9.229844e-11, 9.236236e-11, 
    9.269088e-11, 9.299979e-11, 9.32352e-11, 9.339267e-11, 9.354784e-11, 
    9.401747e-11, 9.42661e-11, 9.482279e-11, 9.472234e-11, 9.489252e-11, 
    9.505514e-11, 9.532813e-11, 9.52832e-11, 9.540347e-11, 9.488805e-11, 
    9.523059e-11, 9.466512e-11, 9.481978e-11, 9.358995e-11, 9.312157e-11, 
    9.292243e-11, 9.274818e-11, 9.232422e-11, 9.261699e-11, 9.250158e-11, 
    9.277618e-11, 9.295065e-11, 9.286436e-11, 9.339698e-11, 9.318991e-11, 
    9.428083e-11, 9.381092e-11, 9.503617e-11, 9.474296e-11, 9.510645e-11, 
    9.492097e-11, 9.523878e-11, 9.495275e-11, 9.544823e-11, 9.555613e-11, 
    9.548239e-11, 9.576563e-11, 9.49369e-11, 9.525514e-11, 9.286194e-11, 
    9.287602e-11, 9.294158e-11, 9.265335e-11, 9.263572e-11, 9.237161e-11, 
    9.260662e-11, 9.27067e-11, 9.296078e-11, 9.311105e-11, 9.325392e-11, 
    9.356804e-11, 9.391886e-11, 9.440947e-11, 9.476197e-11, 9.499826e-11, 
    9.485337e-11, 9.498129e-11, 9.483829e-11, 9.477127e-11, 9.551569e-11, 
    9.509768e-11, 9.572489e-11, 9.569019e-11, 9.540633e-11, 9.56941e-11, 
    9.28859e-11, 9.280491e-11, 9.252371e-11, 9.274378e-11, 9.234285e-11, 
    9.256725e-11, 9.269629e-11, 9.319422e-11, 9.330364e-11, 9.340508e-11, 
    9.360545e-11, 9.386259e-11, 9.43137e-11, 9.470624e-11, 9.50646e-11, 
    9.503834e-11, 9.504759e-11, 9.512763e-11, 9.492934e-11, 9.516019e-11, 
    9.519893e-11, 9.509763e-11, 9.568554e-11, 9.551758e-11, 9.568945e-11, 
    9.558009e-11, 9.283124e-11, 9.296752e-11, 9.289387e-11, 9.303235e-11, 
    9.293479e-11, 9.336858e-11, 9.349865e-11, 9.410731e-11, 9.385753e-11, 
    9.425508e-11, 9.389792e-11, 9.39612e-11, 9.426802e-11, 9.391722e-11, 
    9.468458e-11, 9.41643e-11, 9.513074e-11, 9.461114e-11, 9.516331e-11, 
    9.506305e-11, 9.522905e-11, 9.537773e-11, 9.556478e-11, 9.590991e-11, 
    9.583e-11, 9.611864e-11, 9.317069e-11, 9.334745e-11, 9.33319e-11, 
    9.351689e-11, 9.36537e-11, 9.395026e-11, 9.44259e-11, 9.424705e-11, 
    9.457542e-11, 9.464134e-11, 9.414246e-11, 9.444875e-11, 9.346576e-11, 
    9.362455e-11, 9.353001e-11, 9.318463e-11, 9.428824e-11, 9.372184e-11, 
    9.476779e-11, 9.446093e-11, 9.535653e-11, 9.491111e-11, 9.5786e-11, 
    9.616e-11, 9.651208e-11, 9.692346e-11, 9.344393e-11, 9.332382e-11, 
    9.353889e-11, 9.383644e-11, 9.411256e-11, 9.447964e-11, 9.451721e-11, 
    9.458598e-11, 9.476412e-11, 9.49139e-11, 9.460771e-11, 9.495145e-11, 
    9.366136e-11, 9.433741e-11, 9.327841e-11, 9.359726e-11, 9.38189e-11, 
    9.372169e-11, 9.422661e-11, 9.434561e-11, 9.482921e-11, 9.457922e-11, 
    9.606768e-11, 9.540911e-11, 9.723675e-11, 9.672596e-11, 9.328185e-11, 
    9.344352e-11, 9.400618e-11, 9.373847e-11, 9.450415e-11, 9.469264e-11, 
    9.484587e-11, 9.504172e-11, 9.506288e-11, 9.517893e-11, 9.498876e-11, 
    9.517143e-11, 9.448042e-11, 9.478921e-11, 9.394189e-11, 9.414811e-11, 
    9.405324e-11, 9.394917e-11, 9.427036e-11, 9.461253e-11, 9.461985e-11, 
    9.472957e-11, 9.503872e-11, 9.450726e-11, 9.615264e-11, 9.513643e-11, 
    9.361981e-11, 9.39312e-11, 9.39757e-11, 9.385508e-11, 9.467373e-11, 
    9.43771e-11, 9.517611e-11, 9.496016e-11, 9.531399e-11, 9.513817e-11, 
    9.511229e-11, 9.488647e-11, 9.474588e-11, 9.439069e-11, 9.410171e-11, 
    9.387257e-11, 9.392585e-11, 9.417755e-11, 9.463346e-11, 9.506479e-11, 
    9.49703e-11, 9.52871e-11, 9.444864e-11, 9.48002e-11, 9.466431e-11, 
    9.501865e-11, 9.424229e-11, 9.490333e-11, 9.407332e-11, 9.414609e-11, 
    9.437121e-11, 9.482403e-11, 9.492425e-11, 9.503122e-11, 9.496522e-11, 
    9.464504e-11, 9.459259e-11, 9.436574e-11, 9.430309e-11, 9.413025e-11, 
    9.398714e-11, 9.411789e-11, 9.425519e-11, 9.464518e-11, 9.499664e-11, 
    9.537984e-11, 9.547363e-11, 9.592133e-11, 9.555685e-11, 9.61583e-11, 
    9.564691e-11, 9.65322e-11, 9.494167e-11, 9.563191e-11, 9.438145e-11, 
    9.451617e-11, 9.47598e-11, 9.531868e-11, 9.501698e-11, 9.536982e-11, 
    9.459054e-11, 9.418624e-11, 9.408165e-11, 9.38865e-11, 9.408611e-11, 
    9.406988e-11, 9.42609e-11, 9.419951e-11, 9.465813e-11, 9.441178e-11, 
    9.511164e-11, 9.536704e-11, 9.608839e-11, 9.65306e-11, 9.698082e-11, 
    9.717958e-11, 9.724007e-11, 9.726536e-11 ;

 SOIL3C =
  5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611 ;

 SOIL3C_TO_SOIL1C =
  2.55107e-11, 2.562324e-11, 2.560136e-11, 2.569213e-11, 2.564178e-11, 
    2.570122e-11, 2.553352e-11, 2.56277e-11, 2.556758e-11, 2.552083e-11, 
    2.586829e-11, 2.569618e-11, 2.604711e-11, 2.593733e-11, 2.621312e-11, 
    2.603002e-11, 2.625004e-11, 2.620784e-11, 2.633486e-11, 2.629848e-11, 
    2.646094e-11, 2.635166e-11, 2.654517e-11, 2.643485e-11, 2.64521e-11, 
    2.634806e-11, 2.573082e-11, 2.584686e-11, 2.572395e-11, 2.574049e-11, 
    2.573307e-11, 2.564282e-11, 2.559734e-11, 2.55021e-11, 2.551939e-11, 
    2.558934e-11, 2.574794e-11, 2.56941e-11, 2.582979e-11, 2.582672e-11, 
    2.597779e-11, 2.590968e-11, 2.61636e-11, 2.609143e-11, 2.629999e-11, 
    2.624754e-11, 2.629753e-11, 2.628237e-11, 2.629773e-11, 2.62208e-11, 
    2.625376e-11, 2.618607e-11, 2.592243e-11, 2.599991e-11, 2.576884e-11, 
    2.562991e-11, 2.553764e-11, 2.547217e-11, 2.548143e-11, 2.549907e-11, 
    2.558975e-11, 2.567501e-11, 2.573999e-11, 2.578346e-11, 2.582628e-11, 
    2.595591e-11, 2.602454e-11, 2.617819e-11, 2.615047e-11, 2.619744e-11, 
    2.624232e-11, 2.631767e-11, 2.630527e-11, 2.633847e-11, 2.61962e-11, 
    2.629075e-11, 2.613467e-11, 2.617736e-11, 2.583791e-11, 2.570863e-11, 
    2.565366e-11, 2.560557e-11, 2.548855e-11, 2.556936e-11, 2.55375e-11, 
    2.561329e-11, 2.566145e-11, 2.563763e-11, 2.578465e-11, 2.572749e-11, 
    2.60286e-11, 2.58989e-11, 2.623709e-11, 2.615616e-11, 2.625648e-11, 
    2.620529e-11, 2.629301e-11, 2.621406e-11, 2.635082e-11, 2.63806e-11, 
    2.636025e-11, 2.643843e-11, 2.620969e-11, 2.629753e-11, 2.563697e-11, 
    2.564085e-11, 2.565895e-11, 2.557939e-11, 2.557453e-11, 2.550163e-11, 
    2.556649e-11, 2.559412e-11, 2.566425e-11, 2.570572e-11, 2.574516e-11, 
    2.583186e-11, 2.592869e-11, 2.606411e-11, 2.61614e-11, 2.622662e-11, 
    2.618663e-11, 2.622194e-11, 2.618247e-11, 2.616397e-11, 2.636944e-11, 
    2.625406e-11, 2.642719e-11, 2.641761e-11, 2.633926e-11, 2.641868e-11, 
    2.564358e-11, 2.562122e-11, 2.554361e-11, 2.560435e-11, 2.549369e-11, 
    2.555563e-11, 2.559124e-11, 2.572868e-11, 2.575888e-11, 2.578688e-11, 
    2.584219e-11, 2.591316e-11, 2.603768e-11, 2.614602e-11, 2.624493e-11, 
    2.623769e-11, 2.624024e-11, 2.626233e-11, 2.62076e-11, 2.627132e-11, 
    2.628201e-11, 2.625405e-11, 2.641632e-11, 2.636996e-11, 2.64174e-11, 
    2.638722e-11, 2.562849e-11, 2.566611e-11, 2.564578e-11, 2.5684e-11, 
    2.565707e-11, 2.577681e-11, 2.581271e-11, 2.598071e-11, 2.591176e-11, 
    2.602149e-11, 2.592291e-11, 2.594038e-11, 2.602507e-11, 2.592824e-11, 
    2.614004e-11, 2.599644e-11, 2.626319e-11, 2.611977e-11, 2.627218e-11, 
    2.624451e-11, 2.629033e-11, 2.633136e-11, 2.638299e-11, 2.647825e-11, 
    2.645619e-11, 2.653587e-11, 2.572218e-11, 2.577097e-11, 2.576668e-11, 
    2.581774e-11, 2.585551e-11, 2.593736e-11, 2.606865e-11, 2.601928e-11, 
    2.610991e-11, 2.612811e-11, 2.599041e-11, 2.607495e-11, 2.580363e-11, 
    2.584746e-11, 2.582136e-11, 2.572603e-11, 2.603065e-11, 2.587431e-11, 
    2.616301e-11, 2.607831e-11, 2.632551e-11, 2.620257e-11, 2.644405e-11, 
    2.654728e-11, 2.664446e-11, 2.6758e-11, 2.57976e-11, 2.576445e-11, 
    2.582382e-11, 2.590594e-11, 2.598216e-11, 2.608348e-11, 2.609385e-11, 
    2.611283e-11, 2.6162e-11, 2.620334e-11, 2.611883e-11, 2.62137e-11, 
    2.585762e-11, 2.604422e-11, 2.575192e-11, 2.583993e-11, 2.59011e-11, 
    2.587427e-11, 2.601364e-11, 2.604648e-11, 2.617996e-11, 2.611096e-11, 
    2.65218e-11, 2.634002e-11, 2.684448e-11, 2.670349e-11, 2.575287e-11, 
    2.579749e-11, 2.59528e-11, 2.58789e-11, 2.609024e-11, 2.614227e-11, 
    2.618456e-11, 2.623862e-11, 2.624446e-11, 2.627649e-11, 2.6224e-11, 
    2.627442e-11, 2.608369e-11, 2.616892e-11, 2.593505e-11, 2.599197e-11, 
    2.596578e-11, 2.593706e-11, 2.602571e-11, 2.612015e-11, 2.612218e-11, 
    2.615246e-11, 2.623779e-11, 2.60911e-11, 2.654525e-11, 2.626476e-11, 
    2.584615e-11, 2.59321e-11, 2.594438e-11, 2.591109e-11, 2.613705e-11, 
    2.605517e-11, 2.627571e-11, 2.621611e-11, 2.631377e-11, 2.626524e-11, 
    2.62581e-11, 2.619577e-11, 2.615696e-11, 2.605893e-11, 2.597916e-11, 
    2.591592e-11, 2.593062e-11, 2.60001e-11, 2.612593e-11, 2.624499e-11, 
    2.621891e-11, 2.630635e-11, 2.607492e-11, 2.617196e-11, 2.613445e-11, 
    2.623225e-11, 2.601796e-11, 2.620042e-11, 2.597133e-11, 2.599141e-11, 
    2.605355e-11, 2.617853e-11, 2.62062e-11, 2.623572e-11, 2.62175e-11, 
    2.612913e-11, 2.611465e-11, 2.605204e-11, 2.603475e-11, 2.598704e-11, 
    2.594754e-11, 2.598363e-11, 2.602153e-11, 2.612917e-11, 2.622618e-11, 
    2.633194e-11, 2.635783e-11, 2.648141e-11, 2.63808e-11, 2.654681e-11, 
    2.640566e-11, 2.665001e-11, 2.6211e-11, 2.640152e-11, 2.605638e-11, 
    2.609356e-11, 2.616081e-11, 2.631506e-11, 2.623179e-11, 2.632918e-11, 
    2.611409e-11, 2.600249e-11, 2.597363e-11, 2.591976e-11, 2.597486e-11, 
    2.597038e-11, 2.60231e-11, 2.600616e-11, 2.613274e-11, 2.606475e-11, 
    2.625792e-11, 2.632841e-11, 2.652751e-11, 2.664957e-11, 2.677383e-11, 
    2.68287e-11, 2.684539e-11, 2.685237e-11 ;

 SOIL3C_vr =
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  -1.027984e-20, 2.569961e-21, 1.003089e-36, -7.709882e-21, 0, -2.569961e-21, 
    2.569961e-20, 2.569961e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -1.28498e-20, 1.798972e-20, 1.798972e-20, 7.709882e-21, -2.312965e-20, 
    -2.569961e-21, 5.139921e-21, -1.003089e-36, -5.139921e-21, -1.003089e-36, 
    -7.709882e-21, 7.709882e-21, 7.709882e-21, -1.541976e-20, -1.027984e-20, 
    5.139921e-21, 7.709882e-21, -1.003089e-36, 2.569961e-21, -7.709882e-21, 
    -7.709882e-21, 2.569961e-21, 1.027984e-20, -1.027984e-20, 0, 
    -1.28498e-20, -5.139921e-21, 1.027984e-20, -7.709882e-21, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, -1.28498e-20, 2.569961e-21, 
    7.709882e-21, 1.027984e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, 
    -1.541976e-20, 7.709882e-21, -7.709882e-21, -7.709882e-21, 5.139921e-21, 
    -1.027984e-20, -2.569961e-21, -7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -1.798972e-20, -1.027984e-20, 1.027984e-20, -1.541976e-20, 5.139921e-21, 
    1.003089e-36, -5.139921e-21, -7.709882e-21, -1.027984e-20, 0, 0, 
    1.027984e-20, -1.798972e-20, 2.569961e-21, -1.541976e-20, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 1.027984e-20, -7.709882e-21, 1.027984e-20, 1.003089e-36, 
    2.569961e-21, 1.28498e-20, 5.139921e-21, 1.027984e-20, -7.709882e-21, 
    1.027984e-20, 1.28498e-20, -1.541976e-20, 7.709882e-21, 5.139921e-21, 
    7.709882e-21, 1.541976e-20, -5.139921e-21, -1.027984e-20, 2.569961e-21, 
    -2.569961e-21, 1.003089e-36, 0, 1.027984e-20, -7.709882e-21, 0, 
    7.709882e-21, -7.709882e-21, -2.312965e-20, -5.139921e-21, 0, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    7.709882e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, -7.709882e-21, 
    5.139921e-21, 1.003089e-36, -1.798972e-20, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, 7.709882e-21, 5.139921e-21, 
    1.003089e-36, -1.541976e-20, 2.569961e-21, 5.139921e-21, -1.28498e-20, 
    -5.139921e-21, 2.569961e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, 7.709882e-21, 1.28498e-20, 
    1.027984e-20, 2.569961e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, -7.709882e-21, 1.541976e-20, 1.003089e-36, -1.541976e-20, 
    5.139921e-21, -2.569961e-21, 5.139921e-21, 1.027984e-20, 7.709882e-21, 
    -5.139921e-21, 7.709882e-21, -2.569961e-21, -1.003089e-36, -1.28498e-20, 
    2.569961e-21, -1.027984e-20, 7.709882e-21, -1.027984e-20, -1.027984e-20, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, 1.027984e-20, 7.709882e-21, 
    -1.027984e-20, 1.027984e-20, -1.798972e-20, -1.027984e-20, -1.541976e-20, 
    -5.139921e-21, -1.28498e-20, -5.139921e-21, 5.139921e-21, 7.709882e-21, 
    -7.709882e-21, 2.569961e-21, -1.541976e-20, 1.28498e-20, 0, 
    -2.569961e-21, -5.139921e-21, 1.28498e-20, 5.139921e-21, 5.139921e-21, 0, 
    -7.709882e-21, 2.312965e-20, 1.541976e-20, 7.709882e-21, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, 7.709882e-21, -1.027984e-20, 
    -7.709882e-21, 2.569961e-21, 1.28498e-20, 1.027984e-20, -5.139921e-21, 
    -7.709882e-21, -7.709882e-21, 0, -1.027984e-20, 1.027984e-20, 
    1.027984e-20, 2.055969e-20, -1.027984e-20, -1.541976e-20, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, 5.139921e-21, -1.003089e-36, 
    -1.541976e-20, 0, 5.139921e-21, 7.709882e-21, -2.055969e-20, 
    -1.541976e-20, 1.28498e-20, -1.027984e-20, -2.569961e-21, 1.003089e-36, 
    -1.027984e-20, 1.027984e-20, -7.709882e-21, -1.541976e-20, 1.003089e-36, 
    0, -1.027984e-20, 1.027984e-20, 1.541976e-20, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 1.541976e-20, 
    -1.28498e-20, -7.709882e-21, 1.027984e-20, -1.798972e-20, 1.28498e-20, 
    -1.027984e-20, 5.139921e-21, -7.709882e-21, -7.709882e-21, 1.28498e-20, 
    7.709882e-21, -7.709882e-21, -1.027984e-20, 1.541976e-20, 0, 
    -1.28498e-20, 1.28498e-20, 2.055969e-20, -2.312965e-20, -2.312965e-20, 
    -5.139921e-21, 1.027984e-20, -1.027984e-20, -2.826957e-20, -1.28498e-20, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, 2.569961e-21, 
    0, 5.139921e-21, 0, -2.569961e-21, 7.709882e-21, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, 1.027984e-20, 
    7.709882e-21, 2.569961e-21, -2.312965e-20, 2.569961e-21, -1.027984e-20, 
    -7.709882e-21, 1.027984e-20, 7.709882e-21, 1.28498e-20, -7.709882e-21, 0, 
    -7.709882e-21, -7.709882e-21, -2.312965e-20, 1.541976e-20, -2.569961e-21, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 1.541976e-20, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, 2.569961e-21, 
    5.139921e-21, -1.003089e-36, 5.139921e-21, -1.28498e-20, 1.28498e-20, 
    1.027984e-20, -5.139921e-21,
  0, -7.709882e-21, 1.027984e-20, 1.003089e-36, -5.139921e-21, 1.003089e-36, 
    7.709882e-21, 7.709882e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 0, 0, 1.798972e-20, 0, -7.709882e-21, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 1.003089e-36, -2.569961e-21, 5.139921e-21, 
    -1.027984e-20, 1.003089e-36, 2.569961e-21, 2.569961e-21, -1.798972e-20, 
    -2.569961e-21, -7.709882e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, -1.003089e-36, 2.569961e-21, 5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, -1.28498e-20, -1.003089e-36, 
    -2.569961e-21, 1.027984e-20, 2.569961e-21, -5.139921e-21, 1.28498e-20, 
    5.139921e-21, 7.709882e-21, 0, -1.28498e-20, 1.003089e-36, 0, 
    -2.569961e-21, -2.569961e-21, 1.28498e-20, 1.027984e-20, 0, 
    -2.569961e-21, 0, 0, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    1.003089e-36, -7.709882e-21, 1.027984e-20, 5.139921e-21, -2.055969e-20, 
    -5.139921e-21, 0, 2.569961e-21, -7.709882e-21, -1.798972e-20, 
    -1.027984e-20, 7.709882e-21, 1.027984e-20, 2.569961e-21, -1.28498e-20, 
    -7.709882e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, 0, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, -2.569961e-21, 
    7.709882e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -5.139921e-21, -1.003089e-36, -1.28498e-20, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, 1.798972e-20, 5.139921e-21, -7.709882e-21, 5.139921e-21, 
    1.027984e-20, -7.709882e-21, 7.709882e-21, -2.569961e-21, -1.28498e-20, 
    -5.139921e-21, 7.709882e-21, 5.139921e-21, -7.709882e-21, 5.139921e-21, 
    1.027984e-20, 2.569961e-21, 7.709882e-21, -7.709882e-21, -2.569961e-21, 
    1.027984e-20, -1.28498e-20, 5.139921e-21, 0, 1.003089e-36, 7.709882e-21, 
    -1.027984e-20, -2.569961e-21, 1.28498e-20, -2.569961e-21, -1.798972e-20, 
    -1.003089e-36, -1.027984e-20, -2.569961e-21, 7.709882e-21, -1.003089e-36, 
    -1.027984e-20, 5.139921e-21, 1.003089e-36, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, 1.541976e-20, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, 7.709882e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, -1.027984e-20, 5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -1.027984e-20, 1.541976e-20, -7.709882e-21, 
    -7.709882e-21, 7.709882e-21, 0, 2.569961e-21, -7.709882e-21, 0, 
    5.139921e-21, -1.027984e-20, 1.003089e-36, 5.139921e-21, -2.569961e-21, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, 7.709882e-21, -1.027984e-20, 
    2.569961e-21, -7.709882e-21, 1.28498e-20, 2.569961e-21, 7.709882e-21, 
    -5.139921e-21, 7.709882e-21, -7.709882e-21, -7.709882e-21, 7.709882e-21, 
    1.28498e-20, 5.139921e-21, 1.003089e-36, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 1.003089e-36, -1.541976e-20, -7.709882e-21, -7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 1.027984e-20, -1.28498e-20, -1.027984e-20, 
    5.139921e-21, 1.28498e-20, -1.541976e-20, -2.569961e-21, -1.28498e-20, 
    1.027984e-20, 7.709882e-21, -7.709882e-21, 2.569961e-21, 1.541976e-20, 
    -1.027984e-20, 2.569961e-21, -2.569961e-21, 7.709882e-21, -1.003089e-36, 
    2.569961e-21, 0, 1.027984e-20, -2.569961e-21, 0, 5.139921e-21, 
    -7.709882e-21, 5.139921e-21, 1.28498e-20, -1.541976e-20, -1.541976e-20, 
    -1.798972e-20, -1.541976e-20, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    0, -2.569961e-21, -7.709882e-21, -2.569961e-21, 1.003089e-36, 
    1.28498e-20, 7.709882e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, 1.003089e-36, -7.709882e-21, 
    -5.139921e-21, 1.541976e-20, 7.709882e-21, -7.709882e-21, 1.027984e-20, 
    2.055969e-20, 0, 5.139921e-21, -5.139921e-21, 1.003089e-36, 0, 0, 
    -2.569961e-21, -2.569961e-21, 7.709882e-21, 5.139921e-21, 0, 
    7.709882e-21, 0, 2.569961e-21, -5.139921e-21, 5.139921e-21, 0, 
    5.139921e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, -2.569961e-21, 
    0, -2.569961e-21, 1.027984e-20, 2.569961e-21, -1.28498e-20, 1.003089e-36, 
    0, -2.569961e-21, -5.139921e-21, -7.709882e-21, 5.139921e-21, 
    5.139921e-21, -1.28498e-20, 1.027984e-20, -1.003089e-36, 7.709882e-21, 
    7.709882e-21, 0, 2.569961e-21, 0, 2.569961e-21, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, -1.541976e-20, 2.569961e-21, 0, 0, 
    -5.139921e-21, -5.139921e-21, 1.003089e-36, 2.569961e-21, 0, 
    -7.709882e-21, 7.709882e-21, 1.28498e-20, 1.541976e-20, -2.569961e-21, 
    -1.003089e-36, -2.569961e-21, -1.28498e-20, 7.709882e-21, 2.569961e-21, 
    7.709882e-21, -1.027984e-20, 0, -7.709882e-21, 0, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21,
  1.28498e-20, 5.139921e-21, 1.027984e-20, -2.569961e-21, -7.709882e-21, 
    7.709882e-21, 1.027984e-20, -1.003089e-36, 2.569961e-21, -1.798972e-20, 
    -5.139921e-21, -1.027984e-20, 1.003089e-36, 1.027984e-20, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, 
    -7.709882e-21, 1.003089e-36, -5.139921e-21, -1.28498e-20, 1.027984e-20, 
    2.569961e-21, 5.139921e-21, 1.798972e-20, 0, 2.312965e-20, -1.28498e-20, 
    -2.055969e-20, 7.709882e-21, 2.569961e-21, 1.027984e-20, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, -2.055969e-20, 7.709882e-21, -7.709882e-21, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, 7.709882e-21, 1.027984e-20, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, 1.003089e-36, 5.139921e-21, 
    -5.139921e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, -2.569961e-21, 
    0, 5.139921e-21, 1.027984e-20, -1.28498e-20, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -7.709882e-21, -1.003089e-36, -1.28498e-20, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 1.28498e-20, 
    -5.139921e-21, -7.709882e-21, 1.28498e-20, 1.28498e-20, -1.28498e-20, 
    1.541976e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -1.003089e-36, -5.139921e-21, 0, 7.709882e-21, -5.139921e-21, 
    1.027984e-20, -1.28498e-20, 2.569961e-21, -5.139921e-21, 0, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 1.28498e-20, -5.139921e-21, -1.003089e-36, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    0, 1.798972e-20, -2.312965e-20, 5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, 1.003089e-36, 1.003089e-36, 
    7.709882e-21, -2.569961e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, 2.569961e-21, 7.709882e-21, -1.003089e-36, 
    7.709882e-21, -7.709882e-21, 1.541976e-20, -7.709882e-21, -2.569961e-21, 
    5.139921e-21, -7.709882e-21, 5.139921e-21, -2.569961e-21, -1.541976e-20, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, 0, 0, 2.055969e-20, 
    -7.709882e-21, -7.709882e-21, -1.027984e-20, -1.798972e-20, 1.541976e-20, 
    -2.569961e-21, 5.139921e-21, 1.003089e-36, -2.569961e-21, 2.569961e-21, 
    0, 7.709882e-21, 7.709882e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, 1.027984e-20, -2.569961e-21, -1.027984e-20, -1.027984e-20, 
    2.569961e-21, 2.569961e-21, 7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -1.28498e-20, 2.569961e-21, -1.027984e-20, 
    -7.709882e-21, -5.139921e-21, -1.027984e-20, 2.569961e-21, 1.541976e-20, 
    -5.139921e-21, 1.28498e-20, 7.709882e-21, 5.139921e-21, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, 1.28498e-20, -1.798972e-20, -5.139921e-21, 
    -2.055969e-20, -1.027984e-20, -1.28498e-20, -1.541976e-20, -2.569961e-21, 
    2.569961e-21, 1.003089e-36, -1.027984e-20, 1.027984e-20, 1.798972e-20, 
    2.569961e-21, 1.28498e-20, 7.709882e-21, 1.027984e-20, 1.28498e-20, 0, 
    1.003089e-36, -1.798972e-20, 0, 2.569961e-21, 1.003089e-36, 
    -5.139921e-21, -7.709882e-21, 5.139921e-21, -5.139921e-21, -2.569961e-21, 
    5.139921e-21, 0, 1.28498e-20, -1.027984e-20, -2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    2.569961e-21, 1.28498e-20, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, -1.027984e-20, -1.027984e-20, 
    2.569961e-21, 1.541976e-20, -2.569961e-21, -1.027984e-20, -7.709882e-21, 
    1.28498e-20, -1.027984e-20, -7.709882e-21, -1.027984e-20, -7.709882e-21, 
    2.569961e-21, 2.569961e-21, 7.709882e-21, -7.709882e-21, -1.003089e-36, 
    5.139921e-21, 1.28498e-20, 7.709882e-21, 2.569961e-21, -1.541976e-20, 0, 
    -2.569961e-21, -5.139921e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, -2.312965e-20, -2.569961e-21, -1.027984e-20, -5.139921e-21, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, -2.055969e-20, 
    2.826957e-20, -1.541976e-20, -5.139921e-21, -1.003089e-36, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, 7.709882e-21, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, 7.709882e-21, 5.139921e-21, 0, 1.28498e-20, 5.139921e-21, 
    -7.709882e-21, -1.541976e-20, 0, 0, -2.569961e-21, -1.798972e-20, 
    -1.027984e-20, 1.003089e-36, 2.569961e-21, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, 1.28498e-20, 7.709882e-21, -1.541976e-20, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 1.027984e-20, -1.027984e-20, 1.28498e-20, 
    1.541976e-20, -2.569961e-21, -7.709882e-21, 2.569961e-21, -1.027984e-20,
  1.003089e-36, 1.027984e-20, -2.569961e-21, 0, 5.139921e-21, 0, 
    1.003089e-36, 5.139921e-21, -1.027984e-20, -7.709882e-21, -7.709882e-21, 
    -1.541976e-20, 1.28498e-20, 5.139921e-21, 7.709882e-21, 7.709882e-21, 
    -1.027984e-20, 1.28498e-20, -5.139921e-21, 7.709882e-21, 1.28498e-20, 
    2.569961e-21, -1.541976e-20, -1.003089e-36, 1.798972e-20, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -1.541976e-20, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, -5.139921e-21, -7.709882e-21, -1.003089e-36, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, 0, -7.709882e-21, 
    -1.28498e-20, -5.139921e-21, -1.798972e-20, 2.569961e-21, -1.798972e-20, 
    -5.139921e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, 1.28498e-20, -2.569961e-21, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, 7.709882e-21, 0, 
    -5.139921e-21, -7.709882e-21, 1.541976e-20, -1.027984e-20, -5.139921e-21, 
    -7.709882e-21, 1.027984e-20, -1.027984e-20, 1.541976e-20, 5.139921e-21, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -1.027984e-20, 2.569961e-20, 5.139921e-21, 1.027984e-20, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 1.541976e-20, 1.541976e-20, 5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    1.541976e-20, -1.541976e-20, 2.055969e-20, -1.541976e-20, -1.541976e-20, 
    7.709882e-21, 5.139921e-21, -1.541976e-20, 1.541976e-20, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    1.003089e-36, -5.139921e-21, 5.139921e-21, 0, -1.003089e-36, 
    -1.798972e-20, 1.003089e-36, -5.139921e-21, 2.569961e-21, -2.312965e-20, 
    0, 2.569961e-21, -3.083953e-20, 0, -1.28498e-20, -1.28498e-20, 
    -1.798972e-20, 7.709882e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 2.312965e-20, -5.139921e-21, 1.28498e-20, 
    1.003089e-36, -7.709882e-21, 5.139921e-21, -5.139921e-21, -1.28498e-20, 
    2.569961e-21, 7.709882e-21, 7.709882e-21, 5.139921e-21, -2.055969e-20, 
    -1.003089e-36, -1.003089e-36, -7.709882e-21, -1.027984e-20, 1.027984e-20, 
    0, 2.312965e-20, 2.569961e-21, -1.003089e-36, 0, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, -2.569961e-21, -1.541976e-20, -1.798972e-20, 
    7.709882e-21, 1.003089e-36, 7.709882e-21, -2.569961e-21, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, -1.798972e-20, 2.569961e-21, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, -1.28498e-20, -1.541976e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 5.139921e-21, -1.003089e-36, -3.340949e-20, 
    -5.139921e-21, -1.027984e-20, 0, 5.139921e-21, 0, 1.003089e-36, 
    5.139921e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, -1.003089e-36, 
    -7.709882e-21, 2.569961e-21, -1.027984e-20, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, -1.027984e-20, 7.709882e-21, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, 0, -1.027984e-20, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, 1.027984e-20, -2.569961e-21, 
    1.027984e-20, -2.569961e-21, -1.027984e-20, 1.28498e-20, -5.139921e-21, 
    1.28498e-20, 0, 2.312965e-20, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    2.569961e-21, -7.709882e-21, -1.28498e-20, -2.569961e-21, 1.027984e-20, 
    -2.569961e-20, 1.003089e-36, 1.027984e-20, 1.027984e-20, -1.28498e-20, 
    -1.28498e-20, 7.709882e-21, 7.709882e-21, 2.569961e-21, -1.027984e-20, 
    1.28498e-20, 1.003089e-36, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    -2.055969e-20, -5.139921e-21, 0, -1.541976e-20, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, -1.003089e-36, 5.139921e-21, 1.003089e-36, 
    5.139921e-21, 0, -1.003089e-36, -7.709882e-21, 1.28498e-20, 1.003089e-36, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, 1.28498e-20, -1.28498e-20, 
    1.541976e-20, 1.541976e-20, -1.28498e-20, 5.139921e-21, 7.709882e-21, 
    2.569961e-21, -1.28498e-20, -1.541976e-20, -7.709882e-21, -1.798972e-20, 
    -1.027984e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, 1.798972e-20, 
    -2.569961e-21, -2.569961e-21, 1.003089e-36, 7.709882e-21, -1.027984e-20, 
    5.139921e-21, 1.798972e-20, 1.027984e-20, -2.055969e-20, 1.798972e-20, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 
    7.709882e-21, 2.569961e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, 0, 
    -1.28498e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -7.709882e-21, 7.709882e-21, -2.569961e-21, 2.569961e-21, -2.312965e-20, 
    2.569961e-21, 2.569961e-21, -1.003089e-36, -5.139921e-21, 0, 
    2.569961e-21, 7.709882e-21, -7.709882e-21, 1.28498e-20, 5.139921e-21, 
    -7.709882e-21, -7.709882e-21, -5.139921e-21, -1.28498e-20, 0, 
    -2.569961e-21,
  7.709882e-21, 5.139921e-21, 1.003089e-36, 1.027984e-20, -7.709882e-21, 0, 
    -2.569961e-21, -1.28498e-20, -1.28498e-20, -1.027984e-20, -2.569961e-20, 
    7.709882e-21, 1.28498e-20, 3.597945e-20, 1.027984e-20, 2.569961e-21, 
    1.541976e-20, -1.541976e-20, -2.312965e-20, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 2.569961e-21, -1.027984e-20, 1.28498e-20, 
    -1.003089e-36, 7.709882e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -1.541976e-20, 0, 7.709882e-21, 2.055969e-20, 2.569961e-21, 1.28498e-20, 
    2.569961e-21, -1.28498e-20, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    7.709882e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 
    -2.312965e-20, 1.027984e-20, -2.055969e-20, -1.027984e-20, -1.541976e-20, 
    1.28498e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 2.569961e-21, 
    1.28498e-20, -1.003089e-36, -1.003089e-36, -1.28498e-20, -1.28498e-20, 
    -1.027984e-20, -1.541976e-20, 2.569961e-21, -7.709882e-21, -1.28498e-20, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 1.28498e-20, 
    -2.569961e-21, -1.28498e-20, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -1.003089e-36, 0, 1.28498e-20, 5.139921e-21, 
    -1.541976e-20, -1.28498e-20, 1.003089e-36, -7.709882e-21, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    0, -7.709882e-21, 1.28498e-20, -2.826957e-20, -7.709882e-21, 
    -1.798972e-20, 5.139921e-21, -5.139921e-21, -1.798972e-20, -1.003089e-36, 
    1.027984e-20, -1.541976e-20, 5.139921e-21, 1.798972e-20, -5.139921e-21, 
    2.569961e-21, 1.027984e-20, -1.541976e-20, -5.139921e-21, -2.569961e-21, 
    1.28498e-20, 2.569961e-21, -5.139921e-21, -2.312965e-20, -5.139921e-21, 
    0, -1.798972e-20, -1.541976e-20, -2.569961e-21, 1.798972e-20, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, 1.027984e-20, -1.003089e-36, 
    1.027984e-20, 0, -2.312965e-20, -5.139921e-21, 0, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, -7.709882e-21, 1.027984e-20, 0, 1.28498e-20, 
    2.569961e-21, -2.569961e-21, 2.312965e-20, 2.569961e-21, 1.541976e-20, 
    1.798972e-20, -2.055969e-20, -7.709882e-21, -1.798972e-20, 2.569961e-21, 
    -1.541976e-20, 1.798972e-20, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 1.798972e-20, -1.003089e-36, -1.027984e-20, 2.569961e-21, 
    -5.139921e-21, -1.28498e-20, 1.28498e-20, 7.709882e-21, -1.003089e-36, 
    1.28498e-20, 2.569961e-21, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    -1.798972e-20, -1.798972e-20, -5.139921e-21, -5.139921e-21, 0, 
    1.28498e-20, -2.569961e-21, -1.541976e-20, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 1.28498e-20, 1.28498e-20, 5.139921e-21, 1.003089e-36, 
    1.027984e-20, 1.28498e-20, 2.569961e-21, -7.709882e-21, 1.027984e-20, 
    5.139921e-21, 1.027984e-20, -1.28498e-20, 1.027984e-20, -1.798972e-20, 
    -5.139921e-21, 1.027984e-20, 7.709882e-21, -2.569961e-21, 1.027984e-20, 
    -7.709882e-21, 7.709882e-21, -5.139921e-21, 1.027984e-20, -2.312965e-20, 
    -1.28498e-20, -5.139921e-21, -1.003089e-36, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, 0, -2.569961e-21, -1.28498e-20, -2.569961e-21, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, -2.569961e-21, 1.798972e-20, 
    -2.569961e-21, -7.709882e-21, 1.541976e-20, 1.027984e-20, 7.709882e-21, 
    7.709882e-21, 1.28498e-20, -1.798972e-20, 2.569961e-21, 7.709882e-21, 
    -1.28498e-20, -2.569961e-20, -1.003089e-36, -1.28498e-20, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, 1.541976e-20, -1.003089e-36, 5.139921e-21, -1.003089e-36, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, -1.28498e-20, 
    -1.003089e-36, -1.027984e-20, 7.709882e-21, -1.541976e-20, 5.139921e-21, 
    1.541976e-20, 5.139921e-21, 1.28498e-20, 1.003089e-36, -7.709882e-21, 
    7.709882e-21, -1.541976e-20, 2.569961e-21, -1.798972e-20, -1.798972e-20, 
    -1.541976e-20, 7.709882e-21, 0, 2.055969e-20, 2.826957e-20, 
    -1.003089e-36, -2.569961e-21, 1.798972e-20, -1.003089e-36, 7.709882e-21, 
    5.139921e-21, -1.798972e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, 
    0, -1.28498e-20, 2.569961e-21, -1.541976e-20, -7.709882e-21, 
    2.569961e-21, -1.28498e-20, -2.826957e-20, 2.569961e-21, -7.709882e-21, 
    -2.569961e-21, -1.798972e-20, 5.139921e-21, 7.709882e-21, -1.027984e-20, 
    -2.826957e-20, 5.139921e-21, 7.709882e-21, 7.709882e-21, 1.28498e-20, 
    -7.709882e-21, 7.709882e-21, 1.541976e-20, -1.541976e-20, -5.139921e-21, 
    3.009266e-36, -2.569961e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, 2.055969e-20, -7.709882e-21, -7.709882e-21, 
    -1.28498e-20, 0, -5.139921e-21, 2.569961e-21, 1.003089e-36, 1.541976e-20, 
    5.139921e-21, -2.569961e-21, -2.055969e-20, 7.709882e-21, 2.569961e-21, 
    2.055969e-20, 1.027984e-20, -7.709882e-21, -1.541976e-20, 2.055969e-20, 
    -1.798972e-20, 7.709882e-21, 1.027984e-20, 2.569961e-21, -1.541976e-20, 
    1.003089e-36, 1.28498e-20, -1.541976e-20,
  6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.153676e-12, 5.176412e-12, 5.171992e-12, 5.19033e-12, 5.180158e-12, 
    5.192165e-12, 5.158286e-12, 5.177314e-12, 5.165167e-12, 5.155724e-12, 
    5.225918e-12, 5.191148e-12, 5.262042e-12, 5.239865e-12, 5.29558e-12, 
    5.25859e-12, 5.303038e-12, 5.294514e-12, 5.320175e-12, 5.312823e-12, 
    5.345644e-12, 5.323568e-12, 5.362661e-12, 5.340373e-12, 5.343859e-12, 
    5.322839e-12, 5.198146e-12, 5.221588e-12, 5.196757e-12, 5.2001e-12, 
    5.1986e-12, 5.180368e-12, 5.171179e-12, 5.151939e-12, 5.155433e-12, 
    5.169564e-12, 5.201603e-12, 5.190728e-12, 5.218139e-12, 5.21752e-12, 
    5.248038e-12, 5.234278e-12, 5.285576e-12, 5.270996e-12, 5.31313e-12, 
    5.302533e-12, 5.312632e-12, 5.30957e-12, 5.312672e-12, 5.297131e-12, 
    5.303789e-12, 5.290114e-12, 5.236855e-12, 5.252506e-12, 5.205827e-12, 
    5.177759e-12, 5.159121e-12, 5.145894e-12, 5.147763e-12, 5.151328e-12, 
    5.169646e-12, 5.186871e-12, 5.199998e-12, 5.208779e-12, 5.217431e-12, 
    5.243618e-12, 5.257482e-12, 5.288524e-12, 5.282923e-12, 5.292412e-12, 
    5.301479e-12, 5.316701e-12, 5.314196e-12, 5.320902e-12, 5.292163e-12, 
    5.311262e-12, 5.279732e-12, 5.288355e-12, 5.219779e-12, 5.193662e-12, 
    5.182558e-12, 5.172842e-12, 5.149201e-12, 5.165526e-12, 5.159091e-12, 
    5.174403e-12, 5.184132e-12, 5.17932e-12, 5.209019e-12, 5.197473e-12, 
    5.258304e-12, 5.232101e-12, 5.300422e-12, 5.284072e-12, 5.30434e-12, 
    5.293998e-12, 5.311719e-12, 5.29577e-12, 5.323398e-12, 5.329414e-12, 
    5.325303e-12, 5.341097e-12, 5.294886e-12, 5.312632e-12, 5.179185e-12, 
    5.17997e-12, 5.183626e-12, 5.167554e-12, 5.166571e-12, 5.151843e-12, 
    5.164948e-12, 5.170529e-12, 5.184696e-12, 5.193076e-12, 5.201042e-12, 
    5.218557e-12, 5.238119e-12, 5.265476e-12, 5.285132e-12, 5.298307e-12, 
    5.290229e-12, 5.297361e-12, 5.289388e-12, 5.285651e-12, 5.32716e-12, 
    5.303851e-12, 5.338825e-12, 5.33689e-12, 5.321062e-12, 5.337108e-12, 
    5.180521e-12, 5.176005e-12, 5.160325e-12, 5.172596e-12, 5.15024e-12, 
    5.162753e-12, 5.169948e-12, 5.197713e-12, 5.203814e-12, 5.209471e-12, 
    5.220644e-12, 5.234982e-12, 5.260137e-12, 5.282024e-12, 5.302007e-12, 
    5.300543e-12, 5.301058e-12, 5.305522e-12, 5.294465e-12, 5.307337e-12, 
    5.309497e-12, 5.303849e-12, 5.336631e-12, 5.327265e-12, 5.336849e-12, 
    5.330751e-12, 5.177473e-12, 5.185072e-12, 5.180965e-12, 5.188687e-12, 
    5.183247e-12, 5.207436e-12, 5.214689e-12, 5.248628e-12, 5.2347e-12, 
    5.256868e-12, 5.236952e-12, 5.24048e-12, 5.257589e-12, 5.238028e-12, 
    5.280817e-12, 5.251806e-12, 5.305695e-12, 5.276722e-12, 5.307511e-12, 
    5.30192e-12, 5.311177e-12, 5.319467e-12, 5.329897e-12, 5.349142e-12, 
    5.344686e-12, 5.360781e-12, 5.196401e-12, 5.206257e-12, 5.20539e-12, 
    5.215705e-12, 5.223334e-12, 5.239871e-12, 5.266393e-12, 5.256419e-12, 
    5.27473e-12, 5.278406e-12, 5.250588e-12, 5.267667e-12, 5.212854e-12, 
    5.221709e-12, 5.216437e-12, 5.197178e-12, 5.258717e-12, 5.227133e-12, 
    5.285457e-12, 5.268346e-12, 5.318285e-12, 5.293448e-12, 5.342232e-12, 
    5.363087e-12, 5.382719e-12, 5.405658e-12, 5.211637e-12, 5.20494e-12, 
    5.216932e-12, 5.233524e-12, 5.248921e-12, 5.269389e-12, 5.271484e-12, 
    5.275319e-12, 5.285252e-12, 5.293604e-12, 5.276531e-12, 5.295697e-12, 
    5.223761e-12, 5.261458e-12, 5.202408e-12, 5.220187e-12, 5.232546e-12, 
    5.227125e-12, 5.25528e-12, 5.261915e-12, 5.288881e-12, 5.274942e-12, 
    5.357939e-12, 5.321217e-12, 5.423127e-12, 5.394645e-12, 5.2026e-12, 
    5.211615e-12, 5.242989e-12, 5.228061e-12, 5.270756e-12, 5.281266e-12, 
    5.28981e-12, 5.300732e-12, 5.301911e-12, 5.308382e-12, 5.297778e-12, 
    5.307964e-12, 5.269433e-12, 5.286651e-12, 5.239404e-12, 5.250903e-12, 
    5.245613e-12, 5.23981e-12, 5.257719e-12, 5.276799e-12, 5.277208e-12, 
    5.283326e-12, 5.300564e-12, 5.27093e-12, 5.362676e-12, 5.306012e-12, 
    5.221445e-12, 5.238808e-12, 5.241289e-12, 5.234563e-12, 5.280212e-12, 
    5.263671e-12, 5.308225e-12, 5.296183e-12, 5.315913e-12, 5.306109e-12, 
    5.304666e-12, 5.292075e-12, 5.284235e-12, 5.26443e-12, 5.248315e-12, 
    5.235539e-12, 5.23851e-12, 5.252545e-12, 5.277966e-12, 5.302018e-12, 
    5.296749e-12, 5.314414e-12, 5.26766e-12, 5.287264e-12, 5.279686e-12, 
    5.299444e-12, 5.256154e-12, 5.293014e-12, 5.246732e-12, 5.25079e-12, 
    5.263343e-12, 5.288592e-12, 5.294181e-12, 5.300146e-12, 5.296465e-12, 
    5.278612e-12, 5.275687e-12, 5.263038e-12, 5.259545e-12, 5.249907e-12, 
    5.241927e-12, 5.249218e-12, 5.256874e-12, 5.27862e-12, 5.298217e-12, 
    5.319585e-12, 5.324814e-12, 5.349779e-12, 5.329455e-12, 5.362992e-12, 
    5.334477e-12, 5.383841e-12, 5.295152e-12, 5.333641e-12, 5.263914e-12, 
    5.271426e-12, 5.285012e-12, 5.316174e-12, 5.299352e-12, 5.319026e-12, 
    5.275573e-12, 5.253028e-12, 5.247197e-12, 5.236315e-12, 5.247446e-12, 
    5.246541e-12, 5.257192e-12, 5.253769e-12, 5.279342e-12, 5.265605e-12, 
    5.30463e-12, 5.318871e-12, 5.359093e-12, 5.383752e-12, 5.408856e-12, 
    5.419938e-12, 5.423312e-12, 5.424722e-12 ;

 SOIL3N_vr =
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.117974e-11, 3.131729e-11, 3.129055e-11, 3.14015e-11, 3.133995e-11, 
    3.14126e-11, 3.120763e-11, 3.132275e-11, 3.124926e-11, 3.119213e-11, 
    3.16168e-11, 3.140645e-11, 3.183535e-11, 3.170118e-11, 3.203825e-11, 
    3.181447e-11, 3.208338e-11, 3.203181e-11, 3.218706e-11, 3.214258e-11, 
    3.234115e-11, 3.220759e-11, 3.24441e-11, 3.230926e-11, 3.233035e-11, 
    3.220318e-11, 3.144878e-11, 3.159061e-11, 3.144038e-11, 3.14606e-11, 
    3.145153e-11, 3.134122e-11, 3.128563e-11, 3.116923e-11, 3.119037e-11, 
    3.127586e-11, 3.14697e-11, 3.14039e-11, 3.156974e-11, 3.1566e-11, 
    3.175063e-11, 3.166738e-11, 3.197773e-11, 3.188953e-11, 3.214444e-11, 
    3.208033e-11, 3.214142e-11, 3.21229e-11, 3.214166e-11, 3.204764e-11, 
    3.208793e-11, 3.200519e-11, 3.168297e-11, 3.177766e-11, 3.149525e-11, 
    3.132544e-11, 3.121268e-11, 3.113266e-11, 3.114397e-11, 3.116553e-11, 
    3.127636e-11, 3.138057e-11, 3.145999e-11, 3.151311e-11, 3.156546e-11, 
    3.172389e-11, 3.180777e-11, 3.199557e-11, 3.196168e-11, 3.201909e-11, 
    3.207395e-11, 3.216604e-11, 3.215089e-11, 3.219146e-11, 3.201758e-11, 
    3.213314e-11, 3.194238e-11, 3.199455e-11, 3.157967e-11, 3.142165e-11, 
    3.135447e-11, 3.129569e-11, 3.115267e-11, 3.125144e-11, 3.12125e-11, 
    3.130514e-11, 3.1364e-11, 3.133489e-11, 3.151457e-11, 3.144471e-11, 
    3.181274e-11, 3.165421e-11, 3.206755e-11, 3.196864e-11, 3.209126e-11, 
    3.202869e-11, 3.21359e-11, 3.203941e-11, 3.220656e-11, 3.224296e-11, 
    3.221809e-11, 3.231363e-11, 3.203406e-11, 3.214142e-11, 3.133407e-11, 
    3.133882e-11, 3.136094e-11, 3.12637e-11, 3.125775e-11, 3.116865e-11, 
    3.124793e-11, 3.12817e-11, 3.136741e-11, 3.141811e-11, 3.146631e-11, 
    3.157227e-11, 3.169062e-11, 3.185613e-11, 3.197505e-11, 3.205476e-11, 
    3.200588e-11, 3.204903e-11, 3.200079e-11, 3.197819e-11, 3.222932e-11, 
    3.20883e-11, 3.229989e-11, 3.228819e-11, 3.219242e-11, 3.22895e-11, 
    3.134215e-11, 3.131483e-11, 3.121996e-11, 3.12942e-11, 3.115895e-11, 
    3.123465e-11, 3.127818e-11, 3.144616e-11, 3.148308e-11, 3.15173e-11, 
    3.158489e-11, 3.167164e-11, 3.182382e-11, 3.195625e-11, 3.207714e-11, 
    3.206828e-11, 3.20714e-11, 3.209841e-11, 3.203151e-11, 3.210939e-11, 
    3.212246e-11, 3.208829e-11, 3.228662e-11, 3.222995e-11, 3.228794e-11, 
    3.225104e-11, 3.132371e-11, 3.136968e-11, 3.134484e-11, 3.139156e-11, 
    3.135864e-11, 3.150499e-11, 3.154887e-11, 3.17542e-11, 3.166993e-11, 
    3.180405e-11, 3.168356e-11, 3.170491e-11, 3.180841e-11, 3.169007e-11, 
    3.194894e-11, 3.177342e-11, 3.209946e-11, 3.192417e-11, 3.211044e-11, 
    3.207662e-11, 3.213262e-11, 3.218277e-11, 3.224588e-11, 3.236231e-11, 
    3.233535e-11, 3.243272e-11, 3.143823e-11, 3.149786e-11, 3.149261e-11, 
    3.155502e-11, 3.160117e-11, 3.170122e-11, 3.186168e-11, 3.180134e-11, 
    3.191212e-11, 3.193436e-11, 3.176606e-11, 3.186939e-11, 3.153777e-11, 
    3.159134e-11, 3.155945e-11, 3.144293e-11, 3.181523e-11, 3.162416e-11, 
    3.197701e-11, 3.187349e-11, 3.217562e-11, 3.202536e-11, 3.232051e-11, 
    3.244667e-11, 3.256545e-11, 3.270423e-11, 3.15304e-11, 3.148989e-11, 
    3.156244e-11, 3.166282e-11, 3.175597e-11, 3.18798e-11, 3.189248e-11, 
    3.191568e-11, 3.197578e-11, 3.202631e-11, 3.192301e-11, 3.203897e-11, 
    3.160375e-11, 3.183183e-11, 3.147456e-11, 3.158213e-11, 3.16569e-11, 
    3.162411e-11, 3.179444e-11, 3.183459e-11, 3.199773e-11, 3.19134e-11, 
    3.241553e-11, 3.219336e-11, 3.280992e-11, 3.26376e-11, 3.147573e-11, 
    3.153027e-11, 3.172008e-11, 3.162977e-11, 3.188808e-11, 3.195166e-11, 
    3.200335e-11, 3.206943e-11, 3.207656e-11, 3.211571e-11, 3.205156e-11, 
    3.211318e-11, 3.188007e-11, 3.198424e-11, 3.169839e-11, 3.176796e-11, 
    3.173596e-11, 3.170085e-11, 3.18092e-11, 3.192463e-11, 3.192711e-11, 
    3.196412e-11, 3.206841e-11, 3.188912e-11, 3.244419e-11, 3.210137e-11, 
    3.158974e-11, 3.169479e-11, 3.17098e-11, 3.16691e-11, 3.194528e-11, 
    3.184521e-11, 3.211476e-11, 3.204191e-11, 3.216127e-11, 3.210196e-11, 
    3.209323e-11, 3.201705e-11, 3.196962e-11, 3.18498e-11, 3.175231e-11, 
    3.167501e-11, 3.169298e-11, 3.17779e-11, 3.19317e-11, 3.207721e-11, 
    3.204533e-11, 3.21522e-11, 3.186934e-11, 3.198795e-11, 3.194211e-11, 
    3.206164e-11, 3.179973e-11, 3.202274e-11, 3.174273e-11, 3.176728e-11, 
    3.184322e-11, 3.199599e-11, 3.20298e-11, 3.206588e-11, 3.204361e-11, 
    3.19356e-11, 3.191791e-11, 3.184138e-11, 3.182025e-11, 3.176194e-11, 
    3.171366e-11, 3.175777e-11, 3.180409e-11, 3.193565e-11, 3.205421e-11, 
    3.218349e-11, 3.221513e-11, 3.236616e-11, 3.22432e-11, 3.24461e-11, 
    3.227359e-11, 3.257224e-11, 3.203567e-11, 3.226852e-11, 3.184668e-11, 
    3.189213e-11, 3.197432e-11, 3.216286e-11, 3.206108e-11, 3.218011e-11, 
    3.191722e-11, 3.178082e-11, 3.174554e-11, 3.167971e-11, 3.174705e-11, 
    3.174157e-11, 3.180601e-11, 3.17853e-11, 3.194002e-11, 3.185691e-11, 
    3.209301e-11, 3.217917e-11, 3.242252e-11, 3.25717e-11, 3.272358e-11, 
    3.279063e-11, 3.281104e-11, 3.281957e-11 ;

 SOILC =
  17.34481, 17.34479, 17.3448, 17.34479, 17.34479, 17.34479, 17.3448, 
    17.34479, 17.3448, 17.34481, 17.34476, 17.34479, 17.34474, 17.34476, 
    17.34472, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34475, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.34479, 
    17.3448, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34471, 17.34472, 17.34471, 17.34473, 17.34472, 17.34473, 
    17.34473, 17.34477, 17.34478, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.3448, 17.3448, 17.34479, 17.34479, 17.34477, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34472, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.34479, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34478, 17.34478, 17.34477, 17.34476, 17.34474, 17.34473, 
    17.34472, 17.34473, 17.34472, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.34479, 17.3448, 
    17.3448, 17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34477, 
    17.34477, 17.34476, 17.34475, 17.34473, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 
    17.3447, 17.34471, 17.34479, 17.34479, 17.34479, 17.34479, 17.34479, 
    17.34478, 17.34477, 17.34475, 17.34476, 17.34475, 17.34476, 17.34476, 
    17.34475, 17.34476, 17.34473, 17.34475, 17.34472, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34471, 17.34471, 17.34469, 17.3447, 17.34469, 
    17.34478, 17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 
    17.34475, 17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 
    17.34477, 17.34478, 17.34475, 17.34476, 17.34473, 17.34474, 17.34471, 
    17.34473, 17.3447, 17.34469, 17.34468, 17.34466, 17.34477, 17.34478, 
    17.34477, 17.34476, 17.34475, 17.34474, 17.34474, 17.34474, 17.34473, 
    17.34473, 17.34474, 17.34472, 17.34477, 17.34475, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 
    17.34471, 17.34465, 17.34467, 17.34478, 17.34477, 17.34476, 17.34476, 
    17.34474, 17.34473, 17.34473, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34474, 17.34473, 17.34476, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 
    17.34472, 17.34477, 17.34476, 17.34476, 17.34476, 17.34473, 17.34474, 
    17.34472, 17.34472, 17.34471, 17.34472, 17.34472, 17.34473, 17.34473, 
    17.34474, 17.34475, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34474, 17.34473, 17.34473, 17.34472, 17.34475, 
    17.34473, 17.34475, 17.34475, 17.34474, 17.34473, 17.34473, 17.34472, 
    17.34472, 17.34473, 17.34474, 17.34474, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34475, 17.34473, 17.34472, 17.34471, 17.34471, 17.34469, 
    17.34471, 17.34469, 17.3447, 17.34468, 17.34472, 17.3447, 17.34474, 
    17.34474, 17.34473, 17.34471, 17.34472, 17.34471, 17.34474, 17.34475, 
    17.34475, 17.34476, 17.34475, 17.34475, 17.34475, 17.34475, 17.34473, 
    17.34474, 17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34465, 
    17.34465, 17.34465 ;

 SOILC_HR =
  6.195739e-08, 6.223058e-08, 6.217748e-08, 6.239782e-08, 6.22756e-08, 
    6.241988e-08, 6.201279e-08, 6.224143e-08, 6.209547e-08, 6.198199e-08, 
    6.282544e-08, 6.240766e-08, 6.325951e-08, 6.299303e-08, 6.36625e-08, 
    6.321804e-08, 6.375213e-08, 6.364969e-08, 6.395803e-08, 6.38697e-08, 
    6.426407e-08, 6.39988e-08, 6.446854e-08, 6.420073e-08, 6.424262e-08, 
    6.399005e-08, 6.249174e-08, 6.277342e-08, 6.247505e-08, 6.251522e-08, 
    6.24972e-08, 6.227812e-08, 6.216771e-08, 6.193653e-08, 6.19785e-08, 
    6.21483e-08, 6.253328e-08, 6.240261e-08, 6.273198e-08, 6.272454e-08, 
    6.309124e-08, 6.29259e-08, 6.354229e-08, 6.33671e-08, 6.387339e-08, 
    6.374605e-08, 6.38674e-08, 6.38306e-08, 6.386788e-08, 6.368114e-08, 
    6.376114e-08, 6.359683e-08, 6.295686e-08, 6.314493e-08, 6.258403e-08, 
    6.224678e-08, 6.202281e-08, 6.186388e-08, 6.188635e-08, 6.192918e-08, 
    6.21493e-08, 6.235626e-08, 6.2514e-08, 6.261951e-08, 6.272347e-08, 
    6.303814e-08, 6.320472e-08, 6.357771e-08, 6.351041e-08, 6.362443e-08, 
    6.373339e-08, 6.39163e-08, 6.388619e-08, 6.396677e-08, 6.362144e-08, 
    6.385094e-08, 6.347207e-08, 6.357569e-08, 6.275169e-08, 6.243786e-08, 
    6.230444e-08, 6.218769e-08, 6.190362e-08, 6.209979e-08, 6.202245e-08, 
    6.220644e-08, 6.232334e-08, 6.226553e-08, 6.262239e-08, 6.248365e-08, 
    6.321459e-08, 6.289974e-08, 6.372068e-08, 6.352423e-08, 6.376777e-08, 
    6.36435e-08, 6.385643e-08, 6.366479e-08, 6.399677e-08, 6.406906e-08, 
    6.401966e-08, 6.420943e-08, 6.365416e-08, 6.38674e-08, 6.226391e-08, 
    6.227334e-08, 6.231727e-08, 6.212414e-08, 6.211233e-08, 6.193537e-08, 
    6.209284e-08, 6.215989e-08, 6.233013e-08, 6.243081e-08, 6.252654e-08, 
    6.273701e-08, 6.297206e-08, 6.330077e-08, 6.353696e-08, 6.369527e-08, 
    6.35982e-08, 6.368391e-08, 6.35881e-08, 6.354319e-08, 6.404196e-08, 
    6.376189e-08, 6.418213e-08, 6.415888e-08, 6.396869e-08, 6.41615e-08, 
    6.227996e-08, 6.222569e-08, 6.203729e-08, 6.218473e-08, 6.19161e-08, 
    6.206646e-08, 6.215291e-08, 6.248654e-08, 6.255986e-08, 6.262782e-08, 
    6.276207e-08, 6.293436e-08, 6.323661e-08, 6.349962e-08, 6.373973e-08, 
    6.372213e-08, 6.372833e-08, 6.378196e-08, 6.36491e-08, 6.380377e-08, 
    6.382973e-08, 6.376186e-08, 6.415576e-08, 6.404323e-08, 6.415839e-08, 
    6.408511e-08, 6.224334e-08, 6.233464e-08, 6.22853e-08, 6.237808e-08, 
    6.231271e-08, 6.260337e-08, 6.269052e-08, 6.309833e-08, 6.293097e-08, 
    6.319734e-08, 6.295803e-08, 6.300043e-08, 6.320601e-08, 6.297097e-08, 
    6.348511e-08, 6.313651e-08, 6.378404e-08, 6.343591e-08, 6.380586e-08, 
    6.373869e-08, 6.384992e-08, 6.394953e-08, 6.407485e-08, 6.43061e-08, 
    6.425255e-08, 6.444595e-08, 6.247078e-08, 6.25892e-08, 6.257878e-08, 
    6.270273e-08, 6.27944e-08, 6.29931e-08, 6.331179e-08, 6.319195e-08, 
    6.341197e-08, 6.345614e-08, 6.312188e-08, 6.33271e-08, 6.266848e-08, 
    6.277487e-08, 6.271153e-08, 6.248011e-08, 6.321955e-08, 6.284005e-08, 
    6.354086e-08, 6.333526e-08, 6.393532e-08, 6.363688e-08, 6.422307e-08, 
    6.447366e-08, 6.470955e-08, 6.498519e-08, 6.265385e-08, 6.257338e-08, 
    6.271748e-08, 6.291684e-08, 6.310184e-08, 6.33478e-08, 6.337297e-08, 
    6.341904e-08, 6.35384e-08, 6.363876e-08, 6.34336e-08, 6.366392e-08, 
    6.279953e-08, 6.32525e-08, 6.254295e-08, 6.275658e-08, 6.290509e-08, 
    6.283995e-08, 6.317826e-08, 6.325799e-08, 6.358201e-08, 6.341452e-08, 
    6.44118e-08, 6.397055e-08, 6.51951e-08, 6.485286e-08, 6.254526e-08, 
    6.265358e-08, 6.303058e-08, 6.28512e-08, 6.336422e-08, 6.34905e-08, 
    6.359317e-08, 6.37244e-08, 6.373858e-08, 6.381633e-08, 6.368892e-08, 
    6.38113e-08, 6.334832e-08, 6.355521e-08, 6.298749e-08, 6.312566e-08, 
    6.30621e-08, 6.299238e-08, 6.320757e-08, 6.343683e-08, 6.344175e-08, 
    6.351525e-08, 6.372239e-08, 6.33663e-08, 6.446873e-08, 6.378785e-08, 
    6.27717e-08, 6.298033e-08, 6.301015e-08, 6.292932e-08, 6.347784e-08, 
    6.327909e-08, 6.381444e-08, 6.366975e-08, 6.390682e-08, 6.378902e-08, 
    6.377169e-08, 6.362038e-08, 6.352618e-08, 6.32882e-08, 6.309457e-08, 
    6.294105e-08, 6.297675e-08, 6.314539e-08, 6.345086e-08, 6.373985e-08, 
    6.367654e-08, 6.388881e-08, 6.332702e-08, 6.356257e-08, 6.347153e-08, 
    6.370894e-08, 6.318876e-08, 6.363167e-08, 6.307555e-08, 6.312431e-08, 
    6.327515e-08, 6.357854e-08, 6.364569e-08, 6.371736e-08, 6.367314e-08, 
    6.345861e-08, 6.342348e-08, 6.327148e-08, 6.322951e-08, 6.31137e-08, 
    6.301781e-08, 6.310542e-08, 6.319741e-08, 6.345871e-08, 6.369419e-08, 
    6.395094e-08, 6.401378e-08, 6.431375e-08, 6.406955e-08, 6.447252e-08, 
    6.412989e-08, 6.472303e-08, 6.365737e-08, 6.411983e-08, 6.328201e-08, 
    6.337227e-08, 6.353551e-08, 6.390996e-08, 6.370782e-08, 6.394423e-08, 
    6.34221e-08, 6.315121e-08, 6.308114e-08, 6.295038e-08, 6.308413e-08, 
    6.307325e-08, 6.320123e-08, 6.316011e-08, 6.346739e-08, 6.330233e-08, 
    6.377125e-08, 6.394237e-08, 6.442568e-08, 6.472197e-08, 6.502361e-08, 
    6.515678e-08, 6.519732e-08, 6.521426e-08 ;

 SOILC_LOSS =
  6.195739e-08, 6.223058e-08, 6.217748e-08, 6.239782e-08, 6.22756e-08, 
    6.241988e-08, 6.201279e-08, 6.224143e-08, 6.209547e-08, 6.198199e-08, 
    6.282544e-08, 6.240766e-08, 6.325951e-08, 6.299303e-08, 6.36625e-08, 
    6.321804e-08, 6.375213e-08, 6.364969e-08, 6.395803e-08, 6.38697e-08, 
    6.426407e-08, 6.39988e-08, 6.446854e-08, 6.420073e-08, 6.424262e-08, 
    6.399005e-08, 6.249174e-08, 6.277342e-08, 6.247505e-08, 6.251522e-08, 
    6.24972e-08, 6.227812e-08, 6.216771e-08, 6.193653e-08, 6.19785e-08, 
    6.21483e-08, 6.253328e-08, 6.240261e-08, 6.273198e-08, 6.272454e-08, 
    6.309124e-08, 6.29259e-08, 6.354229e-08, 6.33671e-08, 6.387339e-08, 
    6.374605e-08, 6.38674e-08, 6.38306e-08, 6.386788e-08, 6.368114e-08, 
    6.376114e-08, 6.359683e-08, 6.295686e-08, 6.314493e-08, 6.258403e-08, 
    6.224678e-08, 6.202281e-08, 6.186388e-08, 6.188635e-08, 6.192918e-08, 
    6.21493e-08, 6.235626e-08, 6.2514e-08, 6.261951e-08, 6.272347e-08, 
    6.303814e-08, 6.320472e-08, 6.357771e-08, 6.351041e-08, 6.362443e-08, 
    6.373339e-08, 6.39163e-08, 6.388619e-08, 6.396677e-08, 6.362144e-08, 
    6.385094e-08, 6.347207e-08, 6.357569e-08, 6.275169e-08, 6.243786e-08, 
    6.230444e-08, 6.218769e-08, 6.190362e-08, 6.209979e-08, 6.202245e-08, 
    6.220644e-08, 6.232334e-08, 6.226553e-08, 6.262239e-08, 6.248365e-08, 
    6.321459e-08, 6.289974e-08, 6.372068e-08, 6.352423e-08, 6.376777e-08, 
    6.36435e-08, 6.385643e-08, 6.366479e-08, 6.399677e-08, 6.406906e-08, 
    6.401966e-08, 6.420943e-08, 6.365416e-08, 6.38674e-08, 6.226391e-08, 
    6.227334e-08, 6.231727e-08, 6.212414e-08, 6.211233e-08, 6.193537e-08, 
    6.209284e-08, 6.215989e-08, 6.233013e-08, 6.243081e-08, 6.252654e-08, 
    6.273701e-08, 6.297206e-08, 6.330077e-08, 6.353696e-08, 6.369527e-08, 
    6.35982e-08, 6.368391e-08, 6.35881e-08, 6.354319e-08, 6.404196e-08, 
    6.376189e-08, 6.418213e-08, 6.415888e-08, 6.396869e-08, 6.41615e-08, 
    6.227996e-08, 6.222569e-08, 6.203729e-08, 6.218473e-08, 6.19161e-08, 
    6.206646e-08, 6.215291e-08, 6.248654e-08, 6.255986e-08, 6.262782e-08, 
    6.276207e-08, 6.293436e-08, 6.323661e-08, 6.349962e-08, 6.373973e-08, 
    6.372213e-08, 6.372833e-08, 6.378196e-08, 6.36491e-08, 6.380377e-08, 
    6.382973e-08, 6.376186e-08, 6.415576e-08, 6.404323e-08, 6.415839e-08, 
    6.408511e-08, 6.224334e-08, 6.233464e-08, 6.22853e-08, 6.237808e-08, 
    6.231271e-08, 6.260337e-08, 6.269052e-08, 6.309833e-08, 6.293097e-08, 
    6.319734e-08, 6.295803e-08, 6.300043e-08, 6.320601e-08, 6.297097e-08, 
    6.348511e-08, 6.313651e-08, 6.378404e-08, 6.343591e-08, 6.380586e-08, 
    6.373869e-08, 6.384992e-08, 6.394953e-08, 6.407485e-08, 6.43061e-08, 
    6.425255e-08, 6.444595e-08, 6.247078e-08, 6.25892e-08, 6.257878e-08, 
    6.270273e-08, 6.27944e-08, 6.29931e-08, 6.331179e-08, 6.319195e-08, 
    6.341197e-08, 6.345614e-08, 6.312188e-08, 6.33271e-08, 6.266848e-08, 
    6.277487e-08, 6.271153e-08, 6.248011e-08, 6.321955e-08, 6.284005e-08, 
    6.354086e-08, 6.333526e-08, 6.393532e-08, 6.363688e-08, 6.422307e-08, 
    6.447366e-08, 6.470955e-08, 6.498519e-08, 6.265385e-08, 6.257338e-08, 
    6.271748e-08, 6.291684e-08, 6.310184e-08, 6.33478e-08, 6.337297e-08, 
    6.341904e-08, 6.35384e-08, 6.363876e-08, 6.34336e-08, 6.366392e-08, 
    6.279953e-08, 6.32525e-08, 6.254295e-08, 6.275658e-08, 6.290509e-08, 
    6.283995e-08, 6.317826e-08, 6.325799e-08, 6.358201e-08, 6.341452e-08, 
    6.44118e-08, 6.397055e-08, 6.51951e-08, 6.485286e-08, 6.254526e-08, 
    6.265358e-08, 6.303058e-08, 6.28512e-08, 6.336422e-08, 6.34905e-08, 
    6.359317e-08, 6.37244e-08, 6.373858e-08, 6.381633e-08, 6.368892e-08, 
    6.38113e-08, 6.334832e-08, 6.355521e-08, 6.298749e-08, 6.312566e-08, 
    6.30621e-08, 6.299238e-08, 6.320757e-08, 6.343683e-08, 6.344175e-08, 
    6.351525e-08, 6.372239e-08, 6.33663e-08, 6.446873e-08, 6.378785e-08, 
    6.27717e-08, 6.298033e-08, 6.301015e-08, 6.292932e-08, 6.347784e-08, 
    6.327909e-08, 6.381444e-08, 6.366975e-08, 6.390682e-08, 6.378902e-08, 
    6.377169e-08, 6.362038e-08, 6.352618e-08, 6.32882e-08, 6.309457e-08, 
    6.294105e-08, 6.297675e-08, 6.314539e-08, 6.345086e-08, 6.373985e-08, 
    6.367654e-08, 6.388881e-08, 6.332702e-08, 6.356257e-08, 6.347153e-08, 
    6.370894e-08, 6.318876e-08, 6.363167e-08, 6.307555e-08, 6.312431e-08, 
    6.327515e-08, 6.357854e-08, 6.364569e-08, 6.371736e-08, 6.367314e-08, 
    6.345861e-08, 6.342348e-08, 6.327148e-08, 6.322951e-08, 6.31137e-08, 
    6.301781e-08, 6.310542e-08, 6.319741e-08, 6.345871e-08, 6.369419e-08, 
    6.395094e-08, 6.401378e-08, 6.431375e-08, 6.406955e-08, 6.447252e-08, 
    6.412989e-08, 6.472303e-08, 6.365737e-08, 6.411983e-08, 6.328201e-08, 
    6.337227e-08, 6.353551e-08, 6.390996e-08, 6.370782e-08, 6.394423e-08, 
    6.34221e-08, 6.315121e-08, 6.308114e-08, 6.295038e-08, 6.308413e-08, 
    6.307325e-08, 6.320123e-08, 6.316011e-08, 6.346739e-08, 6.330233e-08, 
    6.377125e-08, 6.394237e-08, 6.442568e-08, 6.472197e-08, 6.502361e-08, 
    6.515678e-08, 6.519732e-08, 6.521426e-08 ;

 SOILICE =
  96.04986, 96.50368, 96.41534, 96.78214, 96.57854, 96.81889, 96.14174, 
    96.52174, 96.27904, 96.09063, 97.49641, 96.79852, 98.22427, 97.77689, 
    98.90291, 98.1546, 99.05418, 98.88121, 99.40219, 99.25278, 99.92099, 
    99.4712, 100.2683, 99.81343, 99.88454, 99.45639, 96.93867, 97.40939, 
    96.91084, 96.97787, 96.94778, 96.58277, 96.39918, 96.01519, 96.08482, 
    96.36686, 97.00801, 96.79005, 97.33982, 97.32738, 97.9416, 97.66438, 
    98.70012, 98.40508, 99.25901, 99.04386, 99.24891, 99.1867, 99.24972, 
    98.93429, 99.06937, 98.79205, 97.71628, 98.03174, 97.09269, 96.53072, 
    96.15839, 95.89476, 95.932, 96.00304, 96.36852, 96.71285, 96.97577, 
    97.15189, 97.32559, 97.85267, 98.13219, 98.75986, 98.64637, 98.83865, 
    99.02247, 99.3316, 99.28068, 99.41702, 98.83353, 99.22112, 98.58176, 
    98.7564, 97.37305, 96.84882, 96.62666, 96.43233, 95.96065, 96.28624, 
    96.15781, 96.46348, 96.65803, 96.56177, 97.15671, 96.92516, 98.14877, 
    97.62061, 99.00102, 98.66965, 99.08053, 98.87074, 99.23038, 98.90667, 
    99.46777, 99.59022, 99.50654, 99.82814, 98.88875, 99.24892, 96.55908, 
    96.57478, 96.6479, 96.32672, 96.30708, 96.01329, 96.27467, 96.38611, 
    96.6693, 96.83707, 96.99671, 97.34825, 97.74178, 98.29359, 98.69112, 
    98.95812, 98.79433, 98.93893, 98.77731, 98.7016, 99.54434, 99.07063, 
    99.78185, 99.74241, 99.42027, 99.74685, 96.5858, 96.49549, 96.18242, 
    96.42738, 95.98132, 96.23087, 96.37455, 96.93004, 97.05229, 97.16579, 
    97.39015, 97.67857, 98.18573, 98.62823, 99.03316, 99.00346, 99.01392, 
    99.10452, 98.88021, 99.14137, 99.18526, 99.07056, 99.73713, 99.54643, 
    99.74157, 99.61737, 96.52483, 96.67683, 96.59469, 96.74921, 96.64034, 
    97.12502, 97.27062, 97.95357, 97.67289, 98.11976, 97.71822, 97.78931, 
    98.13443, 97.73988, 98.60384, 98.01768, 99.10804, 98.52103, 99.1449, 
    99.03141, 99.21933, 99.38783, 99.60001, 99.99225, 99.90133, 100.2298, 
    96.90368, 97.10133, 97.08389, 97.29095, 97.44425, 97.77699, 98.31208, 
    98.11065, 98.48059, 98.55497, 97.99299, 98.33784, 97.23373, 97.41165, 
    97.30566, 96.91928, 98.1571, 97.52071, 98.6977, 98.35153, 99.36379, 
    98.85966, 99.85131, 100.2771, 100.6785, 101.1491, 97.20927, 97.07486, 
    97.31557, 97.64927, 97.95939, 98.37263, 98.41495, 98.49251, 98.69353, 
    98.86275, 98.51707, 98.9052, 97.45301, 98.21243, 97.0241, 97.38108, 
    97.62957, 97.52048, 98.08763, 98.2216, 98.7671, 98.48486, 100.1719, 
    99.42349, 101.508, 100.923, 97.02793, 97.20879, 97.83987, 97.53929, 
    98.40023, 98.61285, 98.78586, 99.00733, 99.03123, 99.1626, 98.94738, 
    99.15408, 98.37351, 98.72189, 97.76757, 97.99936, 97.89268, 97.77576, 
    98.13687, 98.52252, 98.53071, 98.65457, 99.0042, 98.40373, 100.2689, 
    99.11472, 97.40624, 97.75568, 97.80558, 97.6701, 98.59152, 98.25708, 
    99.15939, 98.91504, 99.31557, 99.11642, 99.08715, 98.83175, 98.67295, 
    98.27242, 97.9472, 97.68974, 97.74956, 98.0325, 98.54613, 99.03342, 
    98.92657, 99.2851, 98.33766, 98.73433, 98.58092, 98.98119, 98.10531, 
    98.85107, 97.91525, 97.99707, 98.25045, 98.76131, 98.87444, 98.99545, 
    98.92076, 98.55917, 98.49998, 98.24427, 98.17377, 97.97925, 97.81841, 
    97.96537, 98.11986, 98.5593, 98.95633, 99.39024, 99.49657, 100.0054, 
    99.59115, 100.2753, 99.6936, 100.7018, 98.89429, 99.67641, 98.26196, 
    98.41376, 98.68874, 99.32098, 98.97931, 99.37894, 98.49766, 98.0423, 
    97.92461, 97.70538, 97.92963, 97.91138, 98.12622, 98.05714, 98.57391, 
    98.29613, 99.08643, 99.37576, 100.1954, 100.6998, 101.2146, 101.4424, 
    101.5118, 101.5408,
  94.75323, 95.22436, 95.13264, 95.51013, 95.30208, 95.54713, 94.84859, 
    95.24313, 94.99113, 94.79553, 96.22945, 95.52661, 96.9625, 96.51182, 
    97.64631, 96.89234, 97.79875, 97.6244, 98.14948, 97.99887, 98.67258, 
    98.21904, 99.02277, 98.5641, 98.6358, 98.20412, 95.66769, 96.1418, 
    95.63968, 95.70718, 95.67686, 95.30647, 95.11588, 94.71722, 94.78951, 
    95.08231, 95.73753, 95.51806, 96.0716, 96.05908, 96.67772, 96.39848, 
    97.4419, 97.14462, 98.00515, 97.78831, 97.99498, 97.93227, 97.9958, 
    97.67789, 97.81403, 97.53453, 96.45076, 96.76852, 95.82278, 95.25248, 
    94.86589, 94.59222, 94.63088, 94.70463, 95.08403, 95.44034, 95.70503, 
    95.88236, 96.05728, 96.58822, 96.86975, 97.50214, 97.38774, 97.58153, 
    97.76675, 98.07834, 98.027, 98.16444, 97.57635, 97.96699, 97.32263, 
    97.49862, 96.10521, 95.57722, 95.35209, 95.15028, 94.66062, 94.99862, 
    94.8653, 95.1826, 95.3846, 95.28465, 95.88721, 95.65408, 96.88645, 
    96.35442, 97.74513, 97.4112, 97.82526, 97.61383, 97.97632, 97.65004, 
    98.2156, 98.33905, 98.25468, 98.5789, 97.63198, 97.99501, 95.28186, 
    95.29816, 95.37408, 95.04064, 95.02025, 94.71526, 94.98658, 95.10229, 
    95.39629, 95.56541, 95.72613, 96.08011, 96.47647, 97.03233, 97.43283, 
    97.70189, 97.53683, 97.68255, 97.51968, 97.44337, 98.29281, 97.81532, 
    98.53223, 98.49246, 98.16772, 98.49694, 95.3096, 95.21584, 94.89082, 
    95.14512, 94.68208, 94.94113, 95.09031, 95.65903, 95.78208, 95.89639, 
    96.1223, 96.41277, 96.92365, 97.36948, 97.77752, 97.74758, 97.75813, 
    97.84944, 97.62337, 97.88659, 97.93084, 97.81522, 98.48714, 98.29488, 
    98.49162, 98.3664, 95.2463, 95.40408, 95.31882, 95.47695, 95.36625, 
    95.85536, 96.00198, 96.6898, 96.40706, 96.8572, 96.4527, 96.52431, 
    96.87205, 96.47451, 97.34493, 96.75441, 97.853, 97.26153, 97.89014, 
    97.77575, 97.96515, 98.13501, 98.34889, 98.74439, 98.65271, 98.98396, 
    95.63245, 95.83149, 95.8139, 96.02239, 96.17679, 96.51189, 97.05093, 
    96.84798, 97.22069, 97.29564, 96.72945, 97.0769, 95.96479, 96.144, 
    96.03722, 95.64819, 96.89482, 96.25382, 97.43948, 97.09067, 98.11079, 
    97.60271, 98.60227, 99.03165, 99.43649, 99.91122, 95.94016, 95.8048, 
    96.04719, 96.3833, 96.69563, 97.11194, 97.15456, 97.23271, 97.43525, 
    97.60578, 97.25749, 97.64855, 96.18571, 96.95055, 95.75372, 96.11322, 
    96.36344, 96.25356, 96.82479, 96.95975, 97.50942, 97.225, 98.92564, 
    98.17101, 100.2734, 99.68318, 95.75755, 95.93966, 96.57526, 96.2725, 
    97.13973, 97.35397, 97.52829, 97.7515, 97.77557, 97.90799, 97.69107, 
    97.89939, 97.11282, 97.46383, 96.5024, 96.73589, 96.62841, 96.51064, 
    96.8744, 97.26299, 97.27119, 97.39603, 97.74851, 97.14325, 99.02348, 
    97.85987, 96.1385, 96.49048, 96.5407, 96.40423, 97.33248, 96.99551, 
    97.90475, 97.65848, 98.06216, 97.86144, 97.83194, 97.57454, 97.41453, 
    97.01097, 96.68336, 96.424, 96.48426, 96.76929, 97.28677, 97.7778, 
    97.67012, 98.03144, 97.07669, 97.47639, 97.32182, 97.72515, 96.84262, 
    97.59415, 96.65114, 96.73357, 96.98883, 97.50361, 97.61757, 97.73952, 
    97.66424, 97.2999, 97.24025, 96.9826, 96.91159, 96.71561, 96.5536, 
    96.70164, 96.85729, 97.30001, 97.70011, 98.13744, 98.24461, 98.75772, 
    98.34005, 99.03001, 98.44345, 99.46004, 97.63766, 98.42602, 97.00043, 
    97.15337, 97.43048, 98.06769, 97.72325, 98.12609, 97.2379, 96.77918, 
    96.66058, 96.43977, 96.66564, 96.64725, 96.86367, 96.79408, 97.31473, 
    97.03484, 97.83123, 98.12288, 98.94925, 99.45798, 99.97729, 100.2071, 
    100.2771, 100.3064,
  129.942, 130.6547, 130.5159, 131.0834, 130.7723, 131.1393, 130.0862, 
    130.6831, 130.3018, 130.006, 132.1703, 131.1083, 133.2786, 132.5972, 
    134.3131, 133.1725, 134.5439, 134.28, 135.0748, 134.8468, 135.8669, 
    135.1801, 136.3975, 135.7027, 135.8112, 135.1575, 131.3215, 132.0378, 
    131.2791, 131.3811, 131.3353, 130.779, 130.4906, 129.8876, 129.9969, 
    130.4398, 131.427, 131.0954, 131.9318, 131.9128, 132.848, 132.4258, 
    134.0038, 133.5541, 134.8563, 134.5281, 134.8409, 134.746, 134.8421, 
    134.3609, 134.567, 134.144, 132.5049, 132.9853, 131.5558, 130.6973, 
    130.1124, 129.6985, 129.757, 129.8685, 130.4424, 130.978, 131.3779, 
    131.6458, 131.9101, 132.7126, 133.1384, 134.095, 133.9219, 134.2151, 
    134.4954, 134.9671, 134.8894, 135.0974, 134.2073, 134.7985, 133.8234, 
    134.0897, 131.9825, 131.1848, 130.8471, 130.5426, 129.8019, 130.3132, 
    130.1115, 130.5915, 130.8947, 130.7459, 131.6531, 131.3009, 133.1636, 
    132.3592, 134.4627, 133.9574, 134.584, 134.264, 134.8126, 134.3188, 
    135.1749, 135.3618, 135.2341, 135.7251, 134.2915, 134.8409, 130.7417, 
    130.7664, 130.8793, 130.3768, 130.3459, 129.8846, 130.295, 130.47, 
    130.9118, 131.1669, 131.4097, 131.9446, 132.5437, 133.3842, 133.9901, 
    134.3973, 134.1475, 134.368, 134.1215, 134.0061, 135.2918, 134.5689, 
    135.6544, 135.5942, 135.1024, 135.6009, 130.7837, 130.6418, 130.1501, 
    130.5348, 129.8344, 130.2262, 130.4519, 131.3084, 131.4943, 131.667, 
    132.0084, 132.4474, 133.2199, 133.8943, 134.5117, 134.4664, 134.4824, 
    134.6206, 134.2785, 134.6768, 134.7438, 134.5688, 135.5861, 135.295, 
    135.5929, 135.4032, 130.6879, 130.9233, 130.7977, 131.0333, 130.8678, 
    131.605, 131.8265, 132.8663, 132.4388, 133.1194, 132.5078, 132.6161, 
    133.1418, 132.5408, 133.8571, 132.9639, 134.626, 133.7309, 134.6822, 
    134.5091, 134.7957, 135.0529, 135.3767, 135.9757, 135.8369, 136.3387, 
    131.2682, 131.5689, 131.5423, 131.8574, 132.0907, 132.5973, 133.4124, 
    133.1055, 133.6692, 133.7826, 132.9262, 133.4517, 131.7704, 132.0412, 
    131.8798, 131.292, 133.1763, 132.2072, 134.0002, 133.4725, 135.0162, 
    134.2472, 135.7605, 136.4109, 137.0245, 137.7442, 131.7331, 131.5286, 
    131.8949, 132.4029, 132.8751, 133.5047, 133.5691, 133.6874, 133.9938, 
    134.2518, 133.7248, 134.3166, 132.1042, 133.2606, 131.4514, 131.9946, 
    132.3728, 132.2068, 133.0704, 133.2745, 134.106, 133.6757, 136.2503, 
    135.1074, 138.2935, 137.3984, 131.4572, 131.7324, 132.6931, 132.2354, 
    133.5467, 133.8708, 134.1346, 134.4724, 134.5088, 134.7092, 134.3809, 
    134.6962, 133.506, 134.037, 132.5829, 132.936, 132.7734, 132.5954, 
    133.1454, 133.7331, 133.7456, 133.9344, 134.4678, 133.552, 136.3985, 
    134.6363, 132.0329, 132.5649, 132.6408, 132.4345, 133.8383, 133.3286, 
    134.7043, 134.3316, 134.9426, 134.6388, 134.5941, 134.2045, 133.9624, 
    133.3519, 132.8565, 132.4644, 132.5555, 132.9865, 133.7691, 134.5122, 
    134.3492, 134.8961, 133.4514, 134.056, 133.8222, 134.4325, 133.0974, 
    134.2342, 132.8078, 132.9324, 133.3185, 134.0972, 134.2697, 134.4542, 
    134.3403, 133.789, 133.6988, 133.3091, 133.2016, 132.9053, 132.6603, 
    132.8842, 133.1195, 133.7892, 134.3946, 135.0566, 135.2188, 135.9959, 
    135.3633, 136.4084, 135.5199, 137.0601, 134.3, 135.4935, 133.336, 
    133.5673, 133.9865, 134.9509, 134.4296, 135.0394, 133.6952, 133.0014, 
    132.8221, 132.4883, 132.8297, 132.8019, 133.1292, 133.024, 133.8114, 
    133.3881, 134.593, 135.0345, 136.2861, 137.057, 137.8444, 138.193, 
    138.2992, 138.3436,
  195.776, 196.8889, 196.6722, 197.5725, 197.0726, 197.6627, 196.0012, 
    196.9333, 196.3379, 195.8759, 199.3283, 197.6127, 201.121, 200.0186, 
    202.7959, 200.9493, 203.1697, 202.7423, 204.0302, 203.6606, 205.2841, 
    204.2009, 206.116, 205.0266, 205.1968, 204.1643, 197.9569, 199.1142, 
    197.8885, 198.0532, 197.9793, 197.083, 196.6326, 195.6911, 195.8617, 
    196.5533, 198.1273, 197.5919, 198.943, 198.9124, 200.4243, 199.7416, 
    202.295, 201.5669, 203.676, 203.1441, 203.651, 203.4972, 203.6531, 
    202.8734, 203.2072, 202.522, 199.8694, 200.6464, 198.3354, 196.9553, 
    196.0421, 195.396, 195.4872, 195.6613, 196.5573, 197.4023, 198.048, 
    198.4809, 198.908, 200.2053, 200.894, 202.4426, 202.1624, 202.6372, 
    203.0913, 203.8556, 203.7296, 204.0669, 202.6245, 203.5824, 202.0029, 
    202.434, 199.0248, 197.7362, 197.1908, 196.7139, 195.5574, 196.3555, 
    196.0406, 196.7903, 197.2677, 197.0314, 198.4927, 197.9237, 200.9349, 
    199.6339, 203.0383, 202.2198, 203.2348, 202.7164, 203.6053, 202.8052, 
    204.1925, 204.4924, 204.2884, 205.0617, 202.7609, 203.6511, 197.0249, 
    197.0634, 197.2429, 196.4548, 196.4066, 195.6864, 196.3271, 196.6005, 
    197.2954, 197.7074, 198.0995, 198.9637, 199.9322, 201.2919, 202.2728, 
    202.9323, 202.5277, 202.8849, 202.4856, 202.2987, 204.382, 203.2103, 
    204.9509, 204.8565, 204.0749, 204.8672, 197.0904, 196.8688, 196.1009, 
    196.7017, 195.6081, 196.2198, 196.5721, 197.9357, 198.2361, 198.5151, 
    199.0668, 199.7765, 201.026, 202.1176, 203.1177, 203.0443, 203.0701, 
    203.2941, 202.7398, 203.3852, 203.4937, 203.2101, 204.8439, 204.3871, 
    204.8545, 204.5574, 196.9408, 197.3139, 197.1122, 197.4916, 197.2243, 
    198.4149, 198.7728, 200.4538, 199.7625, 200.8633, 199.8741, 200.0492, 
    200.8996, 199.9274, 202.0574, 200.6118, 203.3028, 201.8531, 203.3939, 
    203.1134, 203.5779, 203.9947, 204.5158, 205.4546, 205.2369, 206.0238, 
    197.8709, 198.3566, 198.3137, 198.8228, 199.1999, 200.0188, 201.3375, 
    200.8409, 201.7532, 201.9368, 200.5509, 201.4011, 198.6821, 199.1197, 
    198.859, 197.9093, 200.9554, 199.388, 202.2891, 201.4348, 203.9352, 
    202.6891, 205.1172, 206.1371, 207.0998, 208.2298, 198.6219, 198.2915, 
    198.8833, 199.7044, 200.4681, 201.4869, 201.5912, 201.7826, 202.2788, 
    202.6967, 201.8433, 202.8015, 199.2215, 201.0918, 198.1668, 199.0445, 
    199.6559, 199.3874, 200.7841, 201.1144, 202.4604, 201.7637, 205.8851, 
    204.0829, 209.0928, 207.6868, 198.1762, 198.6208, 200.1737, 199.4337, 
    201.5549, 202.0796, 202.5067, 203.0539, 203.1129, 203.4377, 202.9057, 
    203.4166, 201.489, 202.3488, 199.9956, 200.5666, 200.3038, 200.0158, 
    200.9055, 201.8567, 201.8769, 202.1826, 203.0463, 201.5636, 206.1175, 
    203.3194, 199.1063, 199.9664, 200.0892, 199.7557, 202.027, 201.2019, 
    203.4297, 202.8258, 203.8159, 203.3235, 203.2511, 202.6201, 202.228, 
    201.2397, 200.4381, 199.804, 199.9513, 200.6483, 201.9149, 203.1184, 
    202.8543, 203.7405, 201.4006, 202.3795, 202.0008, 202.9893, 200.8277, 
    202.6679, 200.3593, 200.561, 201.1855, 202.4462, 202.7256, 203.0245, 
    202.84, 201.9471, 201.8011, 201.1703, 200.9965, 200.517, 200.1208, 
    200.4828, 200.8636, 201.9474, 202.9279, 204.0006, 204.2637, 205.4862, 
    204.4948, 206.133, 204.74, 207.1557, 202.7747, 204.6987, 201.2139, 
    201.5883, 202.267, 203.8294, 202.9846, 203.9727, 201.7953, 200.6725, 
    200.3824, 199.8425, 200.3948, 200.3498, 200.8792, 200.709, 201.9835, 
    201.2982, 203.2494, 203.9648, 205.9413, 207.1509, 208.3872, 208.9349, 
    209.1018, 209.1716,
  319.7119, 321.5092, 321.159, 322.6142, 321.8061, 322.7602, 320.0754, 
    321.5808, 320.619, 319.8731, 325.4563, 322.6793, 328.3638, 326.5753, 
    331.0854, 328.085, 331.6935, 330.9982, 333.0882, 332.4926, 335.1112, 
    333.357, 336.4688, 334.6913, 334.9688, 333.2993, 323.2361, 325.1094, 
    323.1255, 323.3919, 323.2723, 321.8229, 321.0949, 319.5747, 319.8502, 
    320.9669, 323.5117, 322.6456, 324.8322, 324.7827, 327.2332, 326.1262, 
    330.271, 329.0879, 332.5176, 331.652, 332.477, 332.2266, 332.4803, 
    331.2115, 331.7545, 330.6401, 326.3333, 327.5936, 323.8485, 321.6164, 
    320.1413, 319.0986, 319.2458, 319.5267, 320.9734, 322.3391, 323.3835, 
    324.084, 324.7755, 326.8779, 327.9954, 330.5109, 330.0554, 330.8272, 
    331.5659, 332.81, 332.6049, 333.146, 330.8067, 332.3651, 329.7962, 
    330.497, 324.9646, 322.879, 321.997, 321.2263, 319.359, 320.6475, 
    320.139, 321.3498, 322.1215, 321.7396, 324.1032, 323.1824, 328.0617, 
    325.9515, 331.4797, 330.1488, 331.7994, 330.9561, 332.4024, 331.1005, 
    333.3436, 333.8207, 333.4946, 334.7487, 331.0285, 332.4771, 321.7289, 
    321.7912, 322.0813, 320.8078, 320.73, 319.5672, 320.6016, 321.0432, 
    322.1662, 322.8324, 323.4668, 324.8658, 326.4351, 328.6413, 330.2349, 
    331.3073, 330.6493, 331.2301, 330.5809, 330.277, 333.6419, 331.7596, 
    334.568, 334.4142, 333.1586, 334.4315, 321.8349, 321.4767, 320.2364, 
    321.2067, 319.4408, 320.4282, 320.9973, 323.2018, 323.6878, 324.1394, 
    325.0327, 326.1828, 328.2096, 329.9826, 331.6089, 331.4895, 331.5316, 
    331.8959, 330.9942, 332.0442, 332.2208, 331.7593, 334.3936, 333.6501, 
    334.4109, 333.9265, 321.5931, 322.1961, 321.8701, 322.4834, 322.0513, 
    323.9771, 324.5566, 327.2811, 326.1602, 327.9456, 326.341, 326.6248, 
    328.0043, 326.4275, 329.8847, 327.5374, 331.9101, 329.5527, 332.0583, 
    331.6019, 332.3579, 333.0323, 333.8589, 335.3895, 335.0344, 336.3183, 
    323.097, 323.8829, 323.8135, 324.6376, 325.2483, 326.5757, 328.7154, 
    327.9091, 329.3905, 329.6887, 327.4386, 328.8186, 324.4097, 325.1184, 
    324.6962, 323.159, 328.095, 325.5531, 330.2614, 328.8734, 332.9388, 
    330.9117, 334.8391, 336.5031, 338.076, 339.9241, 324.3124, 323.7776, 
    324.7357, 326.0659, 327.3044, 328.9579, 329.1274, 329.4383, 330.2446, 
    330.9241, 329.5368, 331.0946, 325.2833, 328.3164, 323.5757, 324.9966, 
    325.9873, 325.5522, 327.8171, 328.3531, 330.5399, 329.4077, 336.0918, 
    333.1712, 341.3375, 339.0357, 323.5909, 324.3105, 326.8268, 325.6272, 
    329.0685, 329.9209, 330.6152, 331.5051, 331.6012, 332.1296, 331.2641, 
    332.0953, 328.9614, 330.3584, 326.5381, 327.4641, 327.0377, 326.5707, 
    328.0141, 329.5586, 329.5915, 330.0883, 331.4925, 329.0825, 336.4711, 
    331.937, 325.0968, 326.4906, 326.6898, 326.149, 329.8354, 328.4951, 
    332.1167, 331.1341, 332.7454, 331.9438, 331.826, 330.7995, 330.162, 
    328.5565, 327.2556, 326.2274, 326.4662, 327.5966, 329.6533, 331.61, 
    331.1805, 332.6227, 328.8178, 330.4084, 329.7928, 331.4, 327.8878, 
    330.8772, 327.1279, 327.455, 328.4686, 330.5167, 330.971, 331.4573, 
    331.1571, 329.7056, 329.4683, 328.4439, 328.1617, 327.3837, 326.7411, 
    327.3282, 327.946, 329.7061, 331.3001, 333.0417, 333.4557, 335.4409, 
    333.8244, 336.4964, 334.2238, 338.1671, 331.0508, 334.1567, 328.5147, 
    329.1227, 330.2254, 332.7672, 331.3924, 332.9977, 329.459, 327.6358, 
    327.1654, 326.2898, 327.1854, 327.1125, 327.9714, 327.6952, 329.7647, 
    328.6515, 331.8232, 332.9854, 336.1836, 338.1594, 340.182, 341.0789, 
    341.3523, 341.4667,
  524.6366, 527.9116, 527.2736, 529.9268, 528.4529, 530.1931, 525.3011, 
    528.0422, 526.2903, 524.9333, 535.1226, 530.0454, 540.4584, 537.174, 
    545.4717, 539.9459, 546.5943, 545.3109, 549.1841, 548.071, 553.0635, 
    549.6988, 555.6735, 552.2574, 552.7902, 549.5883, 531.0621, 534.4874, 
    530.8601, 531.3466, 531.1282, 528.4834, 527.1569, 524.3786, 524.8915, 
    526.9237, 531.5656, 529.9841, 533.9803, 533.8896, 538.3814, 536.3504, 
    543.9698, 541.7906, 548.1174, 546.5177, 548.0422, 547.5793, 548.0482, 
    545.7044, 546.7071, 544.6502, 536.7302, 539.043, 532.181, 528.107, 
    525.4211, 523.4829, 523.7598, 524.2881, 526.9356, 529.4248, 531.3315, 
    532.6116, 533.8766, 537.7291, 539.7812, 544.4119, 543.5723, 544.9954, 
    546.3588, 548.658, 548.2787, 549.2946, 544.9576, 547.8353, 543.0948, 
    544.3863, 534.2224, 530.4101, 528.8008, 527.3962, 523.9728, 526.3422, 
    525.4169, 527.6212, 529.0279, 528.3315, 532.6467, 530.964, 539.9031, 
    536.0302, 546.1996, 543.7444, 546.79, 545.2333, 547.9042, 545.4996, 
    549.6733, 550.5875, 549.9626, 552.3676, 545.3668, 548.0423, 528.3121, 
    528.4256, 528.9547, 526.6341, 526.4925, 524.3644, 526.2587, 527.0626, 
    529.1095, 530.325, 531.4835, 534.0417, 536.9168, 540.9689, 543.9032, 
    545.8812, 544.6672, 545.7389, 544.5411, 543.9807, 550.2448, 546.7166, 
    552.0209, 551.7256, 549.3189, 551.7589, 528.5053, 527.8525, 525.5941, 
    527.3605, 524.1266, 525.9431, 526.9792, 530.9994, 531.8874, 532.7128, 
    534.3473, 536.4542, 540.1749, 543.4381, 546.4382, 546.2177, 546.2953, 
    546.9683, 545.3034, 547.2422, 547.5685, 546.7159, 551.6862, 550.2604, 
    551.7194, 550.7905, 528.0646, 529.164, 528.5696, 529.6881, 528.8999, 
    532.4161, 533.4759, 538.4691, 536.4127, 539.6898, 536.7443, 537.2648, 
    539.7976, 536.9029, 543.2578, 538.9398, 546.9944, 542.6461, 547.2684, 
    546.4252, 547.822, 549.077, 550.6606, 553.5982, 552.9162, 555.384, 
    530.8082, 532.2439, 532.1171, 533.624, 534.742, 537.1746, 541.1051, 
    539.6229, 542.3477, 542.8968, 538.7585, 541.2949, 533.2072, 534.504, 
    533.7313, 530.9214, 539.9643, 535.3001, 543.9519, 541.3958, 548.8979, 
    545.1511, 552.5412, 555.7395, 558.7698, 562.2432, 533.0292, 532.0514, 
    533.8035, 536.2398, 538.5119, 541.5513, 541.8633, 542.4356, 543.9211, 
    545.1741, 542.6169, 545.4887, 534.8058, 540.3714, 531.6825, 534.2811, 
    536.0958, 535.2985, 539.4537, 540.4389, 544.4655, 542.3792, 554.9482, 
    549.3428, 564.8879, 560.5837, 531.7103, 533.0258, 537.6353, 535.436, 
    541.7548, 543.3245, 544.6044, 546.2464, 546.4239, 547.4, 545.8016, 
    547.3367, 541.5578, 544.1308, 537.1057, 538.8053, 538.0225, 537.1656, 
    539.8157, 542.6571, 542.7177, 543.6329, 546.223, 541.7806, 555.6777, 
    547.0439, 534.4647, 537.0185, 537.384, 536.3922, 543.1669, 540.7001, 
    547.3762, 545.5617, 548.5385, 547.0568, 546.8392, 544.9443, 543.7689, 
    540.8129, 538.4224, 536.5359, 536.9738, 539.0486, 542.8314, 546.4401, 
    545.6472, 548.3116, 541.2936, 544.2229, 543.0885, 546.0524, 539.5836, 
    545.0873, 538.188, 538.7885, 540.6512, 544.4225, 545.2607, 546.1582, 
    545.6041, 542.9279, 542.4908, 540.6058, 540.0869, 538.6577, 537.4781, 
    538.5558, 539.6906, 542.9288, 545.868, 549.0949, 549.8881, 553.6968, 
    550.5944, 555.7263, 551.3602, 558.9454, 545.4078, 551.2317, 540.736, 
    541.8547, 543.8856, 548.5788, 546.0385, 549.0107, 542.4736, 539.1206, 
    538.2568, 536.6505, 538.2936, 538.1597, 539.7373, 539.2297, 543.0367, 
    540.9876, 546.8339, 548.987, 555.1248, 558.9306, 562.7255, 564.4036, 
    564.9157, 565.13,
  947.2838, 954.1565, 952.8134, 958.4072, 955.2968, 958.9701, 948.6699, 
    954.4314, 950.7462, 947.8986, 969.2882, 958.658, 980.3278, 973.521, 
    990.7889, 979.2632, 993.1437, 990.4521, 998.593, 996.2479, 1006.801, 
    999.6788, 1012.354, 1005.091, 1006.221, 999.4456, 960.8081, 967.9803, 
    960.3806, 961.4105, 960.9479, 955.3611, 952.5678, 946.7616, 947.811, 
    952.0774, 961.8741, 958.5283, 966.9372, 966.7508, 976.019, 971.82, 
    987.6458, 983.0991, 996.3455, 992.9828, 996.1872, 995.2134, 996.1999, 
    991.2768, 993.3806, 989.0688, 972.6041, 977.39, 963.1785, 954.5679, 
    948.9214, 944.9504, 945.51, 946.5786, 952.1025, 957.3471, 961.3783, 
    964.0917, 966.7241, 974.6688, 978.9212, 988.5703, 986.8152, 989.7914, 
    992.6495, 997.4839, 996.6851, 998.826, 989.7122, 995.752, 985.8182, 
    988.5168, 967.435, 959.4288, 956.0305, 953.0714, 945.9407, 950.8552, 
    948.9126, 953.545, 956.5095, 955.0412, 964.1661, 960.6005, 979.1744, 
    971.1592, 992.3153, 987.1749, 993.5548, 990.2895, 995.897, 990.8477, 
    999.6249, 1001.556, 1000.236, 1005.325, 990.5692, 996.1874, 955.0002, 
    955.2394, 956.3549, 951.4686, 951.171, 946.733, 950.6799, 952.3696, 
    956.6816, 959.2488, 961.7004, 967.0636, 972.9896, 981.389, 987.5067, 
    991.6476, 989.1044, 991.3491, 988.8405, 987.6687, 1000.832, 993.4003, 
    1004.59, 1003.964, 998.8771, 1004.035, 955.4074, 954.032, 949.2844, 
    952.9963, 946.2518, 950.017, 952.194, 960.6753, 962.556, 964.3065, 
    967.6921, 972.0342, 979.7388, 986.535, 992.8161, 992.3533, 992.5162, 
    993.9291, 990.4365, 994.5047, 995.1908, 993.3992, 1003.88, 1000.865, 
    1003.951, 1001.985, 954.4786, 956.7967, 955.5429, 957.9031, 956.2395, 
    963.677, 965.9006, 976.2007, 971.9485, 978.7315, 972.6333, 973.7089, 
    978.9553, 972.9609, 986.1584, 977.1759, 993.9841, 984.882, 994.5598, 
    992.7888, 995.724, 998.3671, 1001.711, 1007.937, 1006.488, 1011.737, 
    960.2707, 963.3118, 963.0428, 966.205, 968.5044, 973.5224, 981.6723, 
    978.5927, 984.2598, 985.405, 976.8003, 982.0673, 965.3487, 968.0146, 
    966.4254, 960.5102, 979.3014, 969.654, 987.6085, 982.2772, 997.9894, 
    990.1175, 1005.693, 1012.495, 1018.976, 1026.654, 964.9781, 962.9037, 
    966.5739, 971.5918, 976.2894, 982.6009, 983.2507, 984.4432, 987.544, 
    990.1655, 984.8212, 990.8247, 968.6357, 980.147, 962.1218, 967.5558, 
    971.2944, 969.6507, 978.2417, 980.2872, 988.6823, 984.3256, 1010.809, 
    998.9277, 1032.464, 1022.954, 962.1808, 964.9708, 974.4749, 969.9339, 
    983.0247, 986.2977, 988.973, 992.4136, 992.7859, 994.8365, 991.4806, 
    994.7034, 982.6144, 987.9824, 973.3799, 976.8972, 975.2761, 973.5038, 
    978.9928, 984.9051, 985.0313, 986.9418, 992.3644, 983.0784, 1012.363, 
    994.088, 967.9336, 973.1998, 973.9554, 971.9064, 985.9686, 980.83, 
    994.7863, 990.9777, 997.2323, 994.1151, 993.6581, 989.6845, 987.2259, 
    981.0647, 976.1041, 972.2029, 973.1074, 977.4017, 985.2687, 992.8201, 
    991.1567, 996.7543, 982.0645, 988.1749, 985.8051, 992.0067, 978.5112, 
    989.9838, 975.6187, 976.8624, 980.7285, 988.5925, 990.3471, 992.2285, 
    991.0666, 985.4698, 984.5582, 980.634, 979.5561, 976.5913, 974.1497, 
    976.3802, 978.7332, 985.4718, 991.6197, 998.4048, 1000.078, 1008.146, 
    1001.57, 1012.467, 1003.19, 1019.352, 990.6552, 1002.918, 980.9048, 
    983.2325, 987.4698, 997.3171, 991.9773, 998.2272, 984.5224, 977.5508, 
    975.761, 972.4395, 975.8372, 975.56, 978.8303, 977.7771, 985.697, 
    981.428, 993.6468, 998.1774, 1011.185, 1019.321, 1027.732, 1031.413, 
    1032.524, 1032.99,
  1829.892, 1849.354, 1845.526, 1861.551, 1852.614, 1863.175, 1833.792, 
    1850.139, 1839.658, 1831.62, 1893.773, 1862.274, 1928.095, 1906.815, 
    1960.692, 1924.742, 1968.122, 1959.633, 1985.508, 1977.993, 2012.213, 
    1989.004, 2030.649, 2006.597, 2010.305, 1988.253, 1868.495, 1889.772, 
    1867.256, 1870.244, 1868.901, 1852.798, 1844.827, 1828.426, 1831.374, 
    1843.433, 1871.592, 1861.9, 1886.59, 1886.023, 1914.58, 1901.557, 
    1950.849, 1936.76, 1978.305, 1967.613, 1977.799, 1974.694, 1977.84, 
    1962.227, 1968.872, 1955.294, 1903.978, 1918.864, 1875.391, 1850.529, 
    1834.501, 1823.355, 1824.92, 1827.913, 1843.505, 1858.498, 1870.151, 
    1878.059, 1885.941, 1910.377, 1923.666, 1953.735, 1948.262, 1957.558, 
    1966.559, 1981.948, 1979.39, 1986.257, 1957.31, 1976.41, 1945.165, 
    1953.568, 1888.107, 1864.501, 1854.716, 1846.261, 1826.125, 1839.966, 
    1834.476, 1847.61, 1856.09, 1851.883, 1878.276, 1867.893, 1924.462, 
    1899.52, 1965.503, 1949.381, 1969.424, 1959.122, 1976.873, 1960.876, 
    1988.83, 1995.075, 1990.802, 2007.362, 1960.001, 1977.8, 1851.765, 
    1852.45, 1855.647, 1841.705, 1840.861, 1828.346, 1839.47, 1844.264, 
    1856.585, 1863.981, 1871.086, 1886.975, 1905.17, 1931.448, 1950.415, 
    1963.396, 1955.406, 1962.455, 1954.58, 1950.92, 1992.729, 1968.935, 
    2004.955, 2002.911, 1986.422, 2003.141, 1852.931, 1848.999, 1835.525, 
    1846.047, 1826.997, 1837.595, 1843.765, 1868.11, 1873.576, 1878.687, 
    1888.892, 1902.217, 1926.239, 1947.39, 1967.086, 1965.623, 1966.137, 
    1970.612, 1959.584, 1972.439, 1974.622, 1968.931, 2002.638, 1992.836, 
    2002.868, 1996.467, 1850.274, 1856.915, 1853.319, 1860.098, 1855.316, 
    1876.847, 1883.437, 1915.147, 1901.953, 1923.07, 1904.068, 1907.397, 
    1923.773, 1905.081, 1946.221, 1918.194, 1970.786, 1942.264, 1972.615, 
    1966.999, 1976.321, 1984.782, 1995.576, 2015.958, 2011.184, 2028.585, 
    1866.937, 1875.78, 1874.995, 1884.362, 1891.373, 1906.819, 1932.345, 
    1922.634, 1940.34, 1943.883, 1917.019, 1933.587, 1881.762, 1889.876, 
    1885.032, 1867.631, 1924.862, 1894.894, 1950.732, 1934.232, 1983.569, 
    1958.582, 2008.57, 2031.12, 2053.035, 2079.241, 1880.653, 1874.59, 
    1885.484, 1900.853, 1915.424, 1935.227, 1937.227, 1940.906, 1950.531, 
    1958.733, 1942.076, 1960.804, 1891.775, 1927.525, 1872.312, 1888.476, 
    1899.937, 1894.884, 1921.533, 1927.967, 1954.085, 1940.543, 2025.486, 
    1986.585, 2099.51, 2066.706, 1872.484, 1880.632, 1909.774, 1895.753, 
    1936.531, 1946.653, 1954.994, 1965.813, 1966.99, 1973.494, 1962.869, 
    1973.071, 1935.268, 1951.899, 1906.378, 1917.322, 1912.265, 1906.762, 
    1923.891, 1942.335, 1942.726, 1948.656, 1965.658, 1936.696, 2030.678, 
    1971.116, 1889.629, 1905.82, 1908.162, 1901.823, 1945.631, 1929.681, 
    1973.335, 1961.286, 1981.141, 1971.202, 1969.752, 1957.223, 1949.54, 
    1930.422, 1914.845, 1902.738, 1905.534, 1918.9, 1943.461, 1967.098, 
    1961.849, 1979.612, 1933.578, 1952.5, 1945.124, 1964.528, 1922.379, 
    1958.162, 1913.332, 1917.214, 1929.36, 1953.804, 1959.303, 1965.228, 
    1961.565, 1944.084, 1941.262, 1929.062, 1925.663, 1916.366, 1908.765, 
    1915.707, 1923.075, 1944.09, 1963.308, 1984.903, 1990.294, 2016.65, 
    1995.122, 2031.026, 2000.387, 2054.322, 1960.271, 1999.501, 1929.917, 
    1937.171, 1950.3, 1981.413, 1964.435, 1984.333, 1941.151, 1919.367, 
    1913.776, 1903.469, 1914.013, 1913.15, 1923.38, 1920.076, 1944.789, 
    1931.571, 1969.716, 1984.172, 2026.741, 2054.214, 2082.901, 2095.762, 
    2099.725, 2101.389,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.536768, 4.555262, 4.551662, 4.566609, 4.558312, 4.568107, 4.540512, 
    4.555998, 4.546107, 4.53843, 4.595716, 4.567276, 4.625376, 4.607146, 
    4.65303, 4.622537, 4.659195, 4.652147, 4.673377, 4.667288, 4.694517, 
    4.676189, 4.70867, 4.690135, 4.693032, 4.675585, 4.572988, 4.592169, 
    4.571854, 4.574585, 4.573359, 4.558485, 4.551003, 4.535356, 4.538193, 
    4.549686, 4.575813, 4.566931, 4.589335, 4.588828, 4.613858, 4.602561, 
    4.644767, 4.632744, 4.667542, 4.658775, 4.66713, 4.664596, 4.667163, 
    4.65431, 4.659814, 4.648513, 4.604676, 4.617531, 4.579264, 4.556363, 
    4.541191, 4.530447, 4.531965, 4.53486, 4.549754, 4.563786, 4.5745, 
    4.581676, 4.588755, 4.610233, 4.621624, 4.647202, 4.642577, 4.650412, 
    4.657903, 4.6705, 4.668425, 4.673981, 4.650204, 4.665998, 4.639945, 
    4.647061, 4.590688, 4.569326, 4.560273, 4.552354, 4.533133, 4.546401, 
    4.541167, 4.553624, 4.561552, 4.557629, 4.581873, 4.572437, 4.6223, 
    4.600777, 4.657029, 4.643526, 4.660269, 4.65172, 4.666376, 4.653184, 
    4.676049, 4.681039, 4.677629, 4.690734, 4.652454, 4.667131, 4.557519, 
    4.558159, 4.561139, 4.54805, 4.54725, 4.535278, 4.545929, 4.55047, 
    4.562011, 4.568848, 4.575353, 4.589678, 4.605715, 4.628201, 4.644401, 
    4.655281, 4.648607, 4.654499, 4.647913, 4.644828, 4.679169, 4.659866, 
    4.688848, 4.687241, 4.674113, 4.687422, 4.558608, 4.554928, 4.54217, 
    4.552152, 4.533976, 4.544145, 4.549999, 4.572636, 4.577618, 4.582243, 
    4.591386, 4.603139, 4.623806, 4.641838, 4.658339, 4.657128, 4.657555, 
    4.661246, 4.652106, 4.662748, 4.664536, 4.659863, 4.687026, 4.679255, 
    4.687206, 4.682146, 4.556124, 4.562318, 4.55897, 4.565267, 4.560831, 
    4.580582, 4.586514, 4.614345, 4.602908, 4.621117, 4.604754, 4.607651, 
    4.621715, 4.605637, 4.640843, 4.616958, 4.66139, 4.637469, 4.662892, 
    4.658267, 4.665925, 4.672791, 4.681437, 4.697421, 4.693717, 4.707103, 
    4.571562, 4.579617, 4.578906, 4.587343, 4.59359, 4.60715, 4.628954, 
    4.620746, 4.635821, 4.638853, 4.615952, 4.630004, 4.585011, 4.592262, 
    4.587943, 4.572198, 4.622639, 4.596706, 4.644669, 4.630562, 4.671812, 
    4.651268, 4.691678, 4.709027, 4.725387, 4.74456, 4.584015, 4.578537, 
    4.588347, 4.601945, 4.614583, 4.631422, 4.633147, 4.636307, 4.644499, 
    4.651395, 4.637308, 4.653124, 4.593947, 4.624894, 4.576469, 4.591016, 
    4.601142, 4.596697, 4.619809, 4.625268, 4.647497, 4.635996, 4.704742, 
    4.674244, 4.759188, 4.735351, 4.576625, 4.583995, 4.609712, 4.597464, 
    4.632547, 4.641211, 4.648261, 4.657286, 4.65826, 4.663613, 4.654843, 
    4.663266, 4.631458, 4.645654, 4.606766, 4.616211, 4.611864, 4.6071, 
    4.621815, 4.63753, 4.637864, 4.642911, 4.657158, 4.632689, 4.708693, 
    4.661662, 4.592041, 4.606281, 4.608315, 4.602794, 4.640342, 4.626713, 
    4.663483, 4.653525, 4.669847, 4.661732, 4.660539, 4.650131, 4.643661, 
    4.627338, 4.614086, 4.603594, 4.606032, 4.617562, 4.638492, 4.65835, 
    4.653995, 4.668605, 4.629997, 4.646161, 4.63991, 4.656221, 4.620529, 
    4.650918, 4.612783, 4.616118, 4.626443, 4.64726, 4.651871, 4.656802, 
    4.653759, 4.639024, 4.636611, 4.626192, 4.623318, 4.615392, 4.608837, 
    4.614826, 4.621121, 4.639029, 4.655208, 4.672889, 4.677222, 4.697956, 
    4.681077, 4.708956, 4.685251, 4.726333, 4.652679, 4.68455, 4.626913, 
    4.633099, 4.644304, 4.670067, 4.656144, 4.672429, 4.636517, 4.617961, 
    4.613165, 4.604232, 4.61337, 4.612626, 4.621381, 4.618566, 4.639624, 
    4.628304, 4.66051, 4.672299, 4.705699, 4.726254, 4.747232, 4.756515, 
    4.759342, 4.760524,
  5.626039, 5.649297, 5.644769, 5.66357, 5.653134, 5.665454, 5.630748, 
    5.650223, 5.637784, 5.628129, 5.700191, 5.66441, 5.737524, 5.714577, 
    5.772345, 5.73395, 5.780109, 5.771232, 5.797972, 5.790303, 5.824607, 
    5.801515, 5.842442, 5.819085, 5.822735, 5.800755, 5.671595, 5.695728, 
    5.670168, 5.673604, 5.672061, 5.653351, 5.64394, 5.624263, 5.627831, 
    5.642285, 5.675149, 5.663976, 5.692163, 5.691525, 5.723025, 5.708807, 
    5.761939, 5.746801, 5.790622, 5.77958, 5.790104, 5.786911, 5.790145, 
    5.773956, 5.780889, 5.766656, 5.711468, 5.727648, 5.679491, 5.650682, 
    5.631601, 5.618092, 5.62, 5.62364, 5.642369, 5.660018, 5.673497, 
    5.682526, 5.691433, 5.718462, 5.732801, 5.765005, 5.759181, 5.769048, 
    5.778482, 5.794349, 5.791735, 5.798733, 5.768785, 5.788677, 5.755867, 
    5.764827, 5.693865, 5.666988, 5.6556, 5.64564, 5.621468, 5.638153, 
    5.631571, 5.647237, 5.657208, 5.652275, 5.682773, 5.670902, 5.733652, 
    5.706561, 5.777381, 5.760376, 5.781462, 5.770695, 5.789153, 5.772539, 
    5.801339, 5.807625, 5.803329, 5.81984, 5.771619, 5.790105, 5.652137, 
    5.652941, 5.65669, 5.640227, 5.639221, 5.624166, 5.637559, 5.643271, 
    5.657786, 5.666387, 5.674571, 5.692595, 5.712776, 5.741081, 5.761477, 
    5.775179, 5.766774, 5.774194, 5.7659, 5.762015, 5.805269, 5.780953, 
    5.817463, 5.815438, 5.7989, 5.815666, 5.653506, 5.648878, 5.632832, 
    5.645386, 5.622528, 5.635315, 5.642679, 5.671152, 5.67742, 5.683239, 
    5.694743, 5.709534, 5.735547, 5.75825, 5.77903, 5.777506, 5.778043, 
    5.782693, 5.771181, 5.784584, 5.786837, 5.78095, 5.815167, 5.805377, 
    5.815395, 5.809019, 5.650382, 5.658173, 5.653962, 5.661882, 5.656302, 
    5.681149, 5.688613, 5.723638, 5.709242, 5.732163, 5.711567, 5.715213, 
    5.732915, 5.712678, 5.756999, 5.726927, 5.782874, 5.752749, 5.784765, 
    5.778941, 5.788586, 5.797235, 5.808127, 5.828266, 5.823598, 5.840467, 
    5.669801, 5.679934, 5.67904, 5.689656, 5.697517, 5.714581, 5.742029, 
    5.731696, 5.750675, 5.754491, 5.72566, 5.743351, 5.686722, 5.695845, 
    5.690411, 5.670601, 5.734078, 5.701437, 5.761815, 5.744053, 5.796001, 
    5.770126, 5.82103, 5.842893, 5.863514, 5.887687, 5.685468, 5.678577, 
    5.690919, 5.708031, 5.723937, 5.745136, 5.747307, 5.751287, 5.761601, 
    5.770285, 5.752547, 5.772463, 5.697966, 5.736917, 5.675974, 5.694278, 
    5.70702, 5.701427, 5.730515, 5.737388, 5.765376, 5.750895, 5.837492, 
    5.799065, 5.906134, 5.876075, 5.676171, 5.685444, 5.717806, 5.702391, 
    5.746552, 5.757461, 5.766339, 5.777705, 5.778931, 5.785674, 5.774628, 
    5.785236, 5.745181, 5.763056, 5.714098, 5.725987, 5.720515, 5.714518, 
    5.733041, 5.752826, 5.753247, 5.759602, 5.777543, 5.746732, 5.842471, 
    5.783216, 5.695569, 5.713488, 5.716048, 5.709099, 5.756367, 5.739208, 
    5.785509, 5.772968, 5.793526, 5.783304, 5.781801, 5.768694, 5.760545, 
    5.739994, 5.723311, 5.710106, 5.713175, 5.727687, 5.754037, 5.779044, 
    5.77356, 5.791961, 5.743342, 5.763694, 5.755823, 5.776363, 5.731422, 
    5.769684, 5.721673, 5.72587, 5.738868, 5.765079, 5.770885, 5.777094, 
    5.773262, 5.754707, 5.75167, 5.738551, 5.734934, 5.724956, 5.716706, 
    5.724244, 5.732168, 5.754714, 5.775087, 5.797358, 5.802817, 5.82894, 
    5.807672, 5.842803, 5.812931, 5.864706, 5.771903, 5.812049, 5.739459, 
    5.747247, 5.761355, 5.793803, 5.776267, 5.796778, 5.751551, 5.72819, 
    5.722154, 5.710909, 5.722411, 5.721475, 5.732495, 5.728951, 5.755463, 
    5.741211, 5.781765, 5.796615, 5.838698, 5.864606, 5.891056, 5.902761, 
    5.906327, 5.907819,
  8.094118, 8.128306, 8.12165, 8.149295, 8.133948, 8.152065, 8.101038, 
    8.129667, 8.111381, 8.097189, 8.203166, 8.150529, 8.258118, 8.224336, 
    8.309403, 8.252855, 8.320842, 8.307764, 8.347167, 8.335863, 8.386434, 
    8.352388, 8.412737, 8.37829, 8.383674, 8.351268, 8.161097, 8.196599, 
    8.158998, 8.164051, 8.161782, 8.134267, 8.120432, 8.091507, 8.096751, 
    8.117997, 8.166325, 8.149891, 8.191352, 8.190413, 8.236772, 8.215843, 
    8.294074, 8.271778, 8.336335, 8.320062, 8.33557, 8.330865, 8.335631, 
    8.311776, 8.321991, 8.301023, 8.21976, 8.243577, 8.17271, 8.130343, 
    8.102293, 8.082438, 8.085243, 8.090592, 8.118122, 8.144072, 8.163894, 
    8.177176, 8.190279, 8.230056, 8.251163, 8.29859, 8.290011, 8.304545, 
    8.318444, 8.341826, 8.337974, 8.348289, 8.304159, 8.333468, 8.285129, 
    8.298328, 8.193857, 8.154321, 8.137574, 8.12293, 8.0874, 8.111923, 
    8.102249, 8.125278, 8.139939, 8.132685, 8.177539, 8.160077, 8.252416, 
    8.212539, 8.316822, 8.291771, 8.322835, 8.306972, 8.334169, 8.309689, 
    8.352129, 8.361395, 8.355062, 8.379404, 8.308333, 8.335571, 8.132482, 
    8.133665, 8.139176, 8.114973, 8.113493, 8.091364, 8.111052, 8.119448, 
    8.140789, 8.153437, 8.165473, 8.191988, 8.221685, 8.263354, 8.293393, 
    8.313579, 8.301196, 8.312127, 8.299909, 8.294186, 8.357923, 8.322086, 
    8.375899, 8.372914, 8.348535, 8.373251, 8.134496, 8.12769, 8.104102, 
    8.122557, 8.088957, 8.107752, 8.118576, 8.160445, 8.169664, 8.178225, 
    8.195149, 8.216914, 8.255207, 8.28864, 8.319253, 8.317007, 8.317798, 
    8.324649, 8.307688, 8.327436, 8.330756, 8.322081, 8.372515, 8.358081, 
    8.37285, 8.36345, 8.129901, 8.141356, 8.135165, 8.146812, 8.138606, 
    8.175149, 8.186131, 8.237674, 8.216486, 8.250224, 8.219907, 8.225273, 
    8.251332, 8.221541, 8.286797, 8.242516, 8.324916, 8.280539, 8.327703, 
    8.31912, 8.333333, 8.34608, 8.362136, 8.391829, 8.384945, 8.409823, 
    8.158458, 8.173363, 8.172048, 8.187665, 8.199231, 8.224343, 8.264751, 
    8.249537, 8.277483, 8.283104, 8.240651, 8.266698, 8.183348, 8.196771, 
    8.188775, 8.159635, 8.253044, 8.205, 8.293891, 8.267732, 8.344262, 
    8.306134, 8.381158, 8.413401, 8.443824, 8.479502, 8.181503, 8.171366, 
    8.189523, 8.214703, 8.238114, 8.269326, 8.272523, 8.278383, 8.293576, 
    8.306368, 8.28024, 8.309577, 8.199891, 8.257224, 8.167538, 8.194465, 
    8.213216, 8.204983, 8.247799, 8.257916, 8.299136, 8.277806, 8.405437, 
    8.348778, 8.506738, 8.46236, 8.167827, 8.181468, 8.22909, 8.206403, 
    8.271412, 8.287477, 8.300555, 8.3173, 8.319107, 8.329042, 8.312767, 
    8.328398, 8.269392, 8.295719, 8.223632, 8.241133, 8.233077, 8.22425, 
    8.251517, 8.280651, 8.281271, 8.290631, 8.317061, 8.271676, 8.412779, 
    8.325419, 8.196363, 8.222733, 8.226501, 8.216275, 8.285866, 8.260596, 
    8.328799, 8.310322, 8.340613, 8.32555, 8.323336, 8.304025, 8.292021, 
    8.261755, 8.237193, 8.217757, 8.222273, 8.243635, 8.282435, 8.319272, 
    8.311193, 8.338308, 8.266685, 8.296659, 8.285065, 8.315323, 8.249133, 
    8.305483, 8.234781, 8.240959, 8.260096, 8.298698, 8.307252, 8.316401, 
    8.310754, 8.283422, 8.278949, 8.259629, 8.254304, 8.239614, 8.227469, 
    8.238565, 8.250232, 8.283431, 8.313443, 8.346262, 8.354307, 8.392823, 
    8.361465, 8.413268, 8.369218, 8.445583, 8.308752, 8.367917, 8.260966, 
    8.272434, 8.293214, 8.341022, 8.315181, 8.345407, 8.278773, 8.244374, 
    8.235489, 8.218939, 8.235868, 8.234489, 8.250712, 8.245497, 8.284535, 
    8.263547, 8.323281, 8.345167, 8.407215, 8.445436, 8.484475, 8.501758, 
    8.507023, 8.509225,
  12.66552, 12.72099, 12.71019, 12.75506, 12.73015, 12.75956, 12.67674, 
    12.7232, 12.69352, 12.6705, 12.84257, 12.75706, 12.93193, 12.87698, 
    13.01541, 12.92337, 13.03404, 13.01274, 13.07694, 13.05852, 13.14096, 
    13.08545, 13.18388, 13.12768, 13.13646, 13.08362, 12.77422, 12.83189, 
    12.77081, 12.77902, 12.77534, 12.73066, 12.70821, 12.66129, 12.66979, 
    12.70426, 12.78271, 12.75603, 12.82337, 12.82185, 12.8972, 12.86318, 
    12.99045, 12.95416, 13.05929, 13.03277, 13.05804, 13.05037, 13.05814, 
    13.01928, 13.03592, 13.00176, 12.86954, 12.90827, 12.79309, 12.72429, 
    12.67878, 12.64658, 12.65113, 12.6598, 12.70446, 12.74658, 12.77876, 
    12.80034, 12.82163, 12.88628, 12.92061, 12.9978, 12.98384, 13.0075, 
    13.03014, 13.06824, 13.06196, 13.07877, 13.00687, 13.05462, 12.97589, 
    12.99738, 12.82744, 12.76322, 12.73603, 12.71226, 12.65462, 12.6944, 
    12.67871, 12.71607, 12.73987, 12.72809, 12.80093, 12.77257, 12.92265, 
    12.8578, 13.0275, 12.9867, 13.03729, 13.01145, 13.05576, 13.01588, 
    13.08503, 13.10013, 13.08981, 13.1295, 13.01367, 13.05804, 12.72777, 
    12.72968, 12.73863, 12.69935, 12.69695, 12.66105, 12.69299, 12.70661, 
    12.74125, 12.76178, 12.78133, 12.8244, 12.87267, 12.94045, 12.98934, 
    13.02221, 13.00205, 13.01985, 12.99995, 12.99063, 13.09447, 13.03607, 
    13.12378, 13.11891, 13.07917, 13.11946, 12.73103, 12.71999, 12.68172, 
    12.71166, 12.65715, 12.68764, 12.7052, 12.77316, 12.78814, 12.80204, 
    12.82954, 12.86492, 12.92719, 12.9816, 13.03146, 13.0278, 13.02909, 
    13.04025, 13.01262, 13.04479, 13.0502, 13.03606, 13.11826, 13.09473, 
    13.11881, 13.10348, 12.72358, 12.74217, 12.73212, 12.75103, 12.73771, 
    12.79704, 12.81489, 12.89867, 12.86422, 12.91909, 12.86978, 12.87851, 
    12.92089, 12.87244, 12.9786, 12.90655, 13.04068, 12.96841, 13.04522, 
    13.03124, 13.05439, 13.07517, 13.10134, 13.14977, 13.13854, 13.17913, 
    12.76994, 12.79414, 12.79201, 12.81738, 12.83617, 12.87699, 12.94272, 
    12.91797, 12.96344, 12.97259, 12.90351, 12.94589, 12.81037, 12.83218, 
    12.81918, 12.77185, 12.92367, 12.84555, 12.99015, 12.94757, 13.0722, 
    13.01009, 13.13236, 13.18496, 13.23463, 13.29292, 12.80737, 12.7909, 
    12.8204, 12.86132, 12.89939, 12.95017, 12.95537, 12.96491, 12.98964, 
    13.01047, 12.96793, 13.0157, 12.83725, 12.93047, 12.78468, 12.82843, 
    12.8589, 12.84552, 12.91514, 12.9316, 12.99869, 12.96397, 13.17197, 
    13.07957, 13.33744, 13.26491, 12.78515, 12.80731, 12.88471, 12.84783, 
    12.95356, 12.97971, 13.001, 13.02827, 13.03122, 13.0474, 13.02089, 
    13.04635, 12.95027, 12.99313, 12.87584, 12.9043, 12.8912, 12.87684, 
    12.92119, 12.9686, 12.96961, 12.98484, 13.02789, 12.95399, 13.18395, 
    13.0415, 12.83151, 12.87438, 12.8805, 12.86388, 12.97709, 12.93596, 
    13.04701, 13.01691, 13.06626, 13.04171, 13.03811, 13.00665, 12.98711, 
    12.93785, 12.89789, 12.86629, 12.87363, 12.90837, 12.9715, 13.03149, 
    13.01833, 13.0625, 12.94587, 12.99466, 12.97578, 13.02505, 12.91731, 
    13.00903, 12.89397, 12.90402, 12.93515, 12.99798, 13.01191, 13.02681, 
    13.01761, 12.97311, 12.96583, 12.93439, 12.92572, 12.90183, 12.88208, 
    12.90012, 12.9191, 12.97312, 13.02199, 13.07546, 13.08858, 13.15139, 
    13.10025, 13.18475, 13.11289, 13.2375, 13.01435, 13.11077, 12.93656, 
    12.95522, 12.98905, 13.06693, 13.02482, 13.07407, 12.96554, 12.90957, 
    12.89512, 12.86821, 12.89573, 12.89349, 12.91988, 12.9114, 12.97492, 
    12.94076, 13.03802, 13.07368, 13.17487, 13.23726, 13.30105, 13.3293, 
    13.33791, 13.34151,
  20.5999, 20.69597, 20.67725, 20.75504, 20.71184, 20.76284, 20.61933, 
    20.6998, 20.64839, 20.60852, 20.90694, 20.75851, 21.06236, 20.96676, 
    21.20783, 21.04745, 21.24033, 21.20317, 21.31522, 21.28305, 21.42712, 
    21.33008, 21.50222, 21.40389, 21.41924, 21.32689, 20.78828, 20.8884, 
    20.78236, 20.7966, 20.79021, 20.71274, 20.67383, 20.59257, 20.6073, 
    20.66698, 20.80301, 20.75671, 20.87359, 20.87094, 21.00193, 20.94276, 
    21.1643, 21.10106, 21.28439, 21.23812, 21.28222, 21.26883, 21.28239, 
    21.21457, 21.2436, 21.18403, 20.95382, 21.02119, 20.82101, 20.7017, 
    20.62286, 20.56712, 20.57499, 20.59, 20.66733, 20.74033, 20.79616, 
    20.8336, 20.87056, 20.98293, 21.04266, 21.17712, 21.15278, 21.19403, 
    21.23352, 21.30001, 21.28905, 21.31841, 21.19294, 21.27624, 21.13892, 
    21.17638, 20.88066, 20.76919, 20.72204, 20.68085, 20.58105, 20.64991, 
    20.62273, 20.68745, 20.7287, 20.70829, 20.83462, 20.78541, 21.04621, 
    20.93342, 21.22891, 21.15777, 21.246, 21.20092, 21.27823, 21.20864, 
    21.32934, 21.35573, 21.3377, 21.40707, 21.20479, 21.28222, 20.70772, 
    20.71104, 20.72655, 20.65848, 20.65433, 20.59217, 20.64746, 20.67106, 
    20.73109, 20.7667, 20.80061, 20.87539, 20.95927, 21.07719, 21.16237, 
    21.21969, 21.18452, 21.21557, 21.18087, 21.16462, 21.34584, 21.24387, 
    21.39707, 21.38856, 21.31911, 21.38952, 20.71338, 20.69424, 20.62794, 
    20.6798, 20.58541, 20.63819, 20.66861, 20.78644, 20.81242, 20.83656, 
    20.88431, 20.94578, 21.05411, 21.14888, 21.23582, 21.22943, 21.23168, 
    21.25116, 21.20296, 21.25908, 21.26852, 21.24385, 21.38742, 21.34629, 
    21.38838, 21.36159, 20.70046, 20.73269, 20.71527, 20.74804, 20.72495, 
    20.82788, 20.85886, 21.00448, 20.94457, 21.04, 20.95424, 20.96941, 
    21.04314, 20.95886, 21.14365, 21.01818, 21.25191, 21.1259, 21.25984, 
    21.23544, 21.27585, 21.31212, 21.35784, 21.44251, 21.42287, 21.4939, 
    20.78084, 20.82285, 20.81914, 20.86319, 20.89583, 20.96678, 21.08115, 
    21.03806, 21.11724, 21.13318, 21.01291, 21.08667, 20.85101, 20.88889, 
    20.86632, 20.78416, 21.04799, 20.91212, 21.16379, 21.0896, 21.30695, 
    21.19854, 21.41207, 21.50412, 21.59113, 21.69336, 20.84581, 20.81722, 
    20.86843, 20.93953, 21.00573, 21.09411, 21.10318, 21.11979, 21.16289, 
    21.19921, 21.12506, 21.20832, 20.8977, 21.05983, 20.80643, 20.88238, 
    20.93533, 20.91208, 21.03314, 21.06179, 21.17867, 21.11815, 21.48136, 
    21.3198, 21.77155, 21.64422, 20.80724, 20.84571, 20.9802, 20.91608, 
    21.10003, 21.14559, 21.1827, 21.23026, 21.2354, 21.26365, 21.21739, 
    21.26181, 21.0943, 21.16897, 20.96477, 21.01427, 20.99148, 20.96652, 
    21.04366, 21.12622, 21.12798, 21.15453, 21.22959, 21.10077, 21.50234, 
    21.25335, 20.88774, 20.96223, 20.97288, 20.94398, 21.14101, 21.06938, 
    21.26296, 21.21044, 21.29656, 21.25372, 21.24742, 21.19255, 21.15848, 
    21.07266, 21.00312, 20.94816, 20.96093, 21.02135, 21.13128, 21.23587, 
    21.21291, 21.29, 21.08663, 21.17164, 21.13874, 21.22465, 21.03692, 
    21.1967, 20.9963, 21.01378, 21.06796, 21.17743, 21.20172, 21.22771, 
    21.21167, 21.13408, 21.12139, 21.06664, 21.05156, 21.00997, 20.97562, 
    21.00701, 21.04003, 21.13411, 21.21931, 21.31264, 21.33555, 21.44535, 
    21.35593, 21.50374, 21.37803, 21.59616, 21.20598, 21.37432, 21.07043, 
    21.10292, 21.16186, 21.29773, 21.22425, 21.31021, 21.1209, 21.02345, 
    20.9983, 20.9515, 20.99937, 20.99547, 21.04139, 21.02662, 21.13724, 
    21.07774, 21.24727, 21.30952, 21.48644, 21.59574, 21.70763, 21.75724, 
    21.77237, 21.7787,
  34.64178, 34.82256, 34.7873, 34.9339, 34.85246, 34.94862, 34.67832, 
    34.82977, 34.73297, 34.65799, 35.22099, 34.94046, 35.51581, 35.33433, 
    35.79281, 35.48749, 35.85484, 35.78393, 35.99794, 35.93644, 36.21229, 
    36.02638, 36.3565, 36.16775, 36.19719, 36.02028, 34.99663, 35.18589, 
    34.98547, 35.01235, 35.00028, 34.85415, 34.78085, 34.62801, 34.65569, 
    34.76797, 35.02445, 34.93707, 35.15787, 35.15286, 35.40105, 35.28883, 
    35.70983, 35.58942, 35.939, 35.85061, 35.93484, 35.90927, 35.93518, 
    35.80567, 35.86108, 35.74743, 35.30981, 35.43761, 35.05846, 34.83335, 
    34.68494, 34.5802, 34.59498, 34.62318, 34.76863, 34.90616, 35.01151, 
    35.08224, 35.15214, 35.365, 35.47839, 35.73426, 35.68786, 35.7665, 
    35.84183, 35.96887, 35.94791, 36.00405, 35.76441, 35.92341, 35.66148, 
    35.73284, 35.17124, 34.96061, 34.87169, 34.79408, 34.60635, 34.73584, 
    34.68471, 34.80651, 34.88423, 34.84576, 35.08418, 34.99121, 35.48513, 
    35.27114, 35.83303, 35.69738, 35.86566, 35.77964, 35.92722, 35.79436, 
    36.02497, 36.07548, 36.04095, 36.17384, 35.78702, 35.93485, 34.84468, 
    34.85096, 34.88018, 34.75196, 34.74414, 34.62726, 34.73122, 34.77564, 
    34.88874, 34.9559, 35.01992, 35.16127, 35.32013, 35.54402, 35.70615, 
    35.81544, 35.74836, 35.80758, 35.74139, 35.71043, 36.05655, 35.8616, 
    36.15468, 36.13837, 36.00539, 36.14021, 34.85536, 34.81929, 34.6945, 
    34.7921, 34.61456, 34.71379, 34.77103, 34.99316, 35.04223, 35.08784, 
    35.17815, 35.29456, 35.50015, 35.68045, 35.84622, 35.83403, 35.83833, 
    35.87551, 35.78352, 35.89064, 35.90867, 35.86156, 36.13618, 36.05741, 
    36.13802, 36.0867, 34.83101, 34.89175, 34.85891, 34.92071, 34.87716, 
    35.07145, 35.13, 35.4059, 35.29227, 35.47334, 35.31059, 35.33936, 
    35.4793, 35.31936, 35.67049, 35.4319, 35.87695, 35.63669, 35.89209, 
    35.8455, 35.92268, 35.99202, 36.07952, 36.24184, 36.20415, 36.3405, 
    34.9826, 35.06193, 35.05492, 35.13819, 35.19995, 35.33437, 35.55154, 
    35.46964, 35.6202, 35.65054, 35.42189, 35.56203, 35.11515, 35.18681, 
    35.14411, 34.98885, 35.48851, 35.2308, 35.70884, 35.5676, 35.98212, 
    35.7751, 36.18343, 36.36015, 36.52758, 36.7248, 35.10532, 35.05129, 
    35.14811, 35.28272, 35.40826, 35.5762, 35.59344, 35.62506, 35.70713, 
    35.77637, 35.63508, 35.79375, 35.20348, 35.511, 35.03091, 35.17449, 
    35.27476, 35.23071, 35.4603, 35.51473, 35.73722, 35.62194, 36.31643, 
    36.00671, 36.876, 36.62993, 35.03245, 35.10513, 35.35983, 35.2383, 
    35.58744, 35.67417, 35.74489, 35.83562, 35.84542, 35.89936, 35.81104, 
    35.89586, 35.57656, 35.71873, 35.33056, 35.42447, 35.38122, 35.33387, 
    35.4803, 35.6373, 35.64064, 35.69121, 35.83433, 35.58887, 36.35673, 
    35.87968, 35.18464, 35.32574, 35.34594, 35.29114, 35.66546, 35.52916, 
    35.89804, 35.79779, 35.96227, 35.8804, 35.86838, 35.76368, 35.69873, 
    35.5354, 35.40332, 35.29908, 35.32327, 35.43792, 35.64693, 35.84632, 
    35.80251, 35.94973, 35.56196, 35.72381, 35.66113, 35.8249, 35.46748, 
    35.77157, 35.39036, 35.42354, 35.52647, 35.73484, 35.78116, 35.83075, 
    35.80013, 35.65226, 35.62811, 35.52395, 35.49529, 35.41631, 35.35114, 
    35.41068, 35.47338, 35.65231, 35.81471, 35.99301, 36.03684, 36.24728, 
    36.07586, 36.35942, 36.11818, 36.53728, 35.78928, 36.11108, 35.53115, 
    35.59296, 35.70518, 35.96449, 35.82413, 35.98836, 35.62716, 35.44189, 
    35.39416, 35.3054, 35.39619, 35.3888, 35.47597, 35.44792, 35.65827, 
    35.54505, 35.86808, 35.98705, 36.32619, 36.53647, 36.75238, 36.84832, 
    36.87759, 36.88984,
  60.67866, 61.07138, 60.99464, 61.31427, 61.13654, 61.34644, 60.75787, 
    61.08709, 60.87651, 60.71379, 61.94415, 61.3286, 62.59654, 62.19429, 
    63.21474, 62.53363, 63.35389, 63.19484, 63.67592, 63.53733, 64.16097, 
    63.74009, 64.48915, 64.05992, 64.12669, 63.72631, 61.45146, 61.86686, 
    61.42703, 61.48588, 61.45945, 61.14022, 60.9806, 60.64882, 60.70879, 
    60.95258, 61.51238, 61.32119, 61.80522, 61.7942, 62.34192, 62.09377, 
    63.02899, 62.76031, 63.54311, 63.34439, 63.53375, 63.4762, 63.5345, 
    63.24357, 63.36789, 63.11309, 62.1401, 62.42293, 61.58691, 61.09489, 
    60.77224, 60.54533, 60.5773, 60.63837, 60.95401, 61.2537, 61.48405, 
    61.6391, 61.79262, 62.26212, 62.51342, 63.08363, 62.97991, 63.15579, 
    63.32469, 63.61038, 63.56317, 63.68969, 63.15111, 63.50803, 62.92099, 
    63.08046, 61.83464, 61.37265, 61.17847, 61.00938, 60.60192, 60.88274, 
    60.77174, 61.03644, 61.20583, 61.12193, 61.64335, 61.4396, 62.52837, 
    62.05472, 63.30494, 63.00117, 63.37819, 63.18523, 63.5166, 63.21821, 
    63.7369, 63.85101, 63.77299, 64.07372, 63.20175, 63.53376, 61.11959, 
    61.13326, 61.197, 60.91779, 60.90078, 60.64719, 60.87272, 60.96927, 
    61.21567, 61.36237, 61.50245, 61.81269, 62.16289, 62.65925, 63.02077, 
    63.26548, 63.11519, 63.24784, 63.0996, 63.03035, 63.80822, 63.36906, 
    64.03029, 63.99333, 63.69271, 63.99749, 61.14286, 61.06427, 60.79298, 
    61.00508, 60.61969, 60.83485, 60.95924, 61.44387, 61.55134, 61.65136, 
    61.84983, 62.10643, 62.56173, 62.96335, 63.33453, 63.30719, 63.31681, 
    63.40031, 63.19391, 63.43432, 63.47487, 63.36899, 63.98838, 63.81017, 
    63.99254, 63.87637, 61.08979, 61.22225, 61.1506, 61.28547, 61.19041, 
    61.6154, 61.74396, 62.35265, 62.10136, 62.5022, 62.14183, 62.20539, 
    62.51543, 62.16119, 62.9411, 62.41028, 63.40356, 62.86567, 63.43758, 
    63.33292, 63.50638, 63.66257, 63.86015, 64.22809, 64.14249, 64.45267, 
    61.42075, 61.59453, 61.57916, 61.76195, 61.89783, 62.19437, 62.67599, 
    62.494, 62.8289, 62.89658, 62.38808, 62.69933, 61.71135, 61.86889, 
    61.77497, 61.43444, 62.53588, 61.96577, 63.02679, 62.71174, 63.64025, 
    63.17506, 64.09548, 64.49747, 64.88044, 65.3342, 61.68975, 61.57121, 
    61.78375, 62.08028, 62.35789, 62.73087, 62.76927, 62.83974, 63.02298, 
    63.1779, 62.86208, 63.21685, 61.9056, 62.58585, 61.52654, 61.84178, 
    62.06271, 61.96557, 62.47326, 62.59414, 63.09025, 62.83279, 64.3978, 
    63.6957, 65.68405, 65.11556, 61.5299, 61.68932, 62.25066, 61.98231, 
    62.75591, 62.94933, 63.10743, 63.31075, 63.33276, 63.45393, 63.25561, 
    63.44606, 62.73167, 63.04889, 62.18595, 62.39381, 62.298, 62.19328, 
    62.51765, 62.86703, 62.87449, 62.9874, 63.30784, 62.75908, 64.48967, 
    63.4097, 61.8641, 62.17531, 62.21996, 62.09887, 62.92989, 62.62622, 
    63.45097, 63.22589, 63.59551, 63.4113, 63.38429, 63.14947, 63.00418, 
    62.64008, 62.34694, 62.1164, 62.16985, 62.42362, 62.88852, 63.33477, 
    63.23648, 63.56726, 62.69917, 63.06026, 62.92022, 63.2867, 62.48919, 
    63.16716, 62.31825, 62.39175, 62.62022, 63.08494, 63.18863, 63.29981, 
    63.23115, 62.90041, 62.84653, 62.61464, 62.55093, 62.37573, 62.23145, 
    62.36326, 62.5023, 62.90052, 63.26383, 63.6648, 63.7637, 64.24046, 
    63.85188, 64.4958, 63.9476, 64.90269, 63.20683, 63.93153, 62.63064, 
    62.7682, 63.0186, 63.60052, 63.28497, 63.6543, 62.84442, 62.43243, 
    62.32666, 62.13037, 62.33117, 62.31479, 62.50804, 62.4458, 62.91383, 
    62.66155, 63.38363, 63.65136, 64.42004, 64.90083, 65.39787, 65.61987, 
    65.68774, 65.71616,
  116.3177, 117.5456, 117.3041, 118.3152, 117.7513, 118.4177, 116.5638, 
    117.5952, 116.9339, 116.4268, 120.3482, 118.3608, 122.5137, 121.1711, 
    124.6258, 122.3021, 125.1096, 124.5568, 126.2418, 125.7524, 127.9808, 
    126.4695, 129.1813, 127.6151, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9487, 118.3372, 119.895, 119.8592, 121.661, 120.8393, 
    123.9848, 123.0674, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7258, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9053, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3958, 122.2342, 124.1728, 123.8164, 124.4217, 
    125.0078, 126.01, 125.8434, 126.2906, 124.4056, 125.6494, 123.6147, 
    124.1619, 119.9907, 118.5013, 117.8839, 117.3505, 116.0801, 116.9533, 
    116.607, 117.4356, 117.9707, 117.7052, 119.3704, 118.7153, 122.2845, 
    120.7108, 124.9391, 123.8893, 125.1945, 124.5236, 125.6795, 124.6378, 
    126.4582, 126.8648, 126.5865, 127.6649, 124.5808, 125.7399, 117.6978, 
    117.741, 117.9427, 117.063, 117.0098, 116.2202, 116.922, 117.2245, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9566, 
    124.8018, 124.2816, 124.7406, 124.2278, 123.9895, 126.712, 125.1626, 
    127.5082, 127.3751, 126.3013, 127.3901, 117.7713, 117.5232, 116.6731, 
    117.337, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.881, 122.3966, 123.7596, 125.0421, 124.9469, 124.9804, 
    125.2718, 124.5536, 125.3908, 125.5329, 125.1623, 127.3573, 126.719, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9218, 
    119.2802, 119.696, 121.6967, 120.8643, 122.1966, 120.9977, 121.2078, 
    122.241, 121.0616, 123.6834, 121.889, 125.2831, 123.4258, 125.4022, 
    125.0365, 125.6436, 126.1945, 126.8974, 128.2247, 127.9138, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1968, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8149, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3097, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4884, 127.7436, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7949, 121.7142, 122.9675, 123.0978, 123.3374, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.014, 
    120.7371, 120.4183, 122.0996, 122.5056, 124.1956, 123.3137, 128.8452, 
    126.3119, 133.7281, 131.5293, 119.005, 119.5191, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2548, 124.9593, 125.0359, 125.4595, 124.7676, 
    125.4319, 122.9702, 124.0532, 121.1435, 121.834, 121.5149, 121.1677, 
    122.2484, 123.4304, 123.4559, 123.842, 124.9492, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1083, 121.256, 120.8561, 123.6451, 122.6137, 
    125.4491, 124.6645, 125.9575, 125.3102, 125.2158, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.043, 
    124.7011, 125.8578, 122.8602, 124.0923, 123.612, 124.8756, 122.153, 
    124.4611, 121.5822, 121.8271, 122.5935, 124.1773, 124.5353, 124.9212, 
    124.6827, 123.5443, 123.3605, 122.5747, 122.3602, 121.7737, 121.2941, 
    121.7321, 122.197, 123.5447, 124.7961, 126.2024, 126.5535, 128.2698, 
    126.8678, 129.2059, 127.2107, 130.7229, 124.5984, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9752, 124.8696, 126.1653, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5902, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6129, 133.4765, 
    133.7426, 133.8544,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02028661, -0.01995555, -0.02001946, -0.01975575, -0.01990158, 
    -0.01972957, -0.02021903, -0.01994251, -0.02011857, -0.02025658, 
    -0.01925455, -0.01974408, -0.01876002, -0.01906207, -0.01831312, 
    -0.01880666, -0.01821532, -0.0183272, -0.01799279, -0.01808791, 
    -0.01766731, -0.01794907, -0.01745352, -0.01773418, -0.01768994, 
    -0.01795844, -0.01964453, -0.01931477, -0.01966425, -0.01961681, 
    -0.01963809, -0.01989855, -0.02003119, -0.02031218, -0.02026086, 
    -0.02005464, -0.01959551, -0.01975011, -0.01936305, -0.0193717, 
    -0.01895016, -0.01913898, -0.01844525, -0.01863963, -0.01808393, 
    -0.01822197, -0.01809038, -0.01813018, -0.01808986, -0.01829278, 
    -0.01820554, -0.01838521, -0.01910346, -0.01888927, -0.01953586, 
    -0.01993605, -0.02020681, -0.02040132, -0.0203737, -0.02032115, 
    -0.02005344, -0.01980523, -0.01961828, -0.01949429, -0.01937295, 
    -0.01901049, -0.01882169, -0.0184062, -0.01848047, -0.01835486, 
    -0.01823577, -0.01803765, -0.0180701, -0.01798338, -0.01835819, 
    -0.01810815, -0.01852292, -0.01840846, -0.01933998, -0.01970828, 
    -0.019867, -0.02000715, -0.02035249, -0.02011332, -0.02020724, 
    -0.0199846, -0.01984449, -0.01991366, -0.01949091, -0.0196541, 
    -0.01881056, -0.01916902, -0.01824961, -0.0184652, -0.01819835, 
    -0.018334, -0.01810222, -0.01831068, -0.01795123, -0.01787397, 
    -0.01792673, -0.01772502, -0.0183223, -0.01809037, -0.0199156, 
    -0.01990429, -0.01985175, -0.02008383, -0.02009813, -0.02031358, 
    -0.02012176, -0.02004066, -0.01983641, -0.01971663, -0.01960349, 
    -0.01935719, -0.01908603, -0.01871374, -0.01845114, -0.01827735, 
    -0.01838371, -0.01828977, -0.01839482, -0.01844428, -0.01790287, 
    -0.01820472, -0.01775388, -0.01777851, -0.01798132, -0.01777573, 
    -0.01989637, -0.01996146, -0.0201892, -0.02001074, -0.02033719, 
    -0.02015374, -0.02004906, -0.01965065, -0.01956429, -0.01948454, 
    -0.01932809, -0.01912927, -0.0187858, -0.01849238, -0.01822887, 
    -0.01824804, -0.01824128, -0.01818292, -0.01832785, -0.01815925, 
    -0.0181311, -0.01820477, -0.01778181, -0.01790155, -0.01777903, 
    -0.01785689, -0.01994028, -0.01983101, -0.01988997, -0.01977925, 
    -0.01985718, -0.01951315, -0.01941125, -0.01894207, -0.01913316, 
    -0.01883004, -0.01910214, -0.01905361, -0.01882019, -0.01908733, 
    -0.01850841, -0.01889875, -0.01818066, -0.01856294, -0.01815698, 
    -0.01823, -0.01810929, -0.01800191, -0.01786781, -0.01762318, 
    -0.01767951, -0.01747704, -0.01966932, -0.01952978, -0.01954205, 
    -0.01939707, -0.0192906, -0.01906201, -0.01870143, -0.01883616, 
    -0.01858964, -0.01854056, -0.01891541, -0.01868428, -0.01943701, 
    -0.01931319, -0.01938682, -0.01965826, -0.01880499, -0.01923778, 
    -0.01844683, -0.01867518, -0.01801717, -0.0183412, -0.01771059, 
    -0.01744816, -0.01720512, -0.01692564, -0.0194541, -0.0195484, 
    -0.01937992, -0.01914935, -0.01893812, -0.01866116, -0.01863308, 
    -0.01858176, -0.01844956, -0.01833919, -0.01856555, -0.01831163, 
    -0.01928455, -0.01876793, -0.01958416, -0.01933439, -0.01916287, 
    -0.01923793, -0.01885163, -0.0187618, -0.01840148, -0.01858681, 
    -0.01751252, -0.01797928, -0.01671622, -0.01705918, -0.01958146, 
    -0.01945443, -0.01901919, -0.01922496, -0.01864284, -0.01850248, 
    -0.01838924, -0.01824554, -0.01823011, -0.01814562, -0.01828429, 
    -0.01815109, -0.01866058, -0.01843101, -0.01906843, -0.01891111, 
    -0.01898332, -0.01906284, -0.01881855, -0.01856195, -0.01855655, 
    -0.01847509, -0.01824757, -0.01864052, -0.01745318, -0.01817637, 
    -0.01931693, -0.01907655, -0.01904252, -0.01913507, -0.0185165, 
    -0.01873809, -0.01814768, -0.01830525, -0.01804786, -0.01817526, 
    -0.01819409, -0.01835935, -0.01846304, -0.01872787, -0.01894637, 
    -0.01912162, -0.01908072, -0.01888875, -0.01854639, -0.0182287, 
    -0.01829778, -0.01806728, -0.0186844, -0.01842288, -0.01852348, 
    -0.01826242, -0.01883974, -0.01834679, -0.01896801, -0.01891266, 
    -0.01874252, -0.01840526, -0.01833159, -0.01825322, -0.01830154, 
    -0.01853779, -0.01857683, -0.01874665, -0.01879381, -0.0189247, 
    -0.01903379, -0.01893408, -0.01882997, -0.01853771, -0.0182785, 
    -0.01800038, -0.01793303, -0.01761506, -0.01787339, -0.01744924, 
    -0.01780907, -0.01719121, -0.01831871, -0.01781984, -0.01873483, 
    -0.01863387, -0.0184527, -0.01804441, -0.01826364, -0.01800755, 
    -0.01857836, -0.01888215, -0.01896166, -0.01911091, -0.01895826, 
    -0.01897063, -0.01882569, -0.01887214, -0.01852809, -0.01871205, 
    -0.01819455, -0.01800957, -0.01749812, -0.01719238, -0.01688715, 
    -0.01675426, -0.01671404, -0.01669725,
  -0.05424561, -0.05319658, -0.05339885, -0.05256495, -0.05302586, 
    -0.05248226, -0.05403123, -0.05315533, -0.05371277, -0.05415035, 
    -0.05098546, -0.05252808, -0.04943406, -0.05038077, -0.04803829, 
    -0.04958008, -0.04773362, -0.04808215, -0.04704147, -0.04733715, 
    -0.04603188, -0.04690566, -0.04537049, -0.04623903, -0.04610197, 
    -0.04693477, -0.05221383, -0.05117485, -0.05227605, -0.05212636, 
    -0.0521935, -0.05301626, -0.05343598, -0.05432675, -0.0541639, 
    -0.05351026, -0.0520592, -0.05254713, -0.05132678, -0.05135401, 
    -0.05002971, -0.05062228, -0.04845035, -0.04905746, -0.04732477, 
    -0.04775432, -0.04734484, -0.04746862, -0.04734323, -0.04797489, 
    -0.04770316, -0.04826302, -0.05051072, -0.04983884, -0.05187109, 
    -0.05313487, -0.05399247, -0.0546098, -0.05452207, -0.05435523, 
    -0.05350646, -0.05272127, -0.05213102, -0.05174008, -0.05135792, 
    -0.05021893, -0.04962715, -0.0483285, -0.04856027, -0.04816839, 
    -0.04779728, -0.04718089, -0.04728178, -0.04701226, -0.04817876, 
    -0.04740009, -0.04869279, -0.04833554, -0.05125417, -0.05241504, 
    -0.05291651, -0.05335989, -0.05445472, -0.05369613, -0.05399383, 
    -0.05328851, -0.05284534, -0.05306406, -0.05172944, -0.05224403, 
    -0.0495923, -0.05071663, -0.04784041, -0.04851261, -0.04768078, 
    -0.04810335, -0.04738167, -0.04803066, -0.04691239, -0.04667253, 
    -0.0468363, -0.04621063, -0.0480669, -0.04734481, -0.05307018, 
    -0.05303444, -0.0528683, -0.05360271, -0.05364801, -0.05433121, 
    -0.05372288, -0.05346599, -0.0528198, -0.0524414, -0.05208435, 
    -0.05130833, -0.050456, -0.04928926, -0.04846873, -0.0479268, 
    -0.04825836, -0.04796551, -0.04829299, -0.04844731, -0.04676223, 
    -0.04770061, -0.04630008, -0.04637643, -0.04700585, -0.04636782, 
    -0.05300936, -0.05321528, -0.05393665, -0.05337124, -0.05440616, 
    -0.05382423, -0.05349258, -0.05223314, -0.05196073, -0.05170936, 
    -0.05121676, -0.05059177, -0.04951476, -0.04859745, -0.0477758, 
    -0.04783551, -0.04781447, -0.04763275, -0.04808418, -0.04755907, 
    -0.0474715, -0.04770077, -0.04638667, -0.04675814, -0.04637806, 
    -0.04661953, -0.05314826, -0.05280274, -0.05298914, -0.05263917, 
    -0.05288545, -0.0517995, -0.05147852, -0.05000434, -0.05060397, 
    -0.0496533, -0.05050656, -0.05035422, -0.04962245, -0.05046008, 
    -0.04864749, -0.04986856, -0.0476257, -0.0488178, -0.04755202, 
    -0.04777932, -0.04740365, -0.04706981, -0.04665342, -0.04589524, 
    -0.04606965, -0.04544317, -0.05229207, -0.05185194, -0.0518906, 
    -0.05143388, -0.05109882, -0.05038058, -0.04925073, -0.04967244, 
    -0.04890121, -0.04874789, -0.04992079, -0.04919709, -0.05155962, 
    -0.05116987, -0.0514016, -0.05225717, -0.04957483, -0.05093272, 
    -0.04845528, -0.04916863, -0.04711725, -0.0481258, -0.04616595, 
    -0.04535395, -0.04460386, -0.04374361, -0.05161346, -0.05191064, 
    -0.05137987, -0.05065484, -0.04999197, -0.04912479, -0.04903701, 
    -0.04887661, -0.0484638, -0.04811953, -0.04882594, -0.04803364, 
    -0.05107979, -0.04945882, -0.05202339, -0.05123658, -0.0506973, 
    -0.0509332, -0.04972091, -0.04943962, -0.04831377, -0.04889238, 
    -0.04555288, -0.04699952, -0.04310065, -0.04415433, -0.05201487, 
    -0.05161452, -0.05024622, -0.05089242, -0.04906751, -0.04862898, 
    -0.0482756, -0.04782772, -0.04777968, -0.04751668, -0.04794845, 
    -0.04753368, -0.04912296, -0.04840591, -0.05040074, -0.0499073, 
    -0.05013369, -0.05038321, -0.04961729, -0.04881472, -0.04879783, 
    -0.04854348, -0.04783406, -0.04906026, -0.04536945, -0.04761238, 
    -0.05118165, -0.05042623, -0.05031943, -0.05060997, -0.04867275, 
    -0.04936545, -0.04752309, -0.04801374, -0.04721263, -0.04760892, 
    -0.04766752, -0.04818238, -0.04850586, -0.04933343, -0.05001784, 
    -0.05056774, -0.05043931, -0.04983722, -0.0487661, -0.04777528, 
    -0.04799047, -0.04727301, -0.04919747, -0.04838054, -0.04869454, 
    -0.04788031, -0.04968368, -0.04814325, -0.05008569, -0.04991214, 
    -0.0493793, -0.04832558, -0.04809585, -0.04785163, -0.04800219, 
    -0.04873925, -0.04886119, -0.0493922, -0.04953984, -0.04994988, 
    -0.05029202, -0.0499793, -0.04965307, -0.04873898, -0.04793041, 
    -0.04706506, -0.04685586, -0.04587012, -0.04667073, -0.04535725, 
    -0.04647119, -0.04456096, -0.0480557, -0.0465046, -0.04935523, 
    -0.04903945, -0.04847359, -0.04720191, -0.04788411, -0.04708736, 
    -0.04886598, -0.04981653, -0.05006577, -0.0505341, -0.05005512, 
    -0.0500939, -0.04963968, -0.04978518, -0.04870894, -0.04928396, 
    -0.04766896, -0.04709362, -0.04550836, -0.04456457, -0.04362532, 
    -0.04321733, -0.04309396, -0.0430425,
  -0.07888652, -0.07723158, -0.0775505, -0.07623623, -0.07696247, -0.076106, 
    -0.07854813, -0.07716656, -0.07804563, -0.07873614, -0.07375098, 
    -0.07617816, -0.07131527, -0.07280098, -0.06912857, -0.07154429, 
    -0.06865185, -0.06919722, -0.06756967, -0.06803183, -0.06599323, 
    -0.06735747, -0.06496184, -0.06631649, -0.06610259, -0.06740295, 
    -0.07568329, -0.07404868, -0.07578127, -0.07554559, -0.07565129, 
    -0.07694734, -0.07760905, -0.07901463, -0.07875753, -0.07772619, 
    -0.07543988, -0.07620817, -0.07428756, -0.07433038, -0.0722498, 
    -0.0731803, -0.06977365, -0.07072483, -0.06801248, -0.06868424, 
    -0.06804386, -0.06823739, -0.06804134, -0.06902935, -0.06860421, 
    -0.06948034, -0.07300506, -0.07195025, -0.07514382, -0.0771343, 
    -0.07848696, -0.0794616, -0.07932305, -0.0790596, -0.0777202, 
    -0.07648248, -0.07555293, -0.07493766, -0.07433654, -0.07254685, 
    -0.07161812, -0.06958286, -0.0699458, -0.06933221, -0.06875145, 
    -0.06778757, -0.06794526, -0.06752402, -0.06934843, -0.06813025, 
    -0.07015339, -0.06959389, -0.07417341, -0.07600013, -0.07679013, 
    -0.07748907, -0.07921669, -0.07801938, -0.0784891, -0.07737651, 
    -0.07667799, -0.07702267, -0.07492092, -0.07573085, -0.07156347, 
    -0.07332853, -0.06881893, -0.06987116, -0.06856919, -0.06923041, 
    -0.06810144, -0.06911663, -0.06736799, -0.0669933, -0.0672491, 
    -0.06627217, -0.06917335, -0.06804381, -0.07703232, -0.07697599, 
    -0.07671416, -0.07787202, -0.07794347, -0.07902166, -0.07806159, 
    -0.07765638, -0.07663774, -0.07604163, -0.07547947, -0.07425856, 
    -0.07291912, -0.07108821, -0.06980244, -0.0689541, -0.06947305, 
    -0.06901468, -0.06952727, -0.06976891, -0.0671334, -0.06860023, 
    -0.06641176, -0.06653097, -0.06751402, -0.06651752, -0.07693646, 
    -0.07726105, -0.07839886, -0.07750696, -0.07914001, -0.07822149, 
    -0.07769831, -0.07571369, -0.07528488, -0.07488934, -0.07411458, 
    -0.07313237, -0.07144184, -0.07000404, -0.06871784, -0.06881125, 
    -0.06877834, -0.06849407, -0.0692004, -0.06837884, -0.0682419, 
    -0.06860047, -0.06654694, -0.06712701, -0.0665335, -0.06691053, 
    -0.0771554, -0.07661085, -0.07690459, -0.07635316, -0.07674117, 
    -0.07503116, -0.07452621, -0.07220999, -0.07315154, -0.07165914, 
    -0.07299853, -0.07275929, -0.07161076, -0.07292552, -0.07008242, 
    -0.0719969, -0.06848305, -0.07034925, -0.06836782, -0.06872335, 
    -0.0681358, -0.06761396, -0.06696346, -0.06578006, -0.06605216, 
    -0.06507512, -0.07580648, -0.07511368, -0.07517452, -0.074456, 
    -0.07392918, -0.07280067, -0.07102779, -0.07168919, -0.07047994, 
    -0.07023972, -0.07207885, -0.07094371, -0.07465377, -0.07404087, 
    -0.07440524, -0.07575153, -0.07153606, -0.07366809, -0.06978138, 
    -0.07089909, -0.0676881, -0.06926554, -0.06620243, -0.06493605, 
    -0.06376769, -0.06242949, -0.07473847, -0.07520604, -0.07437106, 
    -0.07323145, -0.07219058, -0.07083037, -0.07069276, -0.0704414, 
    -0.06979471, -0.06925572, -0.07036201, -0.06912129, -0.07389925, 
    -0.0713541, -0.07538351, -0.07414576, -0.07329817, -0.07366884, 
    -0.07176521, -0.07132399, -0.06955981, -0.07046612, -0.06524616, 
    -0.06750413, -0.06143053, -0.06306817, -0.0753701, -0.07474012, 
    -0.07258969, -0.07360476, -0.07074057, -0.07005343, -0.06950004, 
    -0.06879908, -0.06872392, -0.06831256, -0.06898798, -0.06833914, 
    -0.0708275, -0.06970408, -0.07283233, -0.07205769, -0.07241302, 
    -0.0728048, -0.07160266, -0.07034442, -0.07031796, -0.0699195, 
    -0.06880899, -0.07072921, -0.06496022, -0.06846222, -0.07405937, 
    -0.07287236, -0.07270464, -0.07316097, -0.070122, -0.07120766, 
    -0.06832257, -0.06909016, -0.06783717, -0.06845681, -0.06854846, 
    -0.06935409, -0.06986059, -0.07115748, -0.07223117, -0.07309463, 
    -0.07289291, -0.07194772, -0.07026824, -0.06871704, -0.06905374, 
    -0.06793156, -0.07094429, -0.06966434, -0.07015613, -0.06888136, 
    -0.07170681, -0.06929285, -0.07233769, -0.07206529, -0.0712294, 
    -0.06957829, -0.06921865, -0.06883649, -0.06907208, -0.07022618, 
    -0.07041723, -0.07124963, -0.07148118, -0.07212451, -0.07266161, 
    -0.07217068, -0.07165879, -0.07022575, -0.06895975, -0.06760654, 
    -0.06727967, -0.06574088, -0.06699049, -0.06494121, -0.0666789, 
    -0.06370091, -0.06915583, -0.06673106, -0.07119166, -0.0706966, 
    -0.06981005, -0.06782043, -0.0688873, -0.06764139, -0.07042474, 
    -0.07191525, -0.07230642, -0.0730418, -0.0722897, -0.07235057, 
    -0.07163779, -0.07186606, -0.07017869, -0.07107989, -0.06855072, 
    -0.06765118, -0.06517676, -0.06370652, -0.06224562, -0.06161173, 
    -0.06142015, -0.06134024,
  -0.08614745, -0.08423818, -0.08460601, -0.08309054, -0.08392785, 
    -0.08294041, -0.08575694, -0.0841632, -0.08517716, -0.0859739, 
    -0.08022729, -0.0830236, -0.07742436, -0.07913367, -0.07491082, 
    -0.07768777, -0.07436323, -0.07498969, -0.07312064, -0.07365122, 
    -0.07131182, -0.07287706, -0.07012921, -0.07168259, -0.07143723, 
    -0.07292926, -0.08245321, -0.08057011, -0.08256613, -0.08229453, 
    -0.08241633, -0.0839104, -0.08467355, -0.08629531, -0.08599859, 
    -0.08480866, -0.08217271, -0.08305819, -0.08084521, -0.08089452, 
    -0.07849939, -0.07957028, -0.07565203, -0.07674539, -0.073629, 
    -0.07440042, -0.07366502, -0.07388725, -0.07366213, -0.07479684, 
    -0.07430851, -0.07531499, -0.07936856, -0.07815475, -0.08183157, 
    -0.084126, -0.08568637, -0.08681123, -0.0866513, -0.08634721, 
    -0.08480175, -0.08337442, -0.08230299, -0.08159406, -0.08090162, 
    -0.07884121, -0.07777269, -0.07543279, -0.07584988, -0.07514479, 
    -0.07447762, -0.07337077, -0.07355182, -0.07306824, -0.07516342, 
    -0.07376422, -0.07608847, -0.07544546, -0.08071374, -0.08281839, 
    -0.08372913, -0.08453515, -0.08652852, -0.08514688, -0.08568884, 
    -0.08440533, -0.08359981, -0.08399726, -0.08157476, -0.08250801, 
    -0.07770982, -0.07974092, -0.07455512, -0.0757641, -0.07426829, 
    -0.07502782, -0.07373113, -0.0748971, -0.07288913, -0.07245912, 
    -0.07275269, -0.07163174, -0.07496227, -0.07366496, -0.0840084, 
    -0.08394343, -0.08364152, -0.08497688, -0.08505931, -0.08630342, 
    -0.08519557, -0.08472814, -0.08355342, -0.08286622, -0.08221833, 
    -0.0808118, -0.07926965, -0.07716323, -0.07568512, -0.07471039, 
    -0.0753066, -0.07477998, -0.07536891, -0.07564659, -0.07261991, 
    -0.07430393, -0.07179189, -0.07192864, -0.07305676, -0.07191321, 
    -0.08389786, -0.08427217, -0.08558471, -0.08455578, -0.08644002, 
    -0.08538005, -0.0847765, -0.08248825, -0.08199411, -0.08153838, 
    -0.08064598, -0.07951511, -0.07756992, -0.07591681, -0.07443902, 
    -0.07454631, -0.07450851, -0.07418202, -0.07499335, -0.07404967, 
    -0.07389243, -0.07430421, -0.07194696, -0.07261257, -0.07193154, 
    -0.07236414, -0.08415033, -0.08352242, -0.08386111, -0.08322532, 
    -0.08367268, -0.08170178, -0.08112007, -0.07845359, -0.07953718, 
    -0.07781987, -0.07936104, -0.07908568, -0.07776422, -0.07927702, 
    -0.0760069, -0.07820842, -0.07416935, -0.07631361, -0.07403702, 
    -0.07444534, -0.07377059, -0.07317148, -0.07242487, -0.07106733, 
    -0.0713794, -0.07025906, -0.0825952, -0.08179685, -0.08186694, 
    -0.08103921, -0.08043247, -0.07913332, -0.07709375, -0.07785442, 
    -0.07646386, -0.07618771, -0.0783027, -0.07699706, -0.08126701, 
    -0.08056109, -0.08098073, -0.08253186, -0.0776783, -0.08013185, 
    -0.07566091, -0.07694576, -0.07325658, -0.07506818, -0.07155176, 
    -0.07009964, -0.06876083, -0.0672285, -0.08136457, -0.08190326, 
    -0.08094137, -0.07962915, -0.07843125, -0.07686674, -0.07670853, 
    -0.07641953, -0.07567624, -0.0750569, -0.07632828, -0.07490247, 
    -0.08039802, -0.07746901, -0.08210775, -0.08068188, -0.07970596, 
    -0.08013272, -0.07794188, -0.07743438, -0.0754063, -0.07644796, 
    -0.07045514, -0.0730454, -0.0660854, -0.06795969, -0.0820923, 
    -0.08136648, -0.0788905, -0.08005892, -0.0767635, -0.07597358, 
    -0.07533762, -0.07453232, -0.07444599, -0.07397356, -0.07474931, 
    -0.07400409, -0.07686344, -0.07557207, -0.07916975, -0.07827836, 
    -0.0786872, -0.07913806, -0.0777549, -0.07630806, -0.07627764, 
    -0.07581966, -0.07454372, -0.07675043, -0.07012735, -0.07414544, 
    -0.08058241, -0.07921582, -0.07902279, -0.07954802, -0.07605239, 
    -0.07730061, -0.07398506, -0.07486669, -0.07342772, -0.07413922, 
    -0.07424447, -0.07516993, -0.07575195, -0.07724288, -0.07847796, 
    -0.07947166, -0.07923948, -0.07815184, -0.0762205, -0.0744381, 
    -0.07482486, -0.07353609, -0.07699774, -0.07552642, -0.07609162, 
    -0.07462684, -0.07787471, -0.07509957, -0.07860051, -0.07828709, 
    -0.07732559, -0.07542753, -0.07501432, -0.0745753, -0.07484592, 
    -0.07617214, -0.07639176, -0.07734887, -0.07761516, -0.07835524, 
    -0.07897326, -0.07840835, -0.07781947, -0.07617165, -0.07471689, 
    -0.07316296, -0.07278777, -0.0710224, -0.0724559, -0.07010557, 
    -0.07209837, -0.06868434, -0.07494214, -0.07215822, -0.07728219, 
    -0.07671294, -0.07569387, -0.07340851, -0.07463366, -0.07320297, 
    -0.07640039, -0.07811449, -0.07856454, -0.07941084, -0.07854529, 
    -0.07861535, -0.07779531, -0.07805789, -0.07611755, -0.07715367, 
    -0.07424707, -0.0732142, -0.07037557, -0.06869076, -0.06701805, 
    -0.0662927, -0.06607352, -0.06598211,
  -0.06724854, -0.06570274, -0.06600055, -0.06477354, -0.06545148, -0.064652, 
    -0.06693238, -0.06564203, -0.06646297, -0.06710804, -0.06245522, 
    -0.06471935, -0.06018564, -0.0615697, -0.05815036, -0.06039893, 
    -0.05770696, -0.05821422, -0.0567008, -0.05713043, -0.05523618, 
    -0.05650358, -0.05427864, -0.0555364, -0.05533773, -0.05654585, 
    -0.06425752, -0.0627328, -0.06434895, -0.06412905, -0.06422766, 
    -0.06543735, -0.06605524, -0.06736824, -0.06712802, -0.06616463, 
    -0.0640304, -0.06474736, -0.06295554, -0.06299547, -0.06105611, 
    -0.06192322, -0.05875054, -0.05963586, -0.05711243, -0.05773707, 
    -0.0571416, -0.05732155, -0.05713926, -0.05805806, -0.05766265, 
    -0.05847763, -0.06175989, -0.06077706, -0.06375419, -0.06561191, 
    -0.06687524, -0.06778593, -0.06765645, -0.06741027, -0.06615902, 
    -0.0650034, -0.06413589, -0.06356188, -0.06300122, -0.0613329, 
    -0.06046769, -0.05857301, -0.05891074, -0.05833981, -0.05779958, 
    -0.05690334, -0.05704994, -0.05665838, -0.0583549, -0.05722193, 
    -0.05910393, -0.05858327, -0.0628491, -0.06455319, -0.06529059, 
    -0.06594318, -0.06755706, -0.06643846, -0.06687724, -0.06583808, 
    -0.06518589, -0.06550768, -0.06354626, -0.06430189, -0.06041678, 
    -0.0620614, -0.05786234, -0.05884128, -0.05763008, -0.05824509, 
    -0.05719513, -0.05813925, -0.05651335, -0.05616517, -0.05640287, 
    -0.05549523, -0.05819201, -0.05714156, -0.0655167, -0.06546409, 
    -0.06521966, -0.06630082, -0.06636755, -0.06737481, -0.06647788, 
    -0.06609943, -0.06514832, -0.06459193, -0.06406734, -0.06292849, 
    -0.0616798, -0.0599742, -0.05877733, -0.05798807, -0.05847083, 
    -0.05804441, -0.05852128, -0.05874613, -0.05629535, -0.05765894, 
    -0.0556249, -0.05573562, -0.05664908, -0.05572313, -0.0654272, 
    -0.06573026, -0.06679294, -0.06595989, -0.06748541, -0.06662723, 
    -0.06613858, -0.0642859, -0.06388579, -0.0635168, -0.06279422, 
    -0.06187855, -0.0603035, -0.05896494, -0.05776833, -0.0578552, 
    -0.0578246, -0.05756022, -0.05821718, -0.05745307, -0.05732574, 
    -0.05765917, -0.05575046, -0.05628941, -0.05573798, -0.05608825, 
    -0.06563161, -0.06512322, -0.06539745, -0.06488267, -0.06524488, 
    -0.0636491, -0.06317811, -0.06101903, -0.06189642, -0.06050589, 
    -0.06175381, -0.06153084, -0.06046084, -0.06168577, -0.05903789, 
    -0.06082051, -0.05754997, -0.05928624, -0.05744282, -0.05777345, 
    -0.05722709, -0.05674197, -0.05613744, -0.05503822, -0.0552909, 
    -0.05438378, -0.06437248, -0.06372607, -0.06378283, -0.06311262, 
    -0.06262136, -0.06156942, -0.05991794, -0.06053387, -0.05940789, 
    -0.05918429, -0.06089685, -0.05983965, -0.06329708, -0.0627255, 
    -0.06306528, -0.0643212, -0.06039126, -0.06237794, -0.05875773, 
    -0.0597981, -0.05681088, -0.05827778, -0.05543046, -0.0542547, 
    -0.0531707, -0.05193007, -0.06337607, -0.06381224, -0.0630334, 
    -0.0619709, -0.06100094, -0.05973412, -0.05960601, -0.059372, 
    -0.05877014, -0.05826864, -0.05929811, -0.05814359, -0.06259346, 
    -0.06022179, -0.06397781, -0.0628233, -0.06203309, -0.06237864, 
    -0.06060469, -0.06019375, -0.05855156, -0.05939502, -0.05454254, 
    -0.05663989, -0.05100461, -0.05252206, -0.0639653, -0.06337761, 
    -0.06137281, -0.06231889, -0.05965052, -0.0590109, -0.05849595, 
    -0.05784388, -0.05777398, -0.05739143, -0.05801958, -0.05741615, 
    -0.05973145, -0.05868579, -0.06159892, -0.06087714, -0.06120819, 
    -0.06157326, -0.06045329, -0.05928174, -0.05925711, -0.05888627, 
    -0.05785311, -0.05963994, -0.05427714, -0.05753061, -0.06274275, 
    -0.06163623, -0.06147993, -0.06190521, -0.05907472, -0.06008543, 
    -0.05740075, -0.05811463, -0.05694946, -0.05752557, -0.0576108, 
    -0.05836016, -0.05883145, -0.06003869, -0.06103876, -0.06184337, 
    -0.06165538, -0.0607747, -0.05921084, -0.05776758, -0.05808076, 
    -0.05703721, -0.05984019, -0.05864882, -0.05910648, -0.05792041, 
    -0.06055029, -0.0583032, -0.06113799, -0.06088421, -0.06010567, 
    -0.05856876, -0.05823416, -0.05787868, -0.05809781, -0.05917168, 
    -0.05934951, -0.06012451, -0.06034014, -0.06093939, -0.06143982, 
    -0.0609824, -0.06050557, -0.05917129, -0.05799333, -0.05673507, 
    -0.05643127, -0.05500184, -0.05616255, -0.0542595, -0.05587307, 
    -0.05310878, -0.05817572, -0.05592152, -0.06007052, -0.05960958, 
    -0.05878441, -0.0569339, -0.05792593, -0.05676747, -0.0593565, 
    -0.06074445, -0.06110886, -0.06179413, -0.06109329, -0.06115, -0.060486, 
    -0.06069862, -0.05912748, -0.05996645, -0.0576129, -0.05677657, 
    -0.05447811, -0.05311397, -0.05175968, -0.05117244, -0.050995, -0.05092099,
  -0.06388779, -0.0621957, -0.06252144, -0.0611801, -0.06192096, -0.06104733, 
    -0.06354145, -0.0621293, -0.06302749, -0.06373385, -0.0586514, 
    -0.06112089, -0.05618334, -0.05768753, -0.05397669, -0.05641495, 
    -0.05349682, -0.05404583, -0.05240908, -0.05287334, -0.0508287, 
    -0.05219606, -0.04979744, -0.05115234, -0.05093816, -0.05224171, 
    -0.0606166, -0.05895376, -0.06071641, -0.06047636, -0.060584, 
    -0.06190551, -0.06258127, -0.06401895, -0.06375575, -0.06270096, 
    -0.0603687, -0.06115149, -0.05919647, -0.05923999, -0.05712903, 
    -0.05807219, -0.05462673, -0.05558663, -0.05285389, -0.0535294, 
    -0.05288542, -0.05307996, -0.05288289, -0.05387678, -0.05344888, 
    -0.05433108, -0.05789445, -0.05682573, -0.06006731, -0.06209637, 
    -0.06347887, -0.06447677, -0.06433482, -0.064065, -0.06269484, 
    -0.06143121, -0.06048382, -0.05985753, -0.05924625, -0.05742997, 
    -0.05648964, -0.0544344, -0.05480034, -0.05418182, -0.05359703, 
    -0.05262791, -0.05278634, -0.05236325, -0.05419815, -0.05297225, 
    -0.05500975, -0.05444551, -0.05908048, -0.06093943, -0.06174508, 
    -0.06245868, -0.06422587, -0.06300065, -0.06348106, -0.06234371, 
    -0.06163064, -0.0619824, -0.05984049, -0.06066504, -0.05643434, 
    -0.05822258, -0.05366495, -0.05472506, -0.05341365, -0.05407925, 
    -0.05294329, -0.05396466, -0.05220662, -0.05183069, -0.05208731, 
    -0.05110795, -0.05402179, -0.05288537, -0.06199226, -0.06193475, 
    -0.06166754, -0.06285001, -0.06292304, -0.06402615, -0.0630438, 
    -0.06262963, -0.06158958, -0.06098172, -0.06040901, -0.05916699, 
    -0.05780731, -0.05595379, -0.05465576, -0.05380101, -0.05432372, 
    -0.053862, -0.05437836, -0.05462195, -0.05197123, -0.05344487, 
    -0.05124778, -0.0513672, -0.05235321, -0.05135374, -0.06189441, 
    -0.06222579, -0.06338874, -0.06247696, -0.06414735, -0.06320731, 
    -0.06267247, -0.06064757, -0.06021089, -0.05980837, -0.05902068, 
    -0.05802357, -0.05631131, -0.05485908, -0.05356321, -0.05365722, 
    -0.0536241, -0.05333808, -0.05404903, -0.05322219, -0.05308449, 
    -0.05344511, -0.05138322, -0.05196481, -0.05136975, -0.05174768, 
    -0.06211791, -0.06156215, -0.06186188, -0.06129931, -0.06169511, 
    -0.05995267, -0.05943906, -0.05708872, -0.05804302, -0.05653113, 
    -0.05788783, -0.05764526, -0.05648219, -0.0578138, -0.05493816, 
    -0.05687295, -0.053327, -0.05520742, -0.0532111, -0.05356875, 
    -0.05297783, -0.05245356, -0.05180076, -0.05061536, -0.05088767, 
    -0.04991059, -0.0607421, -0.06003664, -0.06009855, -0.05936768, 
    -0.05883234, -0.05768722, -0.05589272, -0.05656153, -0.05533935, 
    -0.05509686, -0.05695592, -0.05580776, -0.05956877, -0.0589458, 
    -0.05931608, -0.06068612, -0.05640662, -0.05856723, -0.05463452, 
    -0.05576267, -0.05252801, -0.05411465, -0.05103812, -0.04977168, 
    -0.04860621, -0.04727495, -0.0596549, -0.06013064, -0.05928133, 
    -0.05812408, -0.05706906, -0.05569324, -0.05555425, -0.05530042, 
    -0.05464797, -0.05410476, -0.05522029, -0.05396936, -0.05880197, 
    -0.05622259, -0.0603113, -0.05905237, -0.05819177, -0.05856798, 
    -0.05663845, -0.05619214, -0.05441116, -0.05532538, -0.0500815, 
    -0.05234328, -0.04628376, -0.04790984, -0.06029765, -0.05965658, 
    -0.05747337, -0.05850292, -0.05560254, -0.0549089, -0.05435092, 
    -0.05364497, -0.05356933, -0.05315553, -0.05383512, -0.05318226, 
    -0.05569034, -0.05455658, -0.05771931, -0.05693449, -0.05729436, 
    -0.0576914, -0.05647399, -0.05520254, -0.05517583, -0.05477382, 
    -0.05365496, -0.05559106, -0.04979583, -0.05330605, -0.0589646, 
    -0.0577599, -0.05758987, -0.05805258, -0.05497808, -0.05607454, 
    -0.0531656, -0.053938, -0.05267774, -0.0533006, -0.05339279, -0.05420386, 
    -0.0547144, -0.0560238, -0.05711016, -0.05798528, -0.05778073, 
    -0.05682317, -0.05512566, -0.05356241, -0.05390134, -0.05277258, 
    -0.05580835, -0.05451653, -0.05501251, -0.05372779, -0.05657936, 
    -0.05414217, -0.05721804, -0.05694218, -0.05609651, -0.05442979, 
    -0.05406742, -0.05368262, -0.0539198, -0.0550832, -0.05527603, 
    -0.05611696, -0.0563511, -0.05700215, -0.05754625, -0.0570489, 
    -0.05653077, -0.05508277, -0.0538067, -0.0524461, -0.05211798, 
    -0.05057617, -0.05182787, -0.04977684, -0.05151549, -0.0485397, 
    -0.05400415, -0.05156776, -0.05605835, -0.05555812, -0.05466343, 
    -0.05266093, -0.05373377, -0.0524811, -0.05528361, -0.05679031, 
    -0.05718638, -0.0579317, -0.05716944, -0.0572311, -0.05650952, 
    -0.05674051, -0.05503528, -0.05594538, -0.05339506, -0.05249093, 
    -0.05001213, -0.04854528, -0.04709234, -0.04646338, -0.04627346, 
    -0.04619427,
  -0.04035017, -0.03907184, -0.03931778, -0.03830553, -0.03886447, 
    -0.0382054, -0.04008836, -0.03902173, -0.03969999, -0.0402338, 
    -0.03640078, -0.03826088, -0.03454657, -0.03567605, -0.0328932, 
    -0.03472036, -0.03253425, -0.03294493, -0.03172141, -0.03206819, 
    -0.03054259, -0.03156237, -0.02977479, -0.03078379, -0.03062415, 
    -0.03159644, -0.03788066, -0.03662828, -0.0379559, -0.03777496, 
    -0.03785609, -0.03885281, -0.03936297, -0.04044933, -0.04025035, 
    -0.03945336, -0.03769382, -0.03828395, -0.03681095, -0.03684371, 
    -0.03525646, -0.03596519, -0.0333798, -0.03409905, -0.03205366, 
    -0.03255861, -0.03207722, -0.0322226, -0.03207533, -0.03281844, 
    -0.0324984, -0.03315843, -0.03583157, -0.0350287, -0.03746673, 
    -0.03899687, -0.04004107, -0.04079557, -0.04068821, -0.04048416, 
    -0.03944873, -0.03849493, -0.03778059, -0.03730871, -0.03684842, 
    -0.03548251, -0.03477641, -0.03323578, -0.03350982, -0.03304671, 
    -0.03260919, -0.03188484, -0.03200319, -0.03168719, -0.03305893, 
    -0.03214211, -0.03366669, -0.0332441, -0.03672365, -0.03812404, 
    -0.03873174, -0.03927039, -0.04060581, -0.03967972, -0.04004272, 
    -0.03918359, -0.03864539, -0.03891084, -0.03729587, -0.03791717, 
    -0.03473491, -0.03607827, -0.03265998, -0.03345343, -0.03247205, 
    -0.03296995, -0.03212046, -0.0328842, -0.03157025, -0.03128969, 
    -0.03148119, -0.0307507, -0.03292694, -0.03207718, -0.03891828, 
    -0.03887488, -0.03867324, -0.03956592, -0.0396211, -0.04045478, 
    -0.03971232, -0.03939948, -0.03861441, -0.03815593, -0.0377242, 
    -0.03678877, -0.03576607, -0.03437437, -0.03340153, -0.03276176, 
    -0.03315292, -0.03280739, -0.03319383, -0.03337621, -0.03139455, 
    -0.0324954, -0.03085493, -0.03094397, -0.03167969, -0.03093393, 
    -0.03884443, -0.03909456, -0.03997295, -0.03928419, -0.04054642, 
    -0.03983586, -0.03943183, -0.03790401, -0.03757491, -0.03727167, 
    -0.03667865, -0.03592864, -0.03464259, -0.03355382, -0.03258389, 
    -0.0326542, -0.03262943, -0.03241555, -0.03294734, -0.03232891, 
    -0.03222599, -0.03249558, -0.03095591, -0.03138977, -0.03094587, 
    -0.03122775, -0.03901312, -0.03859372, -0.03881989, -0.03839545, 
    -0.03869404, -0.03738037, -0.03699357, -0.03522618, -0.03594326, 
    -0.03480755, -0.03582659, -0.03564429, -0.03477082, -0.03577095, 
    -0.03361305, -0.03506416, -0.03240726, -0.0338148, -0.03232063, 
    -0.03258804, -0.03214628, -0.03175462, -0.03126735, -0.03038366, 
    -0.03058653, -0.02985898, -0.03797527, -0.03744362, -0.03749027, 
    -0.03693983, -0.03653692, -0.03567581, -0.03432857, -0.03483037, 
    -0.03391368, -0.03373196, -0.03512646, -0.03426485, -0.03709124, 
    -0.0366223, -0.03690099, -0.03793306, -0.03471411, -0.03633747, 
    -0.03338563, -0.03423104, -0.03181022, -0.03299643, -0.03069865, 
    -0.02975563, -0.0288894, -0.02790193, -0.03715609, -0.03751444, 
    -0.03687483, -0.0360042, -0.03521141, -0.03417898, -0.03407476, 
    -0.0338845, -0.0333957, -0.03298903, -0.03382445, -0.03288772, 
    -0.03651407, -0.03457602, -0.03765057, -0.0367025, -0.0360551, 
    -0.03633804, -0.03488811, -0.03455317, -0.03321838, -0.03390321, 
    -0.02998617, -0.03167228, -0.02716813, -0.02837259, -0.03764028, 
    -0.03715736, -0.03551513, -0.0362891, -0.03411097, -0.03359114, 
    -0.03317328, -0.03264504, -0.03258847, -0.03227909, -0.03278728, 
    -0.03229907, -0.03417681, -0.03332726, -0.03569993, -0.03511037, 
    -0.03538064, -0.03567896, -0.03476467, -0.03381114, -0.03379113, 
    -0.03348995, -0.03265251, -0.03410236, -0.0297736, -0.03239161, 
    -0.03663645, -0.03573044, -0.03560267, -0.03595044, -0.03364296, 
    -0.03446495, -0.03228661, -0.03286425, -0.03192206, -0.03238753, 
    -0.03245645, -0.0330632, -0.03344545, -0.03442689, -0.03524229, 
    -0.03589985, -0.03574609, -0.03502678, -0.03375353, -0.03258329, 
    -0.03283682, -0.03199291, -0.03426529, -0.03329727, -0.03366876, 
    -0.03270698, -0.03484375, -0.03301704, -0.03532331, -0.03511614, 
    -0.03448142, -0.03323233, -0.03296109, -0.0326732, -0.03285063, 
    -0.03372172, -0.03386622, -0.03449677, -0.03467244, -0.03516117, 
    -0.03556988, -0.03519628, -0.03480728, -0.0337214, -0.03276602, 
    -0.03174906, -0.03150408, -0.03035447, -0.03128758, -0.02975948, 
    -0.03105455, -0.02884002, -0.03291374, -0.03109353, -0.0344528, 
    -0.03407767, -0.03340728, -0.03190951, -0.03271146, -0.0317752, 
    -0.0338719, -0.0350021, -0.03529953, -0.03585957, -0.03528681, 
    -0.03533312, -0.03479134, -0.03496472, -0.03368582, -0.03436807, 
    -0.03245816, -0.03178253, -0.02993454, -0.02884416, -0.02776664, 
    -0.02730101, -0.02716052, -0.02710195,
  -0.01970495, -0.01870051, -0.01889313, -0.01810233, -0.01853834, 
    -0.01802441, -0.01949858, -0.0186613, -0.01919307, -0.01961318, 
    -0.01662921, -0.01806758, -0.01521542, -0.01607413, -0.01397334, 
    -0.01534703, -0.01370616, -0.01401192, -0.01310461, -0.01336065, 
    -0.01224113, -0.01298748, -0.01168475, -0.01241691, -0.01230052, 
    -0.01301256, -0.01777202, -0.01680408, -0.01783044, -0.01768999, 
    -0.01775294, -0.01852923, -0.01892854, -0.0197832, -0.01962623, 
    -0.01899943, -0.01762706, -0.01808554, -0.01694472, -0.01696996, 
    -0.0157542, -0.01629521, -0.01433697, -0.01487742, -0.01334991, 
    -0.01372426, -0.01336733, -0.01347495, -0.01336593, -0.01391762, 
    -0.01367953, -0.01417134, -0.01619298, -0.015581, -0.01745114, 
    -0.01864185, -0.01946134, -0.02005678, -0.01997189, -0.01981069, 
    -0.0189958, -0.0182499, -0.01769435, -0.01732889, -0.01697359, 
    -0.01592643, -0.01538952, -0.01422918, -0.01443441, -0.01408788, 
    -0.01376187, -0.01322516, -0.01331259, -0.01307939, -0.01409701, 
    -0.01341534, -0.01455213, -0.0142354, -0.01687748, -0.01796112, 
    -0.01843466, -0.01885599, -0.01990677, -0.01917714, -0.01946264, 
    -0.01878799, -0.01836725, -0.01857458, -0.01731896, -0.01780037, 
    -0.01535806, -0.0163818, -0.01379965, -0.01439214, -0.01365996, 
    -0.01403058, -0.01339933, -0.01396663, -0.01299328, -0.01278711, 
    -0.01292777, -0.01239277, -0.0139985, -0.0133673, -0.0185804, 
    -0.01854647, -0.01838898, -0.01908777, -0.01913109, -0.0197875, 
    -0.01920275, -0.01895718, -0.01834308, -0.01798592, -0.01765062, 
    -0.01692763, -0.01614291, -0.01508521, -0.01435325, -0.0138754, 
    -0.01416722, -0.01390938, -0.0141978, -0.01433429, -0.0128641, 
    -0.0136773, -0.01246885, -0.01253391, -0.01307387, -0.01252657, 
    -0.01852268, -0.01871829, -0.01940772, -0.0188668, -0.01985986, 
    -0.01929986, -0.01898255, -0.01779014, -0.01753491, -0.01730026, 
    -0.01684284, -0.01626723, -0.01528811, -0.01446741, -0.01374306, 
    -0.01379535, -0.01377692, -0.01361802, -0.01401371, -0.01355374, 
    -0.01347746, -0.01367744, -0.01254264, -0.01286059, -0.0125353, 
    -0.01274168, -0.01865457, -0.01832693, -0.0185035, -0.01817236, 
    -0.01840522, -0.01738431, -0.01708551, -0.01573116, -0.01627842, 
    -0.01541313, -0.01618917, -0.01604987, -0.01538528, -0.01614663, 
    -0.01451186, -0.01560794, -0.01361187, -0.01466342, -0.0135476, 
    -0.01374614, -0.01341843, -0.01312909, -0.01277073, -0.01212556, 
    -0.01227312, -0.01174552, -0.01784549, -0.01743325, -0.01746936, 
    -0.01704405, -0.01673382, -0.01607395, -0.01505061, -0.01543043, 
    -0.0147378, -0.01460116, -0.0156553, -0.0150025, -0.01716087, 
    -0.01679948, -0.0170141, -0.0178127, -0.01534229, -0.01658059, 
    -0.01434134, -0.01497698, -0.0131701, -0.01405035, -0.01235481, 
    -0.01167093, -0.01104941, -0.0103492, -0.01721095, -0.01748808, 
    -0.01699394, -0.01632508, -0.01571992, -0.0149377, -0.01485912, 
    -0.01471585, -0.01434888, -0.01404482, -0.01467068, -0.01396925, 
    -0.01671625, -0.01523771, -0.01759354, -0.01686119, -0.01636406, 
    -0.01658102, -0.01547424, -0.01522042, -0.01421617, -0.01472993, 
    -0.01183743, -0.0130684, -0.009834953, -0.01068181, -0.01758556, 
    -0.01721193, -0.0159513, -0.01654346, -0.01488641, -0.01449541, 
    -0.01418244, -0.01378853, -0.01374646, -0.0135168, -0.01389441, 
    -0.01353161, -0.01493606, -0.01429764, -0.01609237, -0.01564306, 
    -0.01584878, -0.01607635, -0.01538061, -0.01466068, -0.01464562, 
    -0.01441952, -0.01379409, -0.01487992, -0.01168389, -0.01360025, 
    -0.01681037, -0.01611568, -0.0160181, -0.01628392, -0.01453431, 
    -0.01515368, -0.01352238, -0.01395176, -0.01325265, -0.01359722, 
    -0.01364838, -0.0141002, -0.01438616, -0.0151249, -0.01574342, 
    -0.01624521, -0.01612764, -0.01557954, -0.01461737, -0.01374261, 
    -0.01393131, -0.01330499, -0.01500283, -0.01427519, -0.01455368, 
    -0.01383462, -0.01544059, -0.01406572, -0.01580511, -0.01564746, 
    -0.01516614, -0.0142266, -0.01402398, -0.01380948, -0.01394161, 
    -0.01459346, -0.0147021, -0.01517775, -0.01531073, -0.0156817, 
    -0.01599308, -0.01570841, -0.01541293, -0.01459322, -0.01387857, 
    -0.01312499, -0.0129446, -0.01210436, -0.01278557, -0.0116737, 
    -0.0126148, -0.01101418, -0.01398866, -0.01264334, -0.0151445, 
    -0.01486131, -0.01435756, -0.01324338, -0.01383795, -0.01314426, 
    -0.01470637, -0.01556079, -0.01578699, -0.0162144, -0.01577731, 
    -0.01581258, -0.01540083, -0.0155324, -0.01456649, -0.01508045, 
    -0.01364964, -0.01314967, -0.01180011, -0.01101713, -0.01025399, 
    -0.009927681, -0.009829647, -0.009788836,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  365.2442, 367.1049, 366.7426, 368.2348, 367.4119, 368.3825, 365.6208, 
    367.179, 366.1837, 365.4113, 371.1069, 368.3006, 374.0351, 372.2349, 
    376.7672, 373.7548, 377.3763, 376.6797, 378.7781, 378.1762, 380.8652, 
    379.0562, 382.2616, 380.4327, 380.7185, 378.9965, 368.864, 370.7569, 
    368.7521, 369.0215, 368.9005, 367.4292, 366.6764, 365.1021, 365.3875, 
    366.5439, 369.1428, 368.2665, 370.4768, 370.4268, 372.8975, 371.7822, 
    375.9505, 374.7627, 378.2013, 377.3347, 378.1606, 377.91, 378.1639, 
    376.8934, 377.4374, 376.3206, 371.991, 373.2602, 369.4832, 367.2159, 
    365.6891, 364.6084, 364.7611, 365.0523, 366.5507, 367.9562, 369.0131, 
    369.7211, 370.4196, 372.5399, 373.6645, 376.1911, 375.734, 376.5083, 
    377.2485, 378.4938, 378.2886, 378.8379, 376.4877, 378.0487, 375.4739, 
    376.1771, 370.6107, 368.5027, 367.6084, 366.8123, 364.8785, 366.2133, 
    365.6868, 366.94, 367.7354, 367.3431, 369.7405, 368.8096, 373.7313, 
    371.6062, 377.1622, 375.8278, 377.4824, 376.6375, 378.086, 376.7822, 
    379.0424, 379.5354, 379.1986, 380.4917, 376.71, 378.1607, 367.3321, 
    367.3964, 367.6943, 366.3793, 366.2987, 365.0943, 366.1658, 366.6228, 
    367.781, 368.4555, 369.0973, 370.5107, 372.0937, 374.314, 375.9142, 
    376.9894, 376.3298, 376.9121, 376.2612, 375.9564, 379.351, 377.4426, 
    380.3056, 380.1471, 378.851, 380.1649, 367.4416, 367.0713, 365.7876, 
    366.7919, 364.9633, 365.9863, 366.5754, 368.8293, 369.3207, 369.7771, 
    370.6793, 371.8393, 373.8799, 375.661, 377.2916, 377.1719, 377.2141, 
    377.579, 376.6756, 377.7274, 377.9043, 377.4422, 380.1259, 379.3593, 
    380.1437, 379.6445, 367.1916, 367.8115, 367.4781, 368.1024, 367.6637, 
    369.6132, 370.1987, 372.9457, 371.8165, 373.6144, 371.9988, 372.2848, 
    373.6736, 372.0859, 375.5629, 373.2038, 377.5932, 375.2296, 377.7416, 
    377.2845, 378.0414, 378.7203, 379.5747, 381.1516, 380.786, 382.1069, 
    368.7233, 369.5179, 369.4477, 370.2803, 370.8969, 372.2352, 374.3884, 
    373.5777, 375.0667, 375.3661, 373.1042, 374.4921, 370.0502, 370.7658, 
    370.3395, 368.786, 373.7647, 371.2044, 375.9407, 374.5471, 378.6235, 
    376.593, 380.5849, 382.297, 383.9117, 385.8053, 369.9519, 369.4114, 
    370.3793, 371.7215, 372.9691, 374.6321, 374.8024, 375.1147, 375.9239, 
    376.6053, 375.2136, 376.7762, 370.9323, 373.9874, 369.2074, 370.6429, 
    371.6422, 371.2034, 373.485, 374.0242, 376.2202, 375.0838, 381.8742, 
    378.8641, 387.2502, 384.8956, 369.2227, 369.9499, 372.4882, 371.2791, 
    374.7432, 375.5991, 376.2957, 377.1876, 377.2838, 377.813, 376.9461, 
    377.7786, 374.6357, 376.0381, 372.1973, 373.1299, 372.7006, 372.2302, 
    373.6832, 375.2355, 375.2684, 375.7671, 377.1754, 374.7573, 382.2642, 
    377.6204, 370.7439, 372.1496, 372.3502, 371.8052, 375.5132, 374.167, 
    377.8, 376.8159, 378.4291, 377.627, 377.5091, 376.4805, 375.8411, 
    374.2288, 372.92, 371.8842, 372.1248, 373.2633, 375.3305, 377.2927, 
    376.8624, 378.3064, 374.4913, 376.0882, 375.4706, 377.0823, 373.5562, 
    376.5586, 372.7914, 373.1207, 374.1403, 376.1969, 376.6524, 377.1397, 
    376.8389, 375.3831, 375.1447, 374.1154, 373.8317, 373.0489, 372.4018, 
    372.9931, 373.6148, 375.3835, 376.9822, 378.73, 379.1584, 381.2046, 
    379.5393, 382.2902, 379.9514, 384.0054, 376.7325, 379.882, 374.1866, 
    374.7976, 375.9048, 378.4511, 377.0747, 378.6846, 375.1354, 373.3028, 
    372.8291, 371.9471, 372.8493, 372.7759, 373.6404, 373.3624, 375.4424, 
    374.3242, 377.5062, 378.6718, 381.9684, 383.9973, 386.069, 386.986, 
    387.2654, 387.3822 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.195739e-08, 6.223058e-08, 6.217748e-08, 6.239782e-08, 6.22756e-08, 
    6.241988e-08, 6.201279e-08, 6.224143e-08, 6.209547e-08, 6.198199e-08, 
    6.282544e-08, 6.240766e-08, 6.325951e-08, 6.299303e-08, 6.36625e-08, 
    6.321804e-08, 6.375213e-08, 6.364969e-08, 6.395803e-08, 6.38697e-08, 
    6.426407e-08, 6.39988e-08, 6.446854e-08, 6.420073e-08, 6.424262e-08, 
    6.399005e-08, 6.249174e-08, 6.277342e-08, 6.247505e-08, 6.251522e-08, 
    6.24972e-08, 6.227812e-08, 6.216771e-08, 6.193653e-08, 6.19785e-08, 
    6.21483e-08, 6.253328e-08, 6.240261e-08, 6.273198e-08, 6.272454e-08, 
    6.309124e-08, 6.29259e-08, 6.354229e-08, 6.33671e-08, 6.387339e-08, 
    6.374605e-08, 6.38674e-08, 6.38306e-08, 6.386788e-08, 6.368114e-08, 
    6.376114e-08, 6.359683e-08, 6.295686e-08, 6.314493e-08, 6.258403e-08, 
    6.224678e-08, 6.202281e-08, 6.186388e-08, 6.188635e-08, 6.192918e-08, 
    6.21493e-08, 6.235626e-08, 6.2514e-08, 6.261951e-08, 6.272347e-08, 
    6.303814e-08, 6.320472e-08, 6.357771e-08, 6.351041e-08, 6.362443e-08, 
    6.373339e-08, 6.39163e-08, 6.388619e-08, 6.396677e-08, 6.362144e-08, 
    6.385094e-08, 6.347207e-08, 6.357569e-08, 6.275169e-08, 6.243786e-08, 
    6.230444e-08, 6.218769e-08, 6.190362e-08, 6.209979e-08, 6.202245e-08, 
    6.220644e-08, 6.232334e-08, 6.226553e-08, 6.262239e-08, 6.248365e-08, 
    6.321459e-08, 6.289974e-08, 6.372068e-08, 6.352423e-08, 6.376777e-08, 
    6.36435e-08, 6.385643e-08, 6.366479e-08, 6.399677e-08, 6.406906e-08, 
    6.401966e-08, 6.420943e-08, 6.365416e-08, 6.38674e-08, 6.226391e-08, 
    6.227334e-08, 6.231727e-08, 6.212414e-08, 6.211233e-08, 6.193537e-08, 
    6.209284e-08, 6.215989e-08, 6.233013e-08, 6.243081e-08, 6.252654e-08, 
    6.273701e-08, 6.297206e-08, 6.330077e-08, 6.353696e-08, 6.369527e-08, 
    6.35982e-08, 6.368391e-08, 6.35881e-08, 6.354319e-08, 6.404196e-08, 
    6.376189e-08, 6.418213e-08, 6.415888e-08, 6.396869e-08, 6.41615e-08, 
    6.227996e-08, 6.222569e-08, 6.203729e-08, 6.218473e-08, 6.19161e-08, 
    6.206646e-08, 6.215291e-08, 6.248654e-08, 6.255986e-08, 6.262782e-08, 
    6.276207e-08, 6.293436e-08, 6.323661e-08, 6.349962e-08, 6.373973e-08, 
    6.372213e-08, 6.372833e-08, 6.378196e-08, 6.36491e-08, 6.380377e-08, 
    6.382973e-08, 6.376186e-08, 6.415576e-08, 6.404323e-08, 6.415839e-08, 
    6.408511e-08, 6.224334e-08, 6.233464e-08, 6.22853e-08, 6.237808e-08, 
    6.231271e-08, 6.260337e-08, 6.269052e-08, 6.309833e-08, 6.293097e-08, 
    6.319734e-08, 6.295803e-08, 6.300043e-08, 6.320601e-08, 6.297097e-08, 
    6.348511e-08, 6.313651e-08, 6.378404e-08, 6.343591e-08, 6.380586e-08, 
    6.373869e-08, 6.384992e-08, 6.394953e-08, 6.407485e-08, 6.43061e-08, 
    6.425255e-08, 6.444595e-08, 6.247078e-08, 6.25892e-08, 6.257878e-08, 
    6.270273e-08, 6.27944e-08, 6.29931e-08, 6.331179e-08, 6.319195e-08, 
    6.341197e-08, 6.345614e-08, 6.312188e-08, 6.33271e-08, 6.266848e-08, 
    6.277487e-08, 6.271153e-08, 6.248011e-08, 6.321955e-08, 6.284005e-08, 
    6.354086e-08, 6.333526e-08, 6.393532e-08, 6.363688e-08, 6.422307e-08, 
    6.447366e-08, 6.470955e-08, 6.498519e-08, 6.265385e-08, 6.257338e-08, 
    6.271748e-08, 6.291684e-08, 6.310184e-08, 6.33478e-08, 6.337297e-08, 
    6.341904e-08, 6.35384e-08, 6.363876e-08, 6.34336e-08, 6.366392e-08, 
    6.279953e-08, 6.32525e-08, 6.254295e-08, 6.275658e-08, 6.290509e-08, 
    6.283995e-08, 6.317826e-08, 6.325799e-08, 6.358201e-08, 6.341452e-08, 
    6.44118e-08, 6.397055e-08, 6.51951e-08, 6.485286e-08, 6.254526e-08, 
    6.265358e-08, 6.303058e-08, 6.28512e-08, 6.336422e-08, 6.34905e-08, 
    6.359317e-08, 6.37244e-08, 6.373858e-08, 6.381633e-08, 6.368892e-08, 
    6.38113e-08, 6.334832e-08, 6.355521e-08, 6.298749e-08, 6.312566e-08, 
    6.30621e-08, 6.299238e-08, 6.320757e-08, 6.343683e-08, 6.344175e-08, 
    6.351525e-08, 6.372239e-08, 6.33663e-08, 6.446873e-08, 6.378785e-08, 
    6.27717e-08, 6.298033e-08, 6.301015e-08, 6.292932e-08, 6.347784e-08, 
    6.327909e-08, 6.381444e-08, 6.366975e-08, 6.390682e-08, 6.378902e-08, 
    6.377169e-08, 6.362038e-08, 6.352618e-08, 6.32882e-08, 6.309457e-08, 
    6.294105e-08, 6.297675e-08, 6.314539e-08, 6.345086e-08, 6.373985e-08, 
    6.367654e-08, 6.388881e-08, 6.332702e-08, 6.356257e-08, 6.347153e-08, 
    6.370894e-08, 6.318876e-08, 6.363167e-08, 6.307555e-08, 6.312431e-08, 
    6.327515e-08, 6.357854e-08, 6.364569e-08, 6.371736e-08, 6.367314e-08, 
    6.345861e-08, 6.342348e-08, 6.327148e-08, 6.322951e-08, 6.31137e-08, 
    6.301781e-08, 6.310542e-08, 6.319741e-08, 6.345871e-08, 6.369419e-08, 
    6.395094e-08, 6.401378e-08, 6.431375e-08, 6.406955e-08, 6.447252e-08, 
    6.412989e-08, 6.472303e-08, 6.365737e-08, 6.411983e-08, 6.328201e-08, 
    6.337227e-08, 6.353551e-08, 6.390996e-08, 6.370782e-08, 6.394423e-08, 
    6.34221e-08, 6.315121e-08, 6.308114e-08, 6.295038e-08, 6.308413e-08, 
    6.307325e-08, 6.320123e-08, 6.316011e-08, 6.346739e-08, 6.330233e-08, 
    6.377125e-08, 6.394237e-08, 6.442568e-08, 6.472197e-08, 6.502361e-08, 
    6.515678e-08, 6.519732e-08, 6.521426e-08 ;

 SOM_C_LEACHED =
  4.749521e-20, 2.166047e-20, -1.5443e-20, 3.091888e-20, 5.600154e-20, 
    -7.154138e-20, -4.697594e-20, 4.344937e-20, -6.619853e-20, 2.113425e-20, 
    9.38818e-20, -4.369452e-21, 2.483236e-21, -1.818978e-20, 6.461718e-21, 
    1.843624e-20, -2.207481e-20, 8.66256e-21, -1.517849e-20, -4.697258e-20, 
    4.014227e-20, 8.518192e-20, 4.188453e-20, 2.628613e-22, 8.571384e-21, 
    3.360362e-20, -7.299773e-21, 8.892071e-20, 5.262637e-20, 4.62866e-20, 
    -5.177333e-20, -4.874709e-21, -1.798419e-20, 2.813031e-21, 6.276247e-20, 
    -1.102318e-20, 2.520449e-20, 3.338248e-20, -5.276766e-20, 4.141299e-20, 
    1.456323e-21, 1.092253e-20, -1.617994e-20, 3.946296e-20, -1.02258e-20, 
    4.858414e-20, -1.168864e-21, 6.216324e-20, -2.215445e-20, 3.98493e-20, 
    -1.365568e-20, -3.206656e-20, 2.867888e-21, -5.232617e-20, 7.779421e-22, 
    -1.377497e-20, -1.830971e-20, 7.491389e-20, -7.106918e-21, -2.678266e-20, 
    -1.836653e-20, 3.114689e-21, 1.257022e-20, -4.296603e-21, 1.697582e-20, 
    2.51177e-20, 5.66486e-21, 4.448435e-20, -5.990359e-20, 3.128637e-20, 
    1.084713e-20, 2.311642e-20, 1.662936e-20, 3.05871e-20, -2.139059e-20, 
    -4.322079e-20, 7.975262e-20, 2.432701e-20, -1.064589e-19, 2.220027e-21, 
    1.365183e-20, 2.736295e-20, -9.893185e-21, -2.739144e-21, 6.772856e-20, 
    1.757309e-20, 1.72866e-20, -4.616588e-20, 4.003124e-21, -2.375419e-20, 
    -3.18227e-20, 1.377744e-21, 1.906382e-20, -3.477706e-21, 4.720942e-20, 
    1.32188e-20, -2.637975e-20, -3.41501e-20, 5.887755e-20, 7.143482e-21, 
    3.456792e-20, 1.012433e-20, -1.720789e-20, -7.556175e-20, -4.954169e-21, 
    2.723969e-20, 2.873187e-20, -6.478546e-20, 2.765847e-20, 4.375514e-20, 
    -2.468175e-20, 7.095256e-21, 5.942253e-21, 2.329869e-20, 2.163406e-20, 
    -6.639218e-20, -4.560883e-20, 5.985361e-20, -3.645683e-21, -1.146184e-20, 
    -3.659372e-20, -3.494866e-20, 4.027081e-22, -4.068109e-20, 4.254388e-20, 
    2.537168e-20, 3.218768e-20, 1.340693e-20, 2.038252e-20, -2.406454e-20, 
    -1.435752e-20, -7.625649e-20, 1.011117e-21, -4.344394e-20, -3.281316e-20, 
    6.349894e-20, 8.266335e-20, 5.788183e-20, 2.222867e-20, 5.093267e-20, 
    2.826611e-21, 3.638511e-20, 8.833497e-20, -5.507633e-20, 2.368254e-20, 
    7.943855e-21, 3.891399e-20, -6.73529e-20, -2.440931e-20, 1.014798e-20, 
    6.627557e-20, 3.647341e-20, 4.994532e-21, -3.796176e-20, -3.633893e-20, 
    -1.765576e-20, -4.706144e-20, -2.31947e-20, 1.471938e-20, 4.957314e-20, 
    2.583095e-21, -6.137184e-20, -2.346723e-20, -4.442645e-20, 5.984098e-20, 
    3.992719e-22, 7.897155e-21, 2.848341e-20, 3.215083e-21, -7.725437e-20, 
    2.033385e-20, -6.737003e-20, 2.252252e-20, -4.729812e-20, -4.240905e-20, 
    -7.467941e-21, -4.495631e-21, -2.419117e-20, 2.741784e-20, 2.703258e-20, 
    -3.234001e-21, 6.164624e-20, -4.243234e-20, 1.754577e-20, -4.405648e-20, 
    -2.315886e-20, -4.229161e-20, 2.63885e-20, -2.589862e-20, 4.330895e-20, 
    -1.421545e-20, 3.69084e-20, 4.315891e-20, 1.184168e-20, -2.952744e-20, 
    -4.051298e-20, 2.78821e-21, 5.249932e-20, 5.824536e-20, -3.804131e-20, 
    -1.104184e-20, -3.210862e-20, -3.590039e-21, -2.05256e-21, -3.442081e-20, 
    1.990942e-20, -1.458731e-20, -5.189758e-20, -1.636599e-20, -7.182393e-20, 
    2.41129e-20, 1.403153e-20, 1.617358e-20, 5.461744e-20, -4.276237e-21, 
    2.078382e-20, 1.44138e-20, -2.016748e-20, 2.956324e-21, -5.42251e-21, 
    3.507831e-20, -8.193112e-20, -1.893679e-20, 4.66239e-20, -3.125427e-20, 
    -3.625079e-20, -1.137528e-20, 4.5789e-20, 2.511889e-20, 3.595631e-20, 
    -3.382989e-20, -2.564093e-20, -2.740858e-20, 2.036961e-20, -3.156308e-20, 
    -2.788025e-20, 1.894174e-20, 5.203101e-21, 5.016755e-21, 4.289247e-20, 
    1.756345e-21, 1.870849e-20, 4.136508e-20, 8.098485e-21, -5.322453e-20, 
    6.125905e-20, 7.007521e-20, 3.772211e-21, -4.863619e-20, 2.517972e-20, 
    -1.685283e-20, 1.784034e-20, -6.904053e-20, -2.651895e-20, -2.95515e-20, 
    2.953848e-20, 4.693839e-20, 1.039058e-19, -1.6398e-20, -2.730491e-20, 
    -1.481401e-20, 3.632383e-20, 4.743778e-20, 3.465815e-20, -2.408741e-20, 
    1.105607e-20, 2.685427e-20, -2.964209e-21, -5.937155e-20, 4.885307e-20, 
    -3.860288e-20, -6.149213e-20, 3.5115e-20, 2.777631e-20, -2.979623e-20, 
    -4.85592e-21, -2.519635e-20, 1.478915e-20, -5.791354e-20, -1.109791e-20, 
    -1.735614e-20, -9.124746e-21, 2.963562e-20, 4.702018e-20, 2.304282e-20, 
    -4.730523e-20, -3.074949e-20, -5.819441e-20, -4.385567e-20, 
    -2.507273e-21, -7.692864e-20, 4.220443e-20, -1.067616e-20, 5.513534e-20, 
    -1.14777e-21, 5.42835e-20, 1.054696e-20, 1.837032e-20, -3.292223e-20, 
    -2.992028e-20, -2.337805e-20, 1.786014e-20, -3.91391e-21, 7.471478e-20, 
    -2.058087e-20, -3.993767e-20, -9.789245e-21, -4.581307e-20, 1.043036e-20, 
    -2.497735e-21, 2.289534e-20, 7.405706e-20, -2.578579e-20, -2.286577e-20, 
    -6.533747e-21, 2.161738e-20, 1.401813e-20, -1.003495e-19, -3.65337e-20, 
    -4.810842e-20, 3.919133e-20, 3.299162e-21, 2.733982e-20, 2.580913e-20, 
    -2.431029e-20, -2.034205e-20, 1.126251e-20, 3.476128e-20, 5.686592e-20, 
    -6.038638e-20, 3.089315e-20, 3.186218e-20, 1.777928e-20, -2.683133e-20, 
    -3.342819e-20, -8.856124e-21, -1.586532e-20, -5.742725e-20 ;

 SR =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999958, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 
    0.9999957, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999957, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999957, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999957, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 
    0.9999957, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.3396233, -0.339628, -0.3396271, -0.339631, -0.3396289, -0.3396314, 
    -0.3396243, -0.3396282, -0.3396257, -0.3396237, -0.3396385, -0.3396312, 
    -0.3396466, -0.3396418, -0.3396539, -0.3396458, -0.3396555, -0.3396538, 
    -0.3396594, -0.3396578, -0.3396648, -0.3396602, -0.3396686, -0.3396638, 
    -0.3396645, -0.33966, -0.3396328, -0.3396376, -0.3396325, -0.3396332, 
    -0.3396329, -0.3396289, -0.3396268, -0.339623, -0.3396237, -0.3396266, 
    -0.3396335, -0.3396312, -0.3396372, -0.339637, -0.3396436, -0.3396406, 
    -0.3396518, -0.3396487, -0.3396579, -0.3396555, -0.3396578, -0.3396571, 
    -0.3396578, -0.3396543, -0.3396558, -0.3396528, -0.3396412, -0.3396446, 
    -0.3396344, -0.3396282, -0.3396244, -0.3396217, -0.3396221, -0.3396228, 
    -0.3396266, -0.3396303, -0.3396332, -0.3396351, -0.339637, -0.3396425, 
    -0.3396456, -0.3396524, -0.3396513, -0.3396533, -0.3396553, -0.3396586, 
    -0.3396581, -0.3396595, -0.3396533, -0.3396574, -0.3396506, -0.3396524, 
    -0.3396372, -0.3396318, -0.3396292, -0.3396273, -0.3396224, -0.3396257, 
    -0.3396244, -0.3396277, -0.3396297, -0.3396287, -0.3396352, -0.3396326, 
    -0.3396458, -0.3396401, -0.3396551, -0.3396515, -0.3396559, -0.3396537, 
    -0.3396575, -0.3396541, -0.3396601, -0.3396614, -0.3396605, -0.339664, 
    -0.3396539, -0.3396577, -0.3396287, -0.3396288, -0.3396297, -0.3396262, 
    -0.339626, -0.3396229, -0.3396257, -0.3396268, -0.3396299, -0.3396317, 
    -0.3396334, -0.3396372, -0.3396414, -0.3396474, -0.3396517, -0.3396546, 
    -0.3396529, -0.3396544, -0.3396527, -0.3396519, -0.3396609, -0.3396558, 
    -0.3396635, -0.3396631, -0.3396595, -0.3396631, -0.339629, -0.339628, 
    -0.3396247, -0.3396273, -0.3396226, -0.3396252, -0.3396266, -0.3396326, 
    -0.339634, -0.3396352, -0.3396377, -0.3396408, -0.3396462, -0.339651, 
    -0.3396554, -0.3396551, -0.3396552, -0.3396562, -0.3396538, -0.3396566, 
    -0.339657, -0.3396558, -0.339663, -0.3396609, -0.3396631, -0.3396617, 
    -0.3396283, -0.3396299, -0.3396291, -0.3396307, -0.3396295, -0.3396347, 
    -0.3396363, -0.3396437, -0.3396407, -0.3396455, -0.3396412, -0.339642, 
    -0.3396455, -0.3396415, -0.3396507, -0.3396443, -0.3396562, -0.3396497, 
    -0.3396566, -0.3396554, -0.3396575, -0.3396592, -0.3396615, -0.3396657, 
    -0.3396647, -0.3396683, -0.3396324, -0.3396345, -0.3396344, -0.3396366, 
    -0.3396382, -0.3396419, -0.3396476, -0.3396455, -0.3396495, -0.3396503, 
    -0.3396442, -0.3396479, -0.3396359, -0.3396378, -0.3396367, -0.3396325, 
    -0.3396459, -0.339639, -0.3396518, -0.3396481, -0.339659, -0.3396535, 
    -0.3396642, -0.3396686, -0.3396731, -0.339678, -0.3396357, -0.3396343, 
    -0.3396369, -0.3396404, -0.3396438, -0.3396483, -0.3396488, -0.3396496, 
    -0.3396518, -0.3396536, -0.3396498, -0.3396541, -0.3396381, -0.3396465, 
    -0.3396337, -0.3396375, -0.3396402, -0.3396391, -0.3396452, -0.3396467, 
    -0.3396525, -0.3396495, -0.3396675, -0.3396595, -0.3396819, -0.3396756, 
    -0.3396338, -0.3396357, -0.3396425, -0.3396393, -0.3396486, -0.3396509, 
    -0.3396528, -0.3396551, -0.3396554, -0.3396568, -0.3396545, -0.3396567, 
    -0.3396483, -0.3396521, -0.3396418, -0.3396443, -0.3396431, -0.3396419, 
    -0.3396458, -0.3396498, -0.33965, -0.3396513, -0.3396547, -0.3396486, 
    -0.3396683, -0.339656, -0.3396379, -0.3396415, -0.3396422, -0.3396407, 
    -0.3396506, -0.339647, -0.3396568, -0.3396542, -0.3396585, -0.3396563, 
    -0.339656, -0.3396533, -0.3396515, -0.3396472, -0.3396437, -0.3396409, 
    -0.3396416, -0.3396446, -0.3396501, -0.3396554, -0.3396542, -0.3396581, 
    -0.3396479, -0.3396522, -0.3396505, -0.3396549, -0.3396454, -0.3396531, 
    -0.3396434, -0.3396443, -0.339647, -0.3396524, -0.3396537, -0.339655, 
    -0.3396542, -0.3396502, -0.3396496, -0.3396469, -0.3396461, -0.3396441, 
    -0.3396423, -0.3396439, -0.3396455, -0.3396503, -0.3396546, -0.3396592, 
    -0.3396604, -0.3396657, -0.3396612, -0.3396684, -0.3396621, -0.3396731, 
    -0.3396537, -0.3396621, -0.3396471, -0.3396488, -0.3396516, -0.3396584, 
    -0.3396548, -0.339659, -0.3396496, -0.3396446, -0.3396435, -0.3396411, 
    -0.3396435, -0.3396433, -0.3396457, -0.3396449, -0.3396505, -0.3396475, 
    -0.339656, -0.339659, -0.3396679, -0.3396732, -0.3396789, -0.3396813, 
    -0.339682, -0.3396823 ;

 TAUY =
  -0.3396233, -0.339628, -0.3396271, -0.339631, -0.3396289, -0.3396314, 
    -0.3396243, -0.3396282, -0.3396257, -0.3396237, -0.3396385, -0.3396312, 
    -0.3396466, -0.3396418, -0.3396539, -0.3396458, -0.3396555, -0.3396538, 
    -0.3396594, -0.3396578, -0.3396648, -0.3396602, -0.3396686, -0.3396638, 
    -0.3396645, -0.33966, -0.3396328, -0.3396376, -0.3396325, -0.3396332, 
    -0.3396329, -0.3396289, -0.3396268, -0.339623, -0.3396237, -0.3396266, 
    -0.3396335, -0.3396312, -0.3396372, -0.339637, -0.3396436, -0.3396406, 
    -0.3396518, -0.3396487, -0.3396579, -0.3396555, -0.3396578, -0.3396571, 
    -0.3396578, -0.3396543, -0.3396558, -0.3396528, -0.3396412, -0.3396446, 
    -0.3396344, -0.3396282, -0.3396244, -0.3396217, -0.3396221, -0.3396228, 
    -0.3396266, -0.3396303, -0.3396332, -0.3396351, -0.339637, -0.3396425, 
    -0.3396456, -0.3396524, -0.3396513, -0.3396533, -0.3396553, -0.3396586, 
    -0.3396581, -0.3396595, -0.3396533, -0.3396574, -0.3396506, -0.3396524, 
    -0.3396372, -0.3396318, -0.3396292, -0.3396273, -0.3396224, -0.3396257, 
    -0.3396244, -0.3396277, -0.3396297, -0.3396287, -0.3396352, -0.3396326, 
    -0.3396458, -0.3396401, -0.3396551, -0.3396515, -0.3396559, -0.3396537, 
    -0.3396575, -0.3396541, -0.3396601, -0.3396614, -0.3396605, -0.339664, 
    -0.3396539, -0.3396577, -0.3396287, -0.3396288, -0.3396297, -0.3396262, 
    -0.339626, -0.3396229, -0.3396257, -0.3396268, -0.3396299, -0.3396317, 
    -0.3396334, -0.3396372, -0.3396414, -0.3396474, -0.3396517, -0.3396546, 
    -0.3396529, -0.3396544, -0.3396527, -0.3396519, -0.3396609, -0.3396558, 
    -0.3396635, -0.3396631, -0.3396595, -0.3396631, -0.339629, -0.339628, 
    -0.3396247, -0.3396273, -0.3396226, -0.3396252, -0.3396266, -0.3396326, 
    -0.339634, -0.3396352, -0.3396377, -0.3396408, -0.3396462, -0.339651, 
    -0.3396554, -0.3396551, -0.3396552, -0.3396562, -0.3396538, -0.3396566, 
    -0.339657, -0.3396558, -0.339663, -0.3396609, -0.3396631, -0.3396617, 
    -0.3396283, -0.3396299, -0.3396291, -0.3396307, -0.3396295, -0.3396347, 
    -0.3396363, -0.3396437, -0.3396407, -0.3396455, -0.3396412, -0.339642, 
    -0.3396455, -0.3396415, -0.3396507, -0.3396443, -0.3396562, -0.3396497, 
    -0.3396566, -0.3396554, -0.3396575, -0.3396592, -0.3396615, -0.3396657, 
    -0.3396647, -0.3396683, -0.3396324, -0.3396345, -0.3396344, -0.3396366, 
    -0.3396382, -0.3396419, -0.3396476, -0.3396455, -0.3396495, -0.3396503, 
    -0.3396442, -0.3396479, -0.3396359, -0.3396378, -0.3396367, -0.3396325, 
    -0.3396459, -0.339639, -0.3396518, -0.3396481, -0.339659, -0.3396535, 
    -0.3396642, -0.3396686, -0.3396731, -0.339678, -0.3396357, -0.3396343, 
    -0.3396369, -0.3396404, -0.3396438, -0.3396483, -0.3396488, -0.3396496, 
    -0.3396518, -0.3396536, -0.3396498, -0.3396541, -0.3396381, -0.3396465, 
    -0.3396337, -0.3396375, -0.3396402, -0.3396391, -0.3396452, -0.3396467, 
    -0.3396525, -0.3396495, -0.3396675, -0.3396595, -0.3396819, -0.3396756, 
    -0.3396338, -0.3396357, -0.3396425, -0.3396393, -0.3396486, -0.3396509, 
    -0.3396528, -0.3396551, -0.3396554, -0.3396568, -0.3396545, -0.3396567, 
    -0.3396483, -0.3396521, -0.3396418, -0.3396443, -0.3396431, -0.3396419, 
    -0.3396458, -0.3396498, -0.33965, -0.3396513, -0.3396547, -0.3396486, 
    -0.3396683, -0.339656, -0.3396379, -0.3396415, -0.3396422, -0.3396407, 
    -0.3396506, -0.339647, -0.3396568, -0.3396542, -0.3396585, -0.3396563, 
    -0.339656, -0.3396533, -0.3396515, -0.3396472, -0.3396437, -0.3396409, 
    -0.3396416, -0.3396446, -0.3396501, -0.3396554, -0.3396542, -0.3396581, 
    -0.3396479, -0.3396522, -0.3396505, -0.3396549, -0.3396454, -0.3396531, 
    -0.3396434, -0.3396443, -0.339647, -0.3396524, -0.3396537, -0.339655, 
    -0.3396542, -0.3396502, -0.3396496, -0.3396469, -0.3396461, -0.3396441, 
    -0.3396423, -0.3396439, -0.3396455, -0.3396503, -0.3396546, -0.3396592, 
    -0.3396604, -0.3396657, -0.3396612, -0.3396684, -0.3396621, -0.3396731, 
    -0.3396537, -0.3396621, -0.3396471, -0.3396488, -0.3396516, -0.3396584, 
    -0.3396548, -0.339659, -0.3396496, -0.3396446, -0.3396435, -0.3396411, 
    -0.3396435, -0.3396433, -0.3396457, -0.3396449, -0.3396505, -0.3396475, 
    -0.339656, -0.339659, -0.3396679, -0.3396732, -0.3396789, -0.3396813, 
    -0.339682, -0.3396823 ;

 TBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.8352, 261.8547, 261.8509, 261.8667, 261.8579, 261.8682, 261.8392, 
    261.8555, 261.8451, 261.837, 261.8972, 261.8674, 261.9281, 261.9091, 
    261.9569, 261.9252, 261.9633, 261.956, 261.978, 261.9717, 261.9998, 
    261.9809, 262.0143, 261.9952, 261.9982, 261.9803, 261.8734, 261.8934, 
    261.8722, 261.875, 261.8737, 261.8581, 261.8502, 261.8337, 261.8367, 
    261.8488, 261.8763, 261.867, 261.8905, 261.89, 261.9162, 261.9044, 
    261.9483, 261.9358, 261.9719, 261.9629, 261.9715, 261.9689, 261.9715, 
    261.9582, 261.9639, 261.9522, 261.9066, 261.92, 261.8799, 261.8559, 
    261.8399, 261.8286, 261.8301, 261.8332, 261.8489, 261.8637, 261.875, 
    261.8825, 261.8899, 261.9124, 261.9242, 261.9508, 261.946, 261.9542, 
    261.9619, 261.975, 261.9728, 261.9786, 261.954, 261.9703, 261.9433, 
    261.9507, 261.8919, 261.8695, 261.86, 261.8517, 261.8314, 261.8454, 
    261.8399, 261.853, 261.8614, 261.8572, 261.8827, 261.8728, 261.9249, 
    261.9025, 261.9611, 261.9471, 261.9644, 261.9555, 261.9707, 261.9571, 
    261.9807, 261.9859, 261.9824, 261.9959, 261.9563, 261.9715, 261.8571, 
    261.8578, 261.8609, 261.8471, 261.8463, 261.8336, 261.8449, 261.8497, 
    261.8618, 261.869, 261.8759, 261.8909, 261.9077, 261.9311, 261.9479, 
    261.9592, 261.9523, 261.9584, 261.9516, 261.9484, 261.9839, 261.964, 
    261.9939, 261.9923, 261.9787, 261.9925, 261.8582, 261.8544, 261.8409, 
    261.8515, 261.8323, 261.843, 261.8492, 261.873, 261.8782, 261.8831, 
    261.8927, 261.905, 261.9265, 261.9453, 261.9624, 261.9612, 261.9616, 
    261.9654, 261.9559, 261.967, 261.9688, 261.964, 261.9921, 261.984, 
    261.9922, 261.987, 261.8557, 261.8622, 261.8586, 261.8653, 261.8606, 
    261.8813, 261.8875, 261.9167, 261.9047, 261.9237, 261.9066, 261.9097, 
    261.9243, 261.9076, 261.9442, 261.9194, 261.9656, 261.9407, 261.9671, 
    261.9623, 261.9702, 261.9774, 261.9863, 262.0027, 261.9989, 262.0127, 
    261.8719, 261.8803, 261.8796, 261.8884, 261.895, 261.9091, 261.9319, 
    261.9233, 261.939, 261.9422, 261.9183, 261.933, 261.886, 261.8936, 
    261.8891, 261.8725, 261.9253, 261.8982, 261.9482, 261.9336, 261.9763, 
    261.955, 261.9969, 262.0147, 262.0315, 262.0511, 261.8849, 261.8792, 
    261.8895, 261.9037, 261.9169, 261.9344, 261.9362, 261.9395, 261.9481, 
    261.9552, 261.9406, 261.957, 261.8953, 261.9276, 261.877, 261.8923, 
    261.9029, 261.8982, 261.9224, 261.928, 261.9511, 261.9392, 262.0103, 
    261.9789, 262.066, 262.0417, 261.8772, 261.8849, 261.9118, 261.899, 
    261.9356, 261.9446, 261.952, 261.9613, 261.9623, 261.9679, 261.9588, 
    261.9675, 261.9345, 261.9492, 261.9088, 261.9186, 261.9141, 261.9091, 
    261.9245, 261.9408, 261.9412, 261.9464, 261.9611, 261.9358, 262.0143, 
    261.9658, 261.8934, 261.9082, 261.9104, 261.9046, 261.9437, 261.9296, 
    261.9677, 261.9574, 261.9743, 261.9659, 261.9647, 261.9539, 261.9472, 
    261.9302, 261.9164, 261.9055, 261.908, 261.92, 261.9418, 261.9624, 
    261.9579, 261.973, 261.933, 261.9498, 261.9433, 261.9602, 261.9231, 
    261.9547, 261.915, 261.9185, 261.9293, 261.9509, 261.9557, 261.9608, 
    261.9577, 261.9424, 261.9398, 261.929, 261.926, 261.9178, 261.9109, 
    261.9172, 261.9237, 261.9424, 261.9591, 261.9774, 261.9819, 262.0033, 
    261.9859, 262.0146, 261.9901, 262.0324, 261.9565, 261.9895, 261.9298, 
    261.9362, 261.9478, 261.9745, 261.9601, 261.977, 261.9398, 261.9204, 
    261.9154, 261.9061, 261.9156, 261.9149, 261.924, 261.9211, 261.943, 
    261.9312, 261.9647, 261.9768, 262.0113, 262.0323, 262.0538, 262.0633, 
    262.0662, 262.0674 ;

 TG_R =
  261.8352, 261.8547, 261.8509, 261.8667, 261.8579, 261.8682, 261.8392, 
    261.8555, 261.8451, 261.837, 261.8972, 261.8674, 261.9281, 261.9091, 
    261.9569, 261.9252, 261.9633, 261.956, 261.978, 261.9717, 261.9998, 
    261.9809, 262.0143, 261.9952, 261.9982, 261.9803, 261.8734, 261.8934, 
    261.8722, 261.875, 261.8737, 261.8581, 261.8502, 261.8337, 261.8367, 
    261.8488, 261.8763, 261.867, 261.8905, 261.89, 261.9162, 261.9044, 
    261.9483, 261.9358, 261.9719, 261.9629, 261.9715, 261.9689, 261.9715, 
    261.9582, 261.9639, 261.9522, 261.9066, 261.92, 261.8799, 261.8559, 
    261.8399, 261.8286, 261.8301, 261.8332, 261.8489, 261.8637, 261.875, 
    261.8825, 261.8899, 261.9124, 261.9242, 261.9508, 261.946, 261.9542, 
    261.9619, 261.975, 261.9728, 261.9786, 261.954, 261.9703, 261.9433, 
    261.9507, 261.8919, 261.8695, 261.86, 261.8517, 261.8314, 261.8454, 
    261.8399, 261.853, 261.8614, 261.8572, 261.8827, 261.8728, 261.9249, 
    261.9025, 261.9611, 261.9471, 261.9644, 261.9555, 261.9707, 261.9571, 
    261.9807, 261.9859, 261.9824, 261.9959, 261.9563, 261.9715, 261.8571, 
    261.8578, 261.8609, 261.8471, 261.8463, 261.8336, 261.8449, 261.8497, 
    261.8618, 261.869, 261.8759, 261.8909, 261.9077, 261.9311, 261.9479, 
    261.9592, 261.9523, 261.9584, 261.9516, 261.9484, 261.9839, 261.964, 
    261.9939, 261.9923, 261.9787, 261.9925, 261.8582, 261.8544, 261.8409, 
    261.8515, 261.8323, 261.843, 261.8492, 261.873, 261.8782, 261.8831, 
    261.8927, 261.905, 261.9265, 261.9453, 261.9624, 261.9612, 261.9616, 
    261.9654, 261.9559, 261.967, 261.9688, 261.964, 261.9921, 261.984, 
    261.9922, 261.987, 261.8557, 261.8622, 261.8586, 261.8653, 261.8606, 
    261.8813, 261.8875, 261.9167, 261.9047, 261.9237, 261.9066, 261.9097, 
    261.9243, 261.9076, 261.9442, 261.9194, 261.9656, 261.9407, 261.9671, 
    261.9623, 261.9702, 261.9774, 261.9863, 262.0027, 261.9989, 262.0127, 
    261.8719, 261.8803, 261.8796, 261.8884, 261.895, 261.9091, 261.9319, 
    261.9233, 261.939, 261.9422, 261.9183, 261.933, 261.886, 261.8936, 
    261.8891, 261.8725, 261.9253, 261.8982, 261.9482, 261.9336, 261.9763, 
    261.955, 261.9969, 262.0147, 262.0315, 262.0511, 261.8849, 261.8792, 
    261.8895, 261.9037, 261.9169, 261.9344, 261.9362, 261.9395, 261.9481, 
    261.9552, 261.9406, 261.957, 261.8953, 261.9276, 261.877, 261.8923, 
    261.9029, 261.8982, 261.9224, 261.928, 261.9511, 261.9392, 262.0103, 
    261.9789, 262.066, 262.0417, 261.8772, 261.8849, 261.9118, 261.899, 
    261.9356, 261.9446, 261.952, 261.9613, 261.9623, 261.9679, 261.9588, 
    261.9675, 261.9345, 261.9492, 261.9088, 261.9186, 261.9141, 261.9091, 
    261.9245, 261.9408, 261.9412, 261.9464, 261.9611, 261.9358, 262.0143, 
    261.9658, 261.8934, 261.9082, 261.9104, 261.9046, 261.9437, 261.9296, 
    261.9677, 261.9574, 261.9743, 261.9659, 261.9647, 261.9539, 261.9472, 
    261.9302, 261.9164, 261.9055, 261.908, 261.92, 261.9418, 261.9624, 
    261.9579, 261.973, 261.933, 261.9498, 261.9433, 261.9602, 261.9231, 
    261.9547, 261.915, 261.9185, 261.9293, 261.9509, 261.9557, 261.9608, 
    261.9577, 261.9424, 261.9398, 261.929, 261.926, 261.9178, 261.9109, 
    261.9172, 261.9237, 261.9424, 261.9591, 261.9774, 261.9819, 262.0033, 
    261.9859, 262.0146, 261.9901, 262.0324, 261.9565, 261.9895, 261.9298, 
    261.9362, 261.9478, 261.9745, 261.9601, 261.977, 261.9398, 261.9204, 
    261.9154, 261.9061, 261.9156, 261.9149, 261.924, 261.9211, 261.943, 
    261.9312, 261.9647, 261.9768, 262.0113, 262.0323, 262.0538, 262.0633, 
    262.0662, 262.0674 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  255.214, 255.2139, 255.2139, 255.2138, 255.2139, 255.2138, 255.214, 
    255.2139, 255.2139, 255.214, 255.2136, 255.2138, 255.2134, 255.2135, 
    255.2133, 255.2135, 255.2133, 255.2133, 255.2133, 255.2133, 255.2132, 
    255.2133, 255.2131, 255.2132, 255.2132, 255.2133, 255.2138, 255.2136, 
    255.2138, 255.2137, 255.2137, 255.2138, 255.2139, 255.214, 255.214, 
    255.2139, 255.2137, 255.2138, 255.2137, 255.2137, 255.2135, 255.2136, 
    255.2134, 255.2134, 255.2133, 255.2133, 255.2133, 255.2133, 255.2133, 
    255.2133, 255.2133, 255.2134, 255.2136, 255.2135, 255.2137, 255.2138, 
    255.214, 255.214, 255.214, 255.214, 255.2139, 255.2138, 255.2137, 
    255.2137, 255.2137, 255.2135, 255.2135, 255.2133, 255.2134, 255.2133, 
    255.2133, 255.2133, 255.2133, 255.2133, 255.2134, 255.2133, 255.2134, 
    255.2134, 255.2136, 255.2138, 255.2138, 255.2139, 255.214, 255.2139, 
    255.214, 255.2139, 255.2138, 255.2139, 255.2137, 255.2138, 255.2135, 
    255.2136, 255.2133, 255.2134, 255.2133, 255.2133, 255.2133, 255.2133, 
    255.2133, 255.2132, 255.2132, 255.2132, 255.2133, 255.2133, 255.2139, 
    255.2139, 255.2138, 255.2139, 255.2139, 255.214, 255.2139, 255.2139, 
    255.2138, 255.2138, 255.2137, 255.2137, 255.2135, 255.2134, 255.2134, 
    255.2133, 255.2134, 255.2133, 255.2134, 255.2134, 255.2132, 255.2133, 
    255.2132, 255.2132, 255.2133, 255.2132, 255.2139, 255.2139, 255.214, 
    255.2139, 255.214, 255.2139, 255.2139, 255.2137, 255.2137, 255.2137, 
    255.2137, 255.2136, 255.2135, 255.2134, 255.2133, 255.2133, 255.2133, 
    255.2133, 255.2133, 255.2133, 255.2133, 255.2133, 255.2132, 255.2132, 
    255.2132, 255.2132, 255.2139, 255.2138, 255.2139, 255.2138, 255.2138, 
    255.2137, 255.2137, 255.2135, 255.2136, 255.2135, 255.2136, 255.2135, 
    255.2134, 255.2136, 255.2134, 255.2135, 255.2133, 255.2134, 255.2133, 
    255.2133, 255.2133, 255.2133, 255.2132, 255.2132, 255.2132, 255.2132, 
    255.2138, 255.2137, 255.2137, 255.2137, 255.2136, 255.2136, 255.2134, 
    255.2135, 255.2134, 255.2134, 255.2135, 255.2134, 255.2137, 255.2136, 
    255.2137, 255.2138, 255.2135, 255.2136, 255.2134, 255.2134, 255.2133, 
    255.2133, 255.2132, 255.2131, 255.2131, 255.213, 255.2137, 255.2137, 
    255.2137, 255.2136, 255.2135, 255.2134, 255.2134, 255.2134, 255.2134, 
    255.2133, 255.2134, 255.2133, 255.2136, 255.2135, 255.2137, 255.2136, 
    255.2136, 255.2136, 255.2135, 255.2135, 255.2134, 255.2134, 255.2131, 
    255.2132, 255.213, 255.2131, 255.2137, 255.2137, 255.2135, 255.2136, 
    255.2134, 255.2134, 255.2134, 255.2133, 255.2133, 255.2133, 255.2133, 
    255.2133, 255.2134, 255.2134, 255.2136, 255.2135, 255.2135, 255.2136, 
    255.2135, 255.2134, 255.2134, 255.2134, 255.2133, 255.2134, 255.2131, 
    255.2132, 255.2137, 255.2135, 255.2135, 255.2136, 255.2134, 255.2135, 
    255.2133, 255.2133, 255.2133, 255.2133, 255.2133, 255.2134, 255.2134, 
    255.2135, 255.2135, 255.2136, 255.2136, 255.2135, 255.2134, 255.2133, 
    255.2133, 255.2133, 255.2135, 255.2134, 255.2134, 255.2133, 255.2135, 
    255.2133, 255.2135, 255.2135, 255.2135, 255.2133, 255.2133, 255.2133, 
    255.2133, 255.2134, 255.2134, 255.2135, 255.2135, 255.2135, 255.2136, 
    255.2135, 255.2135, 255.2134, 255.2133, 255.2133, 255.2133, 255.2131, 
    255.2132, 255.2131, 255.2131, 255.213, 255.2133, 255.2132, 255.2135, 
    255.2134, 255.2134, 255.2133, 255.2133, 255.2132, 255.2134, 255.2135, 
    255.2135, 255.2136, 255.2135, 255.2135, 255.2135, 255.2135, 255.2134, 
    255.2135, 255.2133, 255.2133, 255.2132, 255.2131, 255.213, 255.213, 
    255.213, 255.213 ;

 THBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24019, 18.24018, 18.24018, 18.24017, 18.24017, 18.24017, 18.24018, 
    18.24017, 18.24018, 18.24019, 18.24015, 18.24017, 18.24013, 18.24014, 
    18.24011, 18.24013, 18.2401, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24009, 18.24007, 18.24008, 18.24008, 18.24009, 18.24016, 18.24015, 
    18.24016, 18.24016, 18.24016, 18.24017, 18.24018, 18.24019, 18.24019, 
    18.24018, 18.24016, 18.24017, 18.24015, 18.24015, 18.24013, 18.24014, 
    18.24011, 18.24012, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.24011, 18.24014, 18.24013, 18.24016, 18.24017, 18.24018, 
    18.24019, 18.24019, 18.24019, 18.24018, 18.24017, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24013, 18.24011, 18.24011, 18.24011, 18.2401, 
    18.24009, 18.2401, 18.24009, 18.24011, 18.2401, 18.24011, 18.24011, 
    18.24015, 18.24016, 18.24017, 18.24018, 18.24019, 18.24018, 18.24018, 
    18.24018, 18.24017, 18.24017, 18.24016, 18.24016, 18.24013, 18.24014, 
    18.2401, 18.24011, 18.2401, 18.24011, 18.2401, 18.24011, 18.24009, 
    18.24009, 18.24009, 18.24008, 18.24011, 18.2401, 18.24017, 18.24017, 
    18.24017, 18.24018, 18.24018, 18.24019, 18.24018, 18.24018, 18.24017, 
    18.24017, 18.24016, 18.24015, 18.24014, 18.24012, 18.24011, 18.2401, 
    18.24011, 18.2401, 18.24011, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24008, 18.24009, 18.24008, 18.24017, 18.24018, 18.24018, 18.24018, 
    18.24019, 18.24018, 18.24018, 18.24016, 18.24016, 18.24016, 18.24015, 
    18.24014, 18.24013, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.2401, 18.2401, 18.2401, 18.24008, 18.24009, 18.24008, 
    18.24009, 18.24017, 18.24017, 18.24017, 18.24017, 18.24017, 18.24016, 
    18.24015, 18.24013, 18.24014, 18.24013, 18.24014, 18.24014, 18.24013, 
    18.24014, 18.24011, 18.24013, 18.2401, 18.24012, 18.2401, 18.2401, 
    18.2401, 18.24009, 18.24009, 18.24007, 18.24008, 18.24007, 18.24016, 
    18.24016, 18.24016, 18.24015, 18.24015, 18.24014, 18.24012, 18.24013, 
    18.24012, 18.24012, 18.24013, 18.24012, 18.24015, 18.24015, 18.24015, 
    18.24016, 18.24013, 18.24014, 18.24011, 18.24012, 18.24009, 18.24011, 
    18.24008, 18.24007, 18.24006, 18.24004, 18.24015, 18.24016, 18.24015, 
    18.24014, 18.24013, 18.24012, 18.24012, 18.24012, 18.24011, 18.24011, 
    18.24012, 18.24011, 18.24015, 18.24013, 18.24016, 18.24015, 18.24014, 
    18.24014, 18.24013, 18.24013, 18.24011, 18.24012, 18.24007, 18.24009, 
    18.24003, 18.24005, 18.24016, 18.24015, 18.24014, 18.24014, 18.24012, 
    18.24011, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24012, 18.24011, 18.24014, 18.24013, 18.24014, 18.24014, 18.24013, 
    18.24012, 18.24012, 18.24011, 18.2401, 18.24012, 18.24007, 18.2401, 
    18.24015, 18.24014, 18.24014, 18.24014, 18.24011, 18.24012, 18.2401, 
    18.2401, 18.24009, 18.2401, 18.2401, 18.24011, 18.24011, 18.24012, 
    18.24013, 18.24014, 18.24014, 18.24013, 18.24012, 18.2401, 18.2401, 
    18.2401, 18.24012, 18.24011, 18.24011, 18.2401, 18.24013, 18.24011, 
    18.24013, 18.24013, 18.24012, 18.24011, 18.24011, 18.2401, 18.2401, 
    18.24012, 18.24012, 18.24012, 18.24013, 18.24013, 18.24014, 18.24013, 
    18.24013, 18.24012, 18.2401, 18.24009, 18.24009, 18.24007, 18.24009, 
    18.24007, 18.24008, 18.24006, 18.24011, 18.24008, 18.24012, 18.24012, 
    18.24011, 18.24009, 18.2401, 18.24009, 18.24012, 18.24013, 18.24013, 
    18.24014, 18.24013, 18.24013, 18.24013, 18.24013, 18.24012, 18.24012, 
    18.2401, 18.24009, 18.24007, 18.24006, 18.24004, 18.24003, 18.24003, 
    18.24003 ;

 TOTCOLCH4 =
  4.462039e-06, 4.325203e-06, 4.351656e-06, 4.2424e-06, 4.302856e-06, 
    4.231539e-06, 4.434148e-06, 4.319802e-06, 4.392645e-06, 4.449653e-06, 
    4.034039e-06, 4.237558e-06, 3.827714e-06, 3.953823e-06, 3.640763e-06, 
    3.847199e-06, 3.599802e-06, 3.646661e-06, 3.506562e-06, 3.546427e-06, 
    3.370109e-06, 3.488237e-06, 3.280475e-06, 3.398149e-06, 3.379599e-06, 
    3.492165e-06, 4.196245e-06, 4.059115e-06, 4.204432e-06, 4.184731e-06, 
    4.19357e-06, 4.301596e-06, 4.356501e-06, 4.472592e-06, 4.451416e-06, 
    4.366208e-06, 4.175886e-06, 4.240065e-06, 4.079232e-06, 4.082833e-06, 
    3.907129e-06, 3.985898e-06, 3.696084e-06, 3.777397e-06, 3.544759e-06, 
    3.602592e-06, 3.547462e-06, 3.564138e-06, 3.547245e-06, 3.632248e-06, 
    3.595708e-06, 3.67095e-06, 3.971086e-06, 3.881707e-06, 4.1511e-06, 
    4.317118e-06, 4.4291e-06, 4.509345e-06, 4.497961e-06, 4.476291e-06, 
    4.365712e-06, 4.262924e-06, 4.185349e-06, 4.133824e-06, 4.083351e-06, 
    3.932296e-06, 3.85348e-06, 3.679735e-06, 3.710823e-06, 3.658243e-06, 
    3.608371e-06, 3.525364e-06, 3.538964e-06, 3.502619e-06, 3.659637e-06, 
    3.554904e-06, 3.728584e-06, 3.680683e-06, 4.06961e-06, 4.222709e-06, 
    4.288519e-06, 4.346562e-06, 4.489215e-06, 4.390472e-06, 4.429276e-06, 
    4.337232e-06, 4.279199e-06, 4.307859e-06, 4.132419e-06, 4.20022e-06, 
    3.848833e-06, 3.998415e-06, 3.614171e-06, 3.704434e-06, 3.592698e-06, 
    3.649511e-06, 3.552423e-06, 3.639745e-06, 3.489144e-06, 3.456754e-06, 
    3.478871e-06, 3.39431e-06, 3.644614e-06, 3.547456e-06, 4.30866e-06, 
    4.303979e-06, 4.28221e-06, 4.378281e-06, 4.384194e-06, 4.47317e-06, 
    4.393965e-06, 4.360428e-06, 4.275852e-06, 4.226173e-06, 4.179202e-06, 
    4.076791e-06, 3.963815e-06, 3.808378e-06, 3.69855e-06, 3.625787e-06, 
    3.670326e-06, 3.63099e-06, 3.674974e-06, 3.69568e-06, 3.468869e-06, 
    3.595364e-06, 3.40641e-06, 3.416738e-06, 3.501754e-06, 3.415573e-06, 
    4.300694e-06, 4.327653e-06, 4.42183e-06, 4.348049e-06, 4.48291e-06, 
    4.407179e-06, 4.363897e-06, 4.198782e-06, 4.162918e-06, 4.129769e-06, 
    4.064679e-06, 3.981848e-06, 3.838489e-06, 3.715804e-06, 3.605482e-06, 
    3.613512e-06, 3.610684e-06, 3.586234e-06, 3.646935e-06, 3.576316e-06, 
    3.564523e-06, 3.595387e-06, 3.418122e-06, 3.46832e-06, 3.416957e-06, 
    3.449597e-06, 4.318883e-06, 4.273612e-06, 4.298046e-06, 4.252149e-06, 
    4.284455e-06, 4.141656e-06, 4.099282e-06, 3.903747e-06, 3.983467e-06, 
    3.856971e-06, 3.970535e-06, 3.950294e-06, 3.852849e-06, 3.964362e-06, 
    3.722506e-06, 3.885661e-06, 3.585285e-06, 3.745314e-06, 3.575368e-06, 
    3.605956e-06, 3.555387e-06, 3.510384e-06, 3.454176e-06, 3.35161e-06, 
    3.375228e-06, 3.290336e-06, 4.20654e-06, 4.148574e-06, 4.153675e-06, 
    4.093391e-06, 4.049069e-06, 3.9538e-06, 3.803231e-06, 3.859529e-06, 
    3.756492e-06, 3.735963e-06, 3.892628e-06, 3.796062e-06, 4.11e-06, 
    4.058468e-06, 4.089123e-06, 4.201946e-06, 3.846504e-06, 4.027063e-06, 
    3.696745e-06, 3.79226e-06, 3.516781e-06, 3.65252e-06, 3.388262e-06, 
    3.278225e-06, 3.176357e-06, 3.059274e-06, 4.117111e-06, 4.156316e-06, 
    4.086252e-06, 3.990214e-06, 3.902106e-06, 3.786399e-06, 3.774661e-06, 
    3.753197e-06, 3.69789e-06, 3.651684e-06, 3.746411e-06, 3.640146e-06, 
    4.046534e-06, 3.831022e-06, 4.171171e-06, 4.067295e-06, 3.995851e-06, 
    4.027131e-06, 3.865992e-06, 3.828464e-06, 3.677759e-06, 3.75531e-06, 
    3.305207e-06, 3.500896e-06, 2.971638e-06, 3.115202e-06, 4.170052e-06, 
    4.117252e-06, 3.935934e-06, 4.021728e-06, 3.77874e-06, 3.720032e-06, 
    3.67264e-06, 3.612463e-06, 3.606004e-06, 3.570608e-06, 3.628697e-06, 
    3.572899e-06, 3.786154e-06, 3.690125e-06, 3.95648e-06, 3.890829e-06, 
    3.920971e-06, 3.95415e-06, 3.852174e-06, 3.744907e-06, 3.742652e-06, 
    3.70857e-06, 3.613296e-06, 3.777771e-06, 3.280317e-06, 3.583474e-06, 
    4.060034e-06, 3.959858e-06, 3.945671e-06, 3.984267e-06, 3.725897e-06, 
    3.818557e-06, 3.571472e-06, 3.637472e-06, 3.529644e-06, 3.583027e-06, 
    3.590913e-06, 3.660124e-06, 3.703529e-06, 3.814281e-06, 3.905549e-06, 
    3.978661e-06, 3.961605e-06, 3.881492e-06, 3.738398e-06, 3.60541e-06, 
    3.634341e-06, 3.537783e-06, 3.796116e-06, 3.686718e-06, 3.728813e-06, 
    3.619536e-06, 3.861026e-06, 3.654851e-06, 3.914584e-06, 3.891476e-06, 
    3.820408e-06, 3.67934e-06, 3.648503e-06, 3.615678e-06, 3.63592e-06, 
    3.734802e-06, 3.751132e-06, 3.822133e-06, 3.841837e-06, 3.896504e-06, 
    3.942029e-06, 3.900419e-06, 3.856942e-06, 3.734769e-06, 3.626269e-06, 
    3.509742e-06, 3.481515e-06, 3.348199e-06, 3.456504e-06, 3.278662e-06, 
    3.429527e-06, 3.17051e-06, 3.643099e-06, 3.434053e-06, 3.817196e-06, 
    3.774988e-06, 3.699196e-06, 3.528192e-06, 3.620046e-06, 3.512746e-06, 
    3.751775e-06, 3.878732e-06, 3.911933e-06, 3.974194e-06, 3.910515e-06, 
    3.915677e-06, 3.855161e-06, 3.87456e-06, 3.730745e-06, 3.807674e-06, 
    3.591106e-06, 3.513592e-06, 3.299176e-06, 3.171009e-06, 3.043165e-06, 
    2.987551e-06, 2.970728e-06, 2.963709e-06 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24019, 18.24018, 18.24018, 18.24017, 18.24017, 18.24017, 18.24018, 
    18.24017, 18.24018, 18.24019, 18.24015, 18.24017, 18.24013, 18.24014, 
    18.24011, 18.24013, 18.2401, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24009, 18.24007, 18.24008, 18.24008, 18.24009, 18.24016, 18.24015, 
    18.24016, 18.24016, 18.24016, 18.24017, 18.24018, 18.24019, 18.24019, 
    18.24018, 18.24016, 18.24017, 18.24015, 18.24015, 18.24013, 18.24014, 
    18.24011, 18.24012, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.24011, 18.24014, 18.24013, 18.24016, 18.24017, 18.24018, 
    18.24019, 18.24019, 18.24019, 18.24018, 18.24017, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24013, 18.24011, 18.24011, 18.24011, 18.2401, 
    18.24009, 18.2401, 18.24009, 18.24011, 18.2401, 18.24011, 18.24011, 
    18.24015, 18.24016, 18.24017, 18.24018, 18.24019, 18.24018, 18.24018, 
    18.24018, 18.24017, 18.24017, 18.24016, 18.24016, 18.24013, 18.24014, 
    18.2401, 18.24011, 18.2401, 18.24011, 18.2401, 18.24011, 18.24009, 
    18.24009, 18.24009, 18.24008, 18.24011, 18.2401, 18.24017, 18.24017, 
    18.24017, 18.24018, 18.24018, 18.24019, 18.24018, 18.24018, 18.24017, 
    18.24017, 18.24016, 18.24015, 18.24014, 18.24012, 18.24011, 18.2401, 
    18.24011, 18.2401, 18.24011, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24008, 18.24009, 18.24008, 18.24017, 18.24018, 18.24018, 18.24018, 
    18.24019, 18.24018, 18.24018, 18.24016, 18.24016, 18.24016, 18.24015, 
    18.24014, 18.24013, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.2401, 18.2401, 18.2401, 18.24008, 18.24009, 18.24008, 
    18.24009, 18.24017, 18.24017, 18.24017, 18.24017, 18.24017, 18.24016, 
    18.24015, 18.24013, 18.24014, 18.24013, 18.24014, 18.24014, 18.24013, 
    18.24014, 18.24011, 18.24013, 18.2401, 18.24012, 18.2401, 18.2401, 
    18.2401, 18.24009, 18.24009, 18.24007, 18.24008, 18.24007, 18.24016, 
    18.24016, 18.24016, 18.24015, 18.24015, 18.24014, 18.24012, 18.24013, 
    18.24012, 18.24012, 18.24013, 18.24012, 18.24015, 18.24015, 18.24015, 
    18.24016, 18.24013, 18.24014, 18.24011, 18.24012, 18.24009, 18.24011, 
    18.24008, 18.24007, 18.24006, 18.24004, 18.24015, 18.24016, 18.24015, 
    18.24014, 18.24013, 18.24012, 18.24012, 18.24012, 18.24011, 18.24011, 
    18.24012, 18.24011, 18.24015, 18.24013, 18.24016, 18.24015, 18.24014, 
    18.24014, 18.24013, 18.24013, 18.24011, 18.24012, 18.24007, 18.24009, 
    18.24003, 18.24005, 18.24016, 18.24015, 18.24014, 18.24014, 18.24012, 
    18.24011, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24012, 18.24011, 18.24014, 18.24013, 18.24014, 18.24014, 18.24013, 
    18.24012, 18.24012, 18.24011, 18.2401, 18.24012, 18.24007, 18.2401, 
    18.24015, 18.24014, 18.24014, 18.24014, 18.24011, 18.24012, 18.2401, 
    18.2401, 18.24009, 18.2401, 18.2401, 18.24011, 18.24011, 18.24012, 
    18.24013, 18.24014, 18.24014, 18.24013, 18.24012, 18.2401, 18.2401, 
    18.2401, 18.24012, 18.24011, 18.24011, 18.2401, 18.24013, 18.24011, 
    18.24013, 18.24013, 18.24012, 18.24011, 18.24011, 18.2401, 18.2401, 
    18.24012, 18.24012, 18.24012, 18.24013, 18.24013, 18.24014, 18.24013, 
    18.24013, 18.24012, 18.2401, 18.24009, 18.24009, 18.24007, 18.24009, 
    18.24007, 18.24008, 18.24006, 18.24011, 18.24008, 18.24012, 18.24012, 
    18.24011, 18.24009, 18.2401, 18.24009, 18.24012, 18.24013, 18.24013, 
    18.24014, 18.24013, 18.24013, 18.24013, 18.24013, 18.24012, 18.24012, 
    18.2401, 18.24009, 18.24007, 18.24006, 18.24004, 18.24003, 18.24003, 
    18.24003 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976256e-05, 5.976241e-05, 5.976244e-05, 5.976232e-05, 5.976239e-05, 
    5.976231e-05, 5.976253e-05, 5.976241e-05, 5.976249e-05, 5.976254e-05, 
    5.976209e-05, 5.976231e-05, 5.976186e-05, 5.9762e-05, 5.976164e-05, 
    5.976188e-05, 5.976159e-05, 5.976165e-05, 5.976148e-05, 5.976153e-05, 
    5.976132e-05, 5.976146e-05, 5.976121e-05, 5.976135e-05, 5.976133e-05, 
    5.976146e-05, 5.976227e-05, 5.976212e-05, 5.976228e-05, 5.976226e-05, 
    5.976227e-05, 5.976238e-05, 5.976245e-05, 5.976257e-05, 5.976255e-05, 
    5.976246e-05, 5.976225e-05, 5.976232e-05, 5.976214e-05, 5.976214e-05, 
    5.976195e-05, 5.976203e-05, 5.97617e-05, 5.97618e-05, 5.976153e-05, 
    5.976159e-05, 5.976153e-05, 5.976155e-05, 5.976153e-05, 5.976163e-05, 
    5.976159e-05, 5.976167e-05, 5.976202e-05, 5.976192e-05, 5.976222e-05, 
    5.97624e-05, 5.976252e-05, 5.976261e-05, 5.97626e-05, 5.976257e-05, 
    5.976246e-05, 5.976234e-05, 5.976226e-05, 5.97622e-05, 5.976214e-05, 
    5.976198e-05, 5.976189e-05, 5.976169e-05, 5.976172e-05, 5.976166e-05, 
    5.97616e-05, 5.97615e-05, 5.976152e-05, 5.976148e-05, 5.976166e-05, 
    5.976154e-05, 5.976174e-05, 5.976169e-05, 5.976213e-05, 5.97623e-05, 
    5.976237e-05, 5.976243e-05, 5.976259e-05, 5.976248e-05, 5.976252e-05, 
    5.976242e-05, 5.976236e-05, 5.976239e-05, 5.97622e-05, 5.976227e-05, 
    5.976188e-05, 5.976205e-05, 5.976161e-05, 5.976171e-05, 5.976158e-05, 
    5.976165e-05, 5.976154e-05, 5.976164e-05, 5.976146e-05, 5.976142e-05, 
    5.976145e-05, 5.976135e-05, 5.976165e-05, 5.976153e-05, 5.976239e-05, 
    5.976239e-05, 5.976237e-05, 5.976247e-05, 5.976247e-05, 5.976257e-05, 
    5.976249e-05, 5.976245e-05, 5.976236e-05, 5.97623e-05, 5.976225e-05, 
    5.976214e-05, 5.976201e-05, 5.976183e-05, 5.976171e-05, 5.976162e-05, 
    5.976167e-05, 5.976163e-05, 5.976168e-05, 5.97617e-05, 5.976144e-05, 
    5.976159e-05, 5.976136e-05, 5.976137e-05, 5.976147e-05, 5.976137e-05, 
    5.976238e-05, 5.976241e-05, 5.976251e-05, 5.976243e-05, 5.976258e-05, 
    5.97625e-05, 5.976245e-05, 5.976227e-05, 5.976223e-05, 5.97622e-05, 
    5.976213e-05, 5.976203e-05, 5.976187e-05, 5.976173e-05, 5.97616e-05, 
    5.976161e-05, 5.976161e-05, 5.976158e-05, 5.976165e-05, 5.976157e-05, 
    5.976155e-05, 5.976159e-05, 5.976138e-05, 5.976143e-05, 5.976137e-05, 
    5.976141e-05, 5.976241e-05, 5.976235e-05, 5.976238e-05, 5.976233e-05, 
    5.976237e-05, 5.976221e-05, 5.976216e-05, 5.976194e-05, 5.976203e-05, 
    5.976189e-05, 5.976202e-05, 5.976199e-05, 5.976189e-05, 5.976201e-05, 
    5.976174e-05, 5.976192e-05, 5.976158e-05, 5.976176e-05, 5.976156e-05, 
    5.97616e-05, 5.976154e-05, 5.976149e-05, 5.976142e-05, 5.97613e-05, 
    5.976133e-05, 5.976122e-05, 5.976228e-05, 5.976222e-05, 5.976222e-05, 
    5.976215e-05, 5.976211e-05, 5.9762e-05, 5.976183e-05, 5.976189e-05, 
    5.976178e-05, 5.976175e-05, 5.976193e-05, 5.976182e-05, 5.976218e-05, 
    5.976212e-05, 5.976215e-05, 5.976227e-05, 5.976188e-05, 5.976208e-05, 
    5.976171e-05, 5.976182e-05, 5.976149e-05, 5.976165e-05, 5.976134e-05, 
    5.976121e-05, 5.976108e-05, 5.976093e-05, 5.976218e-05, 5.976223e-05, 
    5.976215e-05, 5.976204e-05, 5.976194e-05, 5.976181e-05, 5.976179e-05, 
    5.976177e-05, 5.976171e-05, 5.976165e-05, 5.976176e-05, 5.976164e-05, 
    5.97621e-05, 5.976186e-05, 5.976224e-05, 5.976213e-05, 5.976205e-05, 
    5.976208e-05, 5.97619e-05, 5.976186e-05, 5.976168e-05, 5.976177e-05, 
    5.976124e-05, 5.976147e-05, 5.976082e-05, 5.9761e-05, 5.976224e-05, 
    5.976218e-05, 5.976198e-05, 5.976207e-05, 5.97618e-05, 5.976173e-05, 
    5.976168e-05, 5.976161e-05, 5.97616e-05, 5.976156e-05, 5.976163e-05, 
    5.976156e-05, 5.976181e-05, 5.97617e-05, 5.9762e-05, 5.976193e-05, 
    5.976196e-05, 5.9762e-05, 5.976189e-05, 5.976176e-05, 5.976176e-05, 
    5.976172e-05, 5.976161e-05, 5.97618e-05, 5.976121e-05, 5.976157e-05, 
    5.976212e-05, 5.976201e-05, 5.976199e-05, 5.976203e-05, 5.976174e-05, 
    5.976185e-05, 5.976156e-05, 5.976163e-05, 5.976151e-05, 5.976157e-05, 
    5.976158e-05, 5.976166e-05, 5.976171e-05, 5.976184e-05, 5.976194e-05, 
    5.976203e-05, 5.976201e-05, 5.976192e-05, 5.976175e-05, 5.97616e-05, 
    5.976163e-05, 5.976152e-05, 5.976182e-05, 5.976169e-05, 5.976174e-05, 
    5.976162e-05, 5.97619e-05, 5.976166e-05, 5.976195e-05, 5.976193e-05, 
    5.976185e-05, 5.976169e-05, 5.976165e-05, 5.976161e-05, 5.976163e-05, 
    5.976175e-05, 5.976177e-05, 5.976185e-05, 5.976187e-05, 5.976194e-05, 
    5.976199e-05, 5.976194e-05, 5.976189e-05, 5.976175e-05, 5.976162e-05, 
    5.976149e-05, 5.976145e-05, 5.976129e-05, 5.976142e-05, 5.976121e-05, 
    5.976139e-05, 5.976107e-05, 5.976164e-05, 5.976139e-05, 5.976185e-05, 
    5.976179e-05, 5.976171e-05, 5.976151e-05, 5.976162e-05, 5.976149e-05, 
    5.976177e-05, 5.976191e-05, 5.976195e-05, 5.976202e-05, 5.976195e-05, 
    5.976196e-05, 5.976189e-05, 5.976191e-05, 5.976174e-05, 5.976183e-05, 
    5.976158e-05, 5.976149e-05, 5.976123e-05, 5.976107e-05, 5.976091e-05, 
    5.976084e-05, 5.976082e-05, 5.976081e-05 ;

 TOTLITC_1m =
  5.976256e-05, 5.976241e-05, 5.976244e-05, 5.976232e-05, 5.976239e-05, 
    5.976231e-05, 5.976253e-05, 5.976241e-05, 5.976249e-05, 5.976254e-05, 
    5.976209e-05, 5.976231e-05, 5.976186e-05, 5.9762e-05, 5.976164e-05, 
    5.976188e-05, 5.976159e-05, 5.976165e-05, 5.976148e-05, 5.976153e-05, 
    5.976132e-05, 5.976146e-05, 5.976121e-05, 5.976135e-05, 5.976133e-05, 
    5.976146e-05, 5.976227e-05, 5.976212e-05, 5.976228e-05, 5.976226e-05, 
    5.976227e-05, 5.976238e-05, 5.976245e-05, 5.976257e-05, 5.976255e-05, 
    5.976246e-05, 5.976225e-05, 5.976232e-05, 5.976214e-05, 5.976214e-05, 
    5.976195e-05, 5.976203e-05, 5.97617e-05, 5.97618e-05, 5.976153e-05, 
    5.976159e-05, 5.976153e-05, 5.976155e-05, 5.976153e-05, 5.976163e-05, 
    5.976159e-05, 5.976167e-05, 5.976202e-05, 5.976192e-05, 5.976222e-05, 
    5.97624e-05, 5.976252e-05, 5.976261e-05, 5.97626e-05, 5.976257e-05, 
    5.976246e-05, 5.976234e-05, 5.976226e-05, 5.97622e-05, 5.976214e-05, 
    5.976198e-05, 5.976189e-05, 5.976169e-05, 5.976172e-05, 5.976166e-05, 
    5.97616e-05, 5.97615e-05, 5.976152e-05, 5.976148e-05, 5.976166e-05, 
    5.976154e-05, 5.976174e-05, 5.976169e-05, 5.976213e-05, 5.97623e-05, 
    5.976237e-05, 5.976243e-05, 5.976259e-05, 5.976248e-05, 5.976252e-05, 
    5.976242e-05, 5.976236e-05, 5.976239e-05, 5.97622e-05, 5.976227e-05, 
    5.976188e-05, 5.976205e-05, 5.976161e-05, 5.976171e-05, 5.976158e-05, 
    5.976165e-05, 5.976154e-05, 5.976164e-05, 5.976146e-05, 5.976142e-05, 
    5.976145e-05, 5.976135e-05, 5.976165e-05, 5.976153e-05, 5.976239e-05, 
    5.976239e-05, 5.976237e-05, 5.976247e-05, 5.976247e-05, 5.976257e-05, 
    5.976249e-05, 5.976245e-05, 5.976236e-05, 5.97623e-05, 5.976225e-05, 
    5.976214e-05, 5.976201e-05, 5.976183e-05, 5.976171e-05, 5.976162e-05, 
    5.976167e-05, 5.976163e-05, 5.976168e-05, 5.97617e-05, 5.976144e-05, 
    5.976159e-05, 5.976136e-05, 5.976137e-05, 5.976147e-05, 5.976137e-05, 
    5.976238e-05, 5.976241e-05, 5.976251e-05, 5.976243e-05, 5.976258e-05, 
    5.97625e-05, 5.976245e-05, 5.976227e-05, 5.976223e-05, 5.97622e-05, 
    5.976213e-05, 5.976203e-05, 5.976187e-05, 5.976173e-05, 5.97616e-05, 
    5.976161e-05, 5.976161e-05, 5.976158e-05, 5.976165e-05, 5.976157e-05, 
    5.976155e-05, 5.976159e-05, 5.976138e-05, 5.976143e-05, 5.976137e-05, 
    5.976141e-05, 5.976241e-05, 5.976235e-05, 5.976238e-05, 5.976233e-05, 
    5.976237e-05, 5.976221e-05, 5.976216e-05, 5.976194e-05, 5.976203e-05, 
    5.976189e-05, 5.976202e-05, 5.976199e-05, 5.976189e-05, 5.976201e-05, 
    5.976174e-05, 5.976192e-05, 5.976158e-05, 5.976176e-05, 5.976156e-05, 
    5.97616e-05, 5.976154e-05, 5.976149e-05, 5.976142e-05, 5.97613e-05, 
    5.976133e-05, 5.976122e-05, 5.976228e-05, 5.976222e-05, 5.976222e-05, 
    5.976215e-05, 5.976211e-05, 5.9762e-05, 5.976183e-05, 5.976189e-05, 
    5.976178e-05, 5.976175e-05, 5.976193e-05, 5.976182e-05, 5.976218e-05, 
    5.976212e-05, 5.976215e-05, 5.976227e-05, 5.976188e-05, 5.976208e-05, 
    5.976171e-05, 5.976182e-05, 5.976149e-05, 5.976165e-05, 5.976134e-05, 
    5.976121e-05, 5.976108e-05, 5.976093e-05, 5.976218e-05, 5.976223e-05, 
    5.976215e-05, 5.976204e-05, 5.976194e-05, 5.976181e-05, 5.976179e-05, 
    5.976177e-05, 5.976171e-05, 5.976165e-05, 5.976176e-05, 5.976164e-05, 
    5.97621e-05, 5.976186e-05, 5.976224e-05, 5.976213e-05, 5.976205e-05, 
    5.976208e-05, 5.97619e-05, 5.976186e-05, 5.976168e-05, 5.976177e-05, 
    5.976124e-05, 5.976147e-05, 5.976082e-05, 5.9761e-05, 5.976224e-05, 
    5.976218e-05, 5.976198e-05, 5.976207e-05, 5.97618e-05, 5.976173e-05, 
    5.976168e-05, 5.976161e-05, 5.97616e-05, 5.976156e-05, 5.976163e-05, 
    5.976156e-05, 5.976181e-05, 5.97617e-05, 5.9762e-05, 5.976193e-05, 
    5.976196e-05, 5.9762e-05, 5.976189e-05, 5.976176e-05, 5.976176e-05, 
    5.976172e-05, 5.976161e-05, 5.97618e-05, 5.976121e-05, 5.976157e-05, 
    5.976212e-05, 5.976201e-05, 5.976199e-05, 5.976203e-05, 5.976174e-05, 
    5.976185e-05, 5.976156e-05, 5.976163e-05, 5.976151e-05, 5.976157e-05, 
    5.976158e-05, 5.976166e-05, 5.976171e-05, 5.976184e-05, 5.976194e-05, 
    5.976203e-05, 5.976201e-05, 5.976192e-05, 5.976175e-05, 5.97616e-05, 
    5.976163e-05, 5.976152e-05, 5.976182e-05, 5.976169e-05, 5.976174e-05, 
    5.976162e-05, 5.97619e-05, 5.976166e-05, 5.976195e-05, 5.976193e-05, 
    5.976185e-05, 5.976169e-05, 5.976165e-05, 5.976161e-05, 5.976163e-05, 
    5.976175e-05, 5.976177e-05, 5.976185e-05, 5.976187e-05, 5.976194e-05, 
    5.976199e-05, 5.976194e-05, 5.976189e-05, 5.976175e-05, 5.976162e-05, 
    5.976149e-05, 5.976145e-05, 5.976129e-05, 5.976142e-05, 5.976121e-05, 
    5.976139e-05, 5.976107e-05, 5.976164e-05, 5.976139e-05, 5.976185e-05, 
    5.976179e-05, 5.976171e-05, 5.976151e-05, 5.976162e-05, 5.976149e-05, 
    5.976177e-05, 5.976191e-05, 5.976195e-05, 5.976202e-05, 5.976195e-05, 
    5.976196e-05, 5.976189e-05, 5.976191e-05, 5.976174e-05, 5.976183e-05, 
    5.976158e-05, 5.976149e-05, 5.976123e-05, 5.976107e-05, 5.976091e-05, 
    5.976084e-05, 5.976082e-05, 5.976081e-05 ;

 TOTLITN =
  1.375944e-06, 1.37594e-06, 1.375941e-06, 1.375937e-06, 1.375939e-06, 
    1.375937e-06, 1.375943e-06, 1.37594e-06, 1.375942e-06, 1.375943e-06, 
    1.375931e-06, 1.375937e-06, 1.375924e-06, 1.375928e-06, 1.375918e-06, 
    1.375925e-06, 1.375917e-06, 1.375918e-06, 1.375914e-06, 1.375915e-06, 
    1.375909e-06, 1.375913e-06, 1.375906e-06, 1.37591e-06, 1.375909e-06, 
    1.375913e-06, 1.375936e-06, 1.375931e-06, 1.375936e-06, 1.375935e-06, 
    1.375936e-06, 1.375939e-06, 1.375941e-06, 1.375944e-06, 1.375944e-06, 
    1.375941e-06, 1.375935e-06, 1.375937e-06, 1.375932e-06, 1.375932e-06, 
    1.375927e-06, 1.375929e-06, 1.37592e-06, 1.375922e-06, 1.375915e-06, 
    1.375917e-06, 1.375915e-06, 1.375916e-06, 1.375915e-06, 1.375918e-06, 
    1.375917e-06, 1.375919e-06, 1.375929e-06, 1.375926e-06, 1.375934e-06, 
    1.37594e-06, 1.375943e-06, 1.375945e-06, 1.375945e-06, 1.375944e-06, 
    1.375941e-06, 1.375938e-06, 1.375935e-06, 1.375934e-06, 1.375932e-06, 
    1.375927e-06, 1.375925e-06, 1.375919e-06, 1.37592e-06, 1.375919e-06, 
    1.375917e-06, 1.375914e-06, 1.375915e-06, 1.375913e-06, 1.375919e-06, 
    1.375915e-06, 1.375921e-06, 1.375919e-06, 1.375932e-06, 1.375937e-06, 
    1.375939e-06, 1.37594e-06, 1.375945e-06, 1.375942e-06, 1.375943e-06, 
    1.37594e-06, 1.375938e-06, 1.375939e-06, 1.375934e-06, 1.375936e-06, 
    1.375925e-06, 1.37593e-06, 1.375917e-06, 1.37592e-06, 1.375916e-06, 
    1.375918e-06, 1.375915e-06, 1.375918e-06, 1.375913e-06, 1.375912e-06, 
    1.375913e-06, 1.37591e-06, 1.375918e-06, 1.375915e-06, 1.375939e-06, 
    1.375939e-06, 1.375938e-06, 1.375941e-06, 1.375942e-06, 1.375944e-06, 
    1.375942e-06, 1.375941e-06, 1.375938e-06, 1.375937e-06, 1.375935e-06, 
    1.375932e-06, 1.375928e-06, 1.375923e-06, 1.37592e-06, 1.375918e-06, 
    1.375919e-06, 1.375918e-06, 1.375919e-06, 1.37592e-06, 1.375912e-06, 
    1.375917e-06, 1.37591e-06, 1.375911e-06, 1.375913e-06, 1.375911e-06, 
    1.375939e-06, 1.37594e-06, 1.375943e-06, 1.37594e-06, 1.375945e-06, 
    1.375942e-06, 1.375941e-06, 1.375936e-06, 1.375935e-06, 1.375934e-06, 
    1.375932e-06, 1.375929e-06, 1.375925e-06, 1.375921e-06, 1.375917e-06, 
    1.375917e-06, 1.375917e-06, 1.375916e-06, 1.375918e-06, 1.375916e-06, 
    1.375916e-06, 1.375917e-06, 1.375911e-06, 1.375912e-06, 1.375911e-06, 
    1.375912e-06, 1.37594e-06, 1.375938e-06, 1.375939e-06, 1.375937e-06, 
    1.375938e-06, 1.375934e-06, 1.375933e-06, 1.375927e-06, 1.375929e-06, 
    1.375925e-06, 1.375929e-06, 1.375928e-06, 1.375925e-06, 1.375928e-06, 
    1.375921e-06, 1.375926e-06, 1.375916e-06, 1.375921e-06, 1.375916e-06, 
    1.375917e-06, 1.375915e-06, 1.375914e-06, 1.375912e-06, 1.375908e-06, 
    1.375909e-06, 1.375906e-06, 1.375936e-06, 1.375934e-06, 1.375934e-06, 
    1.375933e-06, 1.375931e-06, 1.375928e-06, 1.375923e-06, 1.375925e-06, 
    1.375922e-06, 1.375921e-06, 1.375926e-06, 1.375923e-06, 1.375933e-06, 
    1.375931e-06, 1.375932e-06, 1.375936e-06, 1.375925e-06, 1.375931e-06, 
    1.37592e-06, 1.375923e-06, 1.375914e-06, 1.375918e-06, 1.37591e-06, 
    1.375906e-06, 1.375902e-06, 1.375898e-06, 1.375933e-06, 1.375935e-06, 
    1.375932e-06, 1.375929e-06, 1.375927e-06, 1.375923e-06, 1.375922e-06, 
    1.375922e-06, 1.37592e-06, 1.375918e-06, 1.375921e-06, 1.375918e-06, 
    1.375931e-06, 1.375924e-06, 1.375935e-06, 1.375932e-06, 1.37593e-06, 
    1.375931e-06, 1.375925e-06, 1.375924e-06, 1.375919e-06, 1.375922e-06, 
    1.375907e-06, 1.375913e-06, 1.375895e-06, 1.3759e-06, 1.375935e-06, 
    1.375933e-06, 1.375928e-06, 1.37593e-06, 1.375923e-06, 1.375921e-06, 
    1.375919e-06, 1.375917e-06, 1.375917e-06, 1.375916e-06, 1.375918e-06, 
    1.375916e-06, 1.375923e-06, 1.37592e-06, 1.375928e-06, 1.375926e-06, 
    1.375927e-06, 1.375928e-06, 1.375925e-06, 1.375921e-06, 1.375921e-06, 
    1.37592e-06, 1.375917e-06, 1.375922e-06, 1.375906e-06, 1.375916e-06, 
    1.375932e-06, 1.375928e-06, 1.375928e-06, 1.375929e-06, 1.375921e-06, 
    1.375924e-06, 1.375916e-06, 1.375918e-06, 1.375914e-06, 1.375916e-06, 
    1.375916e-06, 1.375919e-06, 1.37592e-06, 1.375924e-06, 1.375927e-06, 
    1.375929e-06, 1.375928e-06, 1.375926e-06, 1.375921e-06, 1.375917e-06, 
    1.375918e-06, 1.375915e-06, 1.375923e-06, 1.37592e-06, 1.375921e-06, 
    1.375917e-06, 1.375925e-06, 1.375918e-06, 1.375927e-06, 1.375926e-06, 
    1.375924e-06, 1.375919e-06, 1.375918e-06, 1.375917e-06, 1.375918e-06, 
    1.375921e-06, 1.375922e-06, 1.375924e-06, 1.375925e-06, 1.375926e-06, 
    1.375928e-06, 1.375926e-06, 1.375925e-06, 1.375921e-06, 1.375918e-06, 
    1.375914e-06, 1.375913e-06, 1.375908e-06, 1.375912e-06, 1.375906e-06, 
    1.375911e-06, 1.375902e-06, 1.375918e-06, 1.375911e-06, 1.375924e-06, 
    1.375922e-06, 1.37592e-06, 1.375914e-06, 1.375917e-06, 1.375914e-06, 
    1.375922e-06, 1.375926e-06, 1.375927e-06, 1.375929e-06, 1.375927e-06, 
    1.375927e-06, 1.375925e-06, 1.375926e-06, 1.375921e-06, 1.375923e-06, 
    1.375916e-06, 1.375914e-06, 1.375907e-06, 1.375902e-06, 1.375898e-06, 
    1.375896e-06, 1.375895e-06, 1.375895e-06 ;

 TOTLITN_1m =
  1.375944e-06, 1.37594e-06, 1.375941e-06, 1.375937e-06, 1.375939e-06, 
    1.375937e-06, 1.375943e-06, 1.37594e-06, 1.375942e-06, 1.375943e-06, 
    1.375931e-06, 1.375937e-06, 1.375924e-06, 1.375928e-06, 1.375918e-06, 
    1.375925e-06, 1.375917e-06, 1.375918e-06, 1.375914e-06, 1.375915e-06, 
    1.375909e-06, 1.375913e-06, 1.375906e-06, 1.37591e-06, 1.375909e-06, 
    1.375913e-06, 1.375936e-06, 1.375931e-06, 1.375936e-06, 1.375935e-06, 
    1.375936e-06, 1.375939e-06, 1.375941e-06, 1.375944e-06, 1.375944e-06, 
    1.375941e-06, 1.375935e-06, 1.375937e-06, 1.375932e-06, 1.375932e-06, 
    1.375927e-06, 1.375929e-06, 1.37592e-06, 1.375922e-06, 1.375915e-06, 
    1.375917e-06, 1.375915e-06, 1.375916e-06, 1.375915e-06, 1.375918e-06, 
    1.375917e-06, 1.375919e-06, 1.375929e-06, 1.375926e-06, 1.375934e-06, 
    1.37594e-06, 1.375943e-06, 1.375945e-06, 1.375945e-06, 1.375944e-06, 
    1.375941e-06, 1.375938e-06, 1.375935e-06, 1.375934e-06, 1.375932e-06, 
    1.375927e-06, 1.375925e-06, 1.375919e-06, 1.37592e-06, 1.375919e-06, 
    1.375917e-06, 1.375914e-06, 1.375915e-06, 1.375913e-06, 1.375919e-06, 
    1.375915e-06, 1.375921e-06, 1.375919e-06, 1.375932e-06, 1.375937e-06, 
    1.375939e-06, 1.37594e-06, 1.375945e-06, 1.375942e-06, 1.375943e-06, 
    1.37594e-06, 1.375938e-06, 1.375939e-06, 1.375934e-06, 1.375936e-06, 
    1.375925e-06, 1.37593e-06, 1.375917e-06, 1.37592e-06, 1.375916e-06, 
    1.375918e-06, 1.375915e-06, 1.375918e-06, 1.375913e-06, 1.375912e-06, 
    1.375913e-06, 1.37591e-06, 1.375918e-06, 1.375915e-06, 1.375939e-06, 
    1.375939e-06, 1.375938e-06, 1.375941e-06, 1.375942e-06, 1.375944e-06, 
    1.375942e-06, 1.375941e-06, 1.375938e-06, 1.375937e-06, 1.375935e-06, 
    1.375932e-06, 1.375928e-06, 1.375923e-06, 1.37592e-06, 1.375918e-06, 
    1.375919e-06, 1.375918e-06, 1.375919e-06, 1.37592e-06, 1.375912e-06, 
    1.375917e-06, 1.37591e-06, 1.375911e-06, 1.375913e-06, 1.375911e-06, 
    1.375939e-06, 1.37594e-06, 1.375943e-06, 1.37594e-06, 1.375945e-06, 
    1.375942e-06, 1.375941e-06, 1.375936e-06, 1.375935e-06, 1.375934e-06, 
    1.375932e-06, 1.375929e-06, 1.375925e-06, 1.375921e-06, 1.375917e-06, 
    1.375917e-06, 1.375917e-06, 1.375916e-06, 1.375918e-06, 1.375916e-06, 
    1.375916e-06, 1.375917e-06, 1.375911e-06, 1.375912e-06, 1.375911e-06, 
    1.375912e-06, 1.37594e-06, 1.375938e-06, 1.375939e-06, 1.375937e-06, 
    1.375938e-06, 1.375934e-06, 1.375933e-06, 1.375927e-06, 1.375929e-06, 
    1.375925e-06, 1.375929e-06, 1.375928e-06, 1.375925e-06, 1.375928e-06, 
    1.375921e-06, 1.375926e-06, 1.375916e-06, 1.375921e-06, 1.375916e-06, 
    1.375917e-06, 1.375915e-06, 1.375914e-06, 1.375912e-06, 1.375908e-06, 
    1.375909e-06, 1.375906e-06, 1.375936e-06, 1.375934e-06, 1.375934e-06, 
    1.375933e-06, 1.375931e-06, 1.375928e-06, 1.375923e-06, 1.375925e-06, 
    1.375922e-06, 1.375921e-06, 1.375926e-06, 1.375923e-06, 1.375933e-06, 
    1.375931e-06, 1.375932e-06, 1.375936e-06, 1.375925e-06, 1.375931e-06, 
    1.37592e-06, 1.375923e-06, 1.375914e-06, 1.375918e-06, 1.37591e-06, 
    1.375906e-06, 1.375902e-06, 1.375898e-06, 1.375933e-06, 1.375935e-06, 
    1.375932e-06, 1.375929e-06, 1.375927e-06, 1.375923e-06, 1.375922e-06, 
    1.375922e-06, 1.37592e-06, 1.375918e-06, 1.375921e-06, 1.375918e-06, 
    1.375931e-06, 1.375924e-06, 1.375935e-06, 1.375932e-06, 1.37593e-06, 
    1.375931e-06, 1.375925e-06, 1.375924e-06, 1.375919e-06, 1.375922e-06, 
    1.375907e-06, 1.375913e-06, 1.375895e-06, 1.3759e-06, 1.375935e-06, 
    1.375933e-06, 1.375928e-06, 1.37593e-06, 1.375923e-06, 1.375921e-06, 
    1.375919e-06, 1.375917e-06, 1.375917e-06, 1.375916e-06, 1.375918e-06, 
    1.375916e-06, 1.375923e-06, 1.37592e-06, 1.375928e-06, 1.375926e-06, 
    1.375927e-06, 1.375928e-06, 1.375925e-06, 1.375921e-06, 1.375921e-06, 
    1.37592e-06, 1.375917e-06, 1.375922e-06, 1.375906e-06, 1.375916e-06, 
    1.375932e-06, 1.375928e-06, 1.375928e-06, 1.375929e-06, 1.375921e-06, 
    1.375924e-06, 1.375916e-06, 1.375918e-06, 1.375914e-06, 1.375916e-06, 
    1.375916e-06, 1.375919e-06, 1.37592e-06, 1.375924e-06, 1.375927e-06, 
    1.375929e-06, 1.375928e-06, 1.375926e-06, 1.375921e-06, 1.375917e-06, 
    1.375918e-06, 1.375915e-06, 1.375923e-06, 1.37592e-06, 1.375921e-06, 
    1.375917e-06, 1.375925e-06, 1.375918e-06, 1.375927e-06, 1.375926e-06, 
    1.375924e-06, 1.375919e-06, 1.375918e-06, 1.375917e-06, 1.375918e-06, 
    1.375921e-06, 1.375922e-06, 1.375924e-06, 1.375925e-06, 1.375926e-06, 
    1.375928e-06, 1.375926e-06, 1.375925e-06, 1.375921e-06, 1.375918e-06, 
    1.375914e-06, 1.375913e-06, 1.375908e-06, 1.375912e-06, 1.375906e-06, 
    1.375911e-06, 1.375902e-06, 1.375918e-06, 1.375911e-06, 1.375924e-06, 
    1.375922e-06, 1.37592e-06, 1.375914e-06, 1.375917e-06, 1.375914e-06, 
    1.375922e-06, 1.375926e-06, 1.375927e-06, 1.375929e-06, 1.375927e-06, 
    1.375927e-06, 1.375925e-06, 1.375926e-06, 1.375921e-06, 1.375923e-06, 
    1.375916e-06, 1.375914e-06, 1.375907e-06, 1.375902e-06, 1.375898e-06, 
    1.375896e-06, 1.375895e-06, 1.375895e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34481, 17.34479, 17.3448, 17.34479, 17.34479, 17.34479, 17.3448, 
    17.34479, 17.3448, 17.34481, 17.34476, 17.34479, 17.34474, 17.34476, 
    17.34472, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34475, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.34479, 
    17.3448, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34471, 17.34472, 17.34471, 17.34473, 17.34472, 17.34473, 
    17.34473, 17.34477, 17.34478, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.3448, 17.3448, 17.34479, 17.34479, 17.34477, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34472, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.34479, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34478, 17.34478, 17.34477, 17.34476, 17.34474, 17.34473, 
    17.34472, 17.34473, 17.34472, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.34479, 17.3448, 
    17.3448, 17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34477, 
    17.34477, 17.34476, 17.34475, 17.34473, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 
    17.3447, 17.34471, 17.34479, 17.34479, 17.34479, 17.34479, 17.34479, 
    17.34478, 17.34477, 17.34475, 17.34476, 17.34475, 17.34476, 17.34476, 
    17.34475, 17.34476, 17.34473, 17.34475, 17.34472, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34471, 17.34471, 17.34469, 17.3447, 17.34469, 
    17.34478, 17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 
    17.34475, 17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 
    17.34477, 17.34478, 17.34475, 17.34476, 17.34473, 17.34474, 17.34471, 
    17.34473, 17.3447, 17.34469, 17.34468, 17.34466, 17.34477, 17.34478, 
    17.34477, 17.34476, 17.34475, 17.34474, 17.34474, 17.34474, 17.34473, 
    17.34473, 17.34474, 17.34472, 17.34477, 17.34475, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 
    17.34471, 17.34465, 17.34467, 17.34478, 17.34477, 17.34476, 17.34476, 
    17.34474, 17.34473, 17.34473, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34474, 17.34473, 17.34476, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 
    17.34472, 17.34477, 17.34476, 17.34476, 17.34476, 17.34473, 17.34474, 
    17.34472, 17.34472, 17.34471, 17.34472, 17.34472, 17.34473, 17.34473, 
    17.34474, 17.34475, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34474, 17.34473, 17.34473, 17.34472, 17.34475, 
    17.34473, 17.34475, 17.34475, 17.34474, 17.34473, 17.34473, 17.34472, 
    17.34472, 17.34473, 17.34474, 17.34474, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34475, 17.34473, 17.34472, 17.34471, 17.34471, 17.34469, 
    17.34471, 17.34469, 17.3447, 17.34468, 17.34472, 17.3447, 17.34474, 
    17.34474, 17.34473, 17.34471, 17.34472, 17.34471, 17.34474, 17.34475, 
    17.34475, 17.34476, 17.34475, 17.34475, 17.34475, 17.34475, 17.34473, 
    17.34474, 17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34465, 
    17.34465, 17.34465 ;

 TOTSOMC_1m =
  17.34481, 17.34479, 17.3448, 17.34479, 17.34479, 17.34479, 17.3448, 
    17.34479, 17.3448, 17.34481, 17.34476, 17.34479, 17.34474, 17.34476, 
    17.34472, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34475, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.34479, 
    17.3448, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34471, 17.34472, 17.34471, 17.34473, 17.34472, 17.34473, 
    17.34473, 17.34477, 17.34478, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.3448, 17.3448, 17.34479, 17.34479, 17.34477, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34472, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.34479, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34478, 17.34478, 17.34477, 17.34476, 17.34474, 17.34473, 
    17.34472, 17.34473, 17.34472, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.34479, 17.3448, 
    17.3448, 17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34477, 
    17.34477, 17.34476, 17.34475, 17.34473, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 
    17.3447, 17.34471, 17.34479, 17.34479, 17.34479, 17.34479, 17.34479, 
    17.34478, 17.34477, 17.34475, 17.34476, 17.34475, 17.34476, 17.34476, 
    17.34475, 17.34476, 17.34473, 17.34475, 17.34472, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34471, 17.34471, 17.34469, 17.3447, 17.34469, 
    17.34478, 17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 
    17.34475, 17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 
    17.34477, 17.34478, 17.34475, 17.34476, 17.34473, 17.34474, 17.34471, 
    17.34473, 17.3447, 17.34469, 17.34468, 17.34466, 17.34477, 17.34478, 
    17.34477, 17.34476, 17.34475, 17.34474, 17.34474, 17.34474, 17.34473, 
    17.34473, 17.34474, 17.34472, 17.34477, 17.34475, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 
    17.34471, 17.34465, 17.34467, 17.34478, 17.34477, 17.34476, 17.34476, 
    17.34474, 17.34473, 17.34473, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34474, 17.34473, 17.34476, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 
    17.34472, 17.34477, 17.34476, 17.34476, 17.34476, 17.34473, 17.34474, 
    17.34472, 17.34472, 17.34471, 17.34472, 17.34472, 17.34473, 17.34473, 
    17.34474, 17.34475, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34474, 17.34473, 17.34473, 17.34472, 17.34475, 
    17.34473, 17.34475, 17.34475, 17.34474, 17.34473, 17.34473, 17.34472, 
    17.34472, 17.34473, 17.34474, 17.34474, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34475, 17.34473, 17.34472, 17.34471, 17.34471, 17.34469, 
    17.34471, 17.34469, 17.3447, 17.34468, 17.34472, 17.3447, 17.34474, 
    17.34474, 17.34473, 17.34471, 17.34472, 17.34471, 17.34474, 17.34475, 
    17.34475, 17.34476, 17.34475, 17.34475, 17.34475, 17.34475, 17.34473, 
    17.34474, 17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34465, 
    17.34465, 17.34465 ;

 TOTSOMN =
  1.773786, 1.773784, 1.773785, 1.773783, 1.773784, 1.773783, 1.773786, 
    1.773784, 1.773785, 1.773786, 1.77378, 1.773783, 1.773777, 1.773779, 
    1.773775, 1.773778, 1.773774, 1.773775, 1.773773, 1.773773, 1.773771, 
    1.773772, 1.773769, 1.773771, 1.773771, 1.773772, 1.773782, 1.773781, 
    1.773783, 1.773782, 1.773782, 1.773784, 1.773785, 1.773786, 1.773786, 
    1.773785, 1.773782, 1.773783, 1.773781, 1.773781, 1.773778, 1.77378, 
    1.773775, 1.773777, 1.773773, 1.773774, 1.773773, 1.773773, 1.773773, 
    1.773775, 1.773774, 1.773775, 1.773779, 1.773778, 1.773782, 1.773784, 
    1.773786, 1.773787, 1.773787, 1.773786, 1.773785, 1.773783, 1.773782, 
    1.773782, 1.773781, 1.773779, 1.773778, 1.773775, 1.773776, 1.773775, 
    1.773774, 1.773773, 1.773773, 1.773772, 1.773775, 1.773773, 1.773776, 
    1.773775, 1.773781, 1.773783, 1.773784, 1.773785, 1.773786, 1.773785, 
    1.773786, 1.773784, 1.773784, 1.773784, 1.773782, 1.773782, 1.773778, 
    1.77378, 1.773774, 1.773775, 1.773774, 1.773775, 1.773773, 1.773775, 
    1.773772, 1.773772, 1.773772, 1.773771, 1.773775, 1.773773, 1.773784, 
    1.773784, 1.773784, 1.773785, 1.773785, 1.773786, 1.773785, 1.773785, 
    1.773784, 1.773783, 1.773782, 1.773781, 1.773779, 1.773777, 1.773775, 
    1.773774, 1.773775, 1.773774, 1.773775, 1.773775, 1.773772, 1.773774, 
    1.773771, 1.773771, 1.773772, 1.773771, 1.773784, 1.773784, 1.773786, 
    1.773785, 1.773786, 1.773785, 1.773785, 1.773782, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773777, 1.773776, 1.773774, 1.773774, 1.773774, 
    1.773774, 1.773775, 1.773774, 1.773773, 1.773774, 1.773771, 1.773772, 
    1.773771, 1.773772, 1.773784, 1.773784, 1.773784, 1.773783, 1.773784, 
    1.773782, 1.773781, 1.773778, 1.77378, 1.773778, 1.773779, 1.773779, 
    1.773778, 1.773779, 1.773776, 1.773778, 1.773774, 1.773776, 1.773774, 
    1.773774, 1.773773, 1.773773, 1.773772, 1.77377, 1.773771, 1.773769, 
    1.773783, 1.773782, 1.773782, 1.773781, 1.77378, 1.773779, 1.773777, 
    1.773778, 1.773776, 1.773776, 1.773778, 1.773777, 1.773781, 1.773781, 
    1.773781, 1.773783, 1.773778, 1.77378, 1.773775, 1.773777, 1.773773, 
    1.773775, 1.773771, 1.773769, 1.773767, 1.773766, 1.773781, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773777, 1.773777, 1.773776, 1.773775, 
    1.773775, 1.773776, 1.773775, 1.77378, 1.773777, 1.773782, 1.773781, 
    1.77378, 1.77378, 1.773778, 1.773777, 1.773775, 1.773776, 1.773769, 
    1.773772, 1.773764, 1.773767, 1.773782, 1.773781, 1.773779, 1.77378, 
    1.773777, 1.773776, 1.773775, 1.773774, 1.773774, 1.773774, 1.773774, 
    1.773774, 1.773777, 1.773775, 1.773779, 1.773778, 1.773779, 1.773779, 
    1.773778, 1.773776, 1.773776, 1.773776, 1.773774, 1.773777, 1.773769, 
    1.773774, 1.773781, 1.773779, 1.773779, 1.77378, 1.773776, 1.773777, 
    1.773774, 1.773775, 1.773773, 1.773774, 1.773774, 1.773775, 1.773775, 
    1.773777, 1.773778, 1.77378, 1.773779, 1.773778, 1.773776, 1.773774, 
    1.773775, 1.773773, 1.773777, 1.773775, 1.773776, 1.773774, 1.773778, 
    1.773775, 1.773779, 1.773778, 1.773777, 1.773775, 1.773775, 1.773774, 
    1.773775, 1.773776, 1.773776, 1.773777, 1.773777, 1.773778, 1.773779, 
    1.773778, 1.773778, 1.773776, 1.773774, 1.773773, 1.773772, 1.77377, 
    1.773772, 1.773769, 1.773771, 1.773767, 1.773775, 1.773772, 1.773777, 
    1.773777, 1.773775, 1.773773, 1.773774, 1.773773, 1.773776, 1.773778, 
    1.773779, 1.773779, 1.773778, 1.773779, 1.773778, 1.773778, 1.773776, 
    1.773777, 1.773774, 1.773773, 1.773769, 1.773767, 1.773765, 1.773764, 
    1.773764, 1.773764 ;

 TOTSOMN_1m =
  1.773786, 1.773784, 1.773785, 1.773783, 1.773784, 1.773783, 1.773786, 
    1.773784, 1.773785, 1.773786, 1.77378, 1.773783, 1.773777, 1.773779, 
    1.773775, 1.773778, 1.773774, 1.773775, 1.773773, 1.773773, 1.773771, 
    1.773772, 1.773769, 1.773771, 1.773771, 1.773772, 1.773782, 1.773781, 
    1.773783, 1.773782, 1.773782, 1.773784, 1.773785, 1.773786, 1.773786, 
    1.773785, 1.773782, 1.773783, 1.773781, 1.773781, 1.773778, 1.77378, 
    1.773775, 1.773777, 1.773773, 1.773774, 1.773773, 1.773773, 1.773773, 
    1.773775, 1.773774, 1.773775, 1.773779, 1.773778, 1.773782, 1.773784, 
    1.773786, 1.773787, 1.773787, 1.773786, 1.773785, 1.773783, 1.773782, 
    1.773782, 1.773781, 1.773779, 1.773778, 1.773775, 1.773776, 1.773775, 
    1.773774, 1.773773, 1.773773, 1.773772, 1.773775, 1.773773, 1.773776, 
    1.773775, 1.773781, 1.773783, 1.773784, 1.773785, 1.773786, 1.773785, 
    1.773786, 1.773784, 1.773784, 1.773784, 1.773782, 1.773782, 1.773778, 
    1.77378, 1.773774, 1.773775, 1.773774, 1.773775, 1.773773, 1.773775, 
    1.773772, 1.773772, 1.773772, 1.773771, 1.773775, 1.773773, 1.773784, 
    1.773784, 1.773784, 1.773785, 1.773785, 1.773786, 1.773785, 1.773785, 
    1.773784, 1.773783, 1.773782, 1.773781, 1.773779, 1.773777, 1.773775, 
    1.773774, 1.773775, 1.773774, 1.773775, 1.773775, 1.773772, 1.773774, 
    1.773771, 1.773771, 1.773772, 1.773771, 1.773784, 1.773784, 1.773786, 
    1.773785, 1.773786, 1.773785, 1.773785, 1.773782, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773777, 1.773776, 1.773774, 1.773774, 1.773774, 
    1.773774, 1.773775, 1.773774, 1.773773, 1.773774, 1.773771, 1.773772, 
    1.773771, 1.773772, 1.773784, 1.773784, 1.773784, 1.773783, 1.773784, 
    1.773782, 1.773781, 1.773778, 1.77378, 1.773778, 1.773779, 1.773779, 
    1.773778, 1.773779, 1.773776, 1.773778, 1.773774, 1.773776, 1.773774, 
    1.773774, 1.773773, 1.773773, 1.773772, 1.77377, 1.773771, 1.773769, 
    1.773783, 1.773782, 1.773782, 1.773781, 1.77378, 1.773779, 1.773777, 
    1.773778, 1.773776, 1.773776, 1.773778, 1.773777, 1.773781, 1.773781, 
    1.773781, 1.773783, 1.773778, 1.77378, 1.773775, 1.773777, 1.773773, 
    1.773775, 1.773771, 1.773769, 1.773767, 1.773766, 1.773781, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773777, 1.773777, 1.773776, 1.773775, 
    1.773775, 1.773776, 1.773775, 1.77378, 1.773777, 1.773782, 1.773781, 
    1.77378, 1.77378, 1.773778, 1.773777, 1.773775, 1.773776, 1.773769, 
    1.773772, 1.773764, 1.773767, 1.773782, 1.773781, 1.773779, 1.77378, 
    1.773777, 1.773776, 1.773775, 1.773774, 1.773774, 1.773774, 1.773774, 
    1.773774, 1.773777, 1.773775, 1.773779, 1.773778, 1.773779, 1.773779, 
    1.773778, 1.773776, 1.773776, 1.773776, 1.773774, 1.773777, 1.773769, 
    1.773774, 1.773781, 1.773779, 1.773779, 1.77378, 1.773776, 1.773777, 
    1.773774, 1.773775, 1.773773, 1.773774, 1.773774, 1.773775, 1.773775, 
    1.773777, 1.773778, 1.77378, 1.773779, 1.773778, 1.773776, 1.773774, 
    1.773775, 1.773773, 1.773777, 1.773775, 1.773776, 1.773774, 1.773778, 
    1.773775, 1.773779, 1.773778, 1.773777, 1.773775, 1.773775, 1.773774, 
    1.773775, 1.773776, 1.773776, 1.773777, 1.773777, 1.773778, 1.773779, 
    1.773778, 1.773778, 1.773776, 1.773774, 1.773773, 1.773772, 1.77377, 
    1.773772, 1.773769, 1.773771, 1.773767, 1.773775, 1.773772, 1.773777, 
    1.773777, 1.773775, 1.773773, 1.773774, 1.773773, 1.773776, 1.773778, 
    1.773779, 1.773779, 1.773778, 1.773779, 1.773778, 1.773778, 1.773776, 
    1.773777, 1.773774, 1.773773, 1.773769, 1.773767, 1.773765, 1.773764, 
    1.773764, 1.773764 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  249.9696, 249.9699, 249.9698, 249.9701, 249.9699, 249.9701, 249.9697, 
    249.9699, 249.9698, 249.9697, 249.9704, 249.9701, 249.9709, 249.9706, 
    249.9713, 249.9708, 249.9713, 249.9713, 249.9715, 249.9715, 249.9718, 
    249.9716, 249.972, 249.9718, 249.9718, 249.9716, 249.9702, 249.9704, 
    249.9701, 249.9702, 249.9702, 249.9699, 249.9698, 249.9696, 249.9697, 
    249.9698, 249.9702, 249.9701, 249.9704, 249.9704, 249.9707, 249.9706, 
    249.9711, 249.971, 249.9715, 249.9713, 249.9715, 249.9714, 249.9715, 
    249.9713, 249.9714, 249.9712, 249.9706, 249.9708, 249.9702, 249.9699, 
    249.9697, 249.9696, 249.9696, 249.9696, 249.9698, 249.97, 249.9702, 
    249.9703, 249.9704, 249.9707, 249.9708, 249.9712, 249.9711, 249.9712, 
    249.9713, 249.9715, 249.9715, 249.9716, 249.9712, 249.9714, 249.9711, 
    249.9712, 249.9704, 249.9701, 249.97, 249.9699, 249.9696, 249.9698, 
    249.9697, 249.9699, 249.97, 249.9699, 249.9703, 249.9701, 249.9708, 
    249.9705, 249.9713, 249.9711, 249.9714, 249.9713, 249.9715, 249.9713, 
    249.9716, 249.9716, 249.9716, 249.9718, 249.9713, 249.9715, 249.9699, 
    249.9699, 249.97, 249.9698, 249.9698, 249.9696, 249.9698, 249.9698, 
    249.97, 249.9701, 249.9702, 249.9704, 249.9706, 249.9709, 249.9711, 
    249.9713, 249.9712, 249.9713, 249.9712, 249.9711, 249.9716, 249.9714, 
    249.9718, 249.9717, 249.9716, 249.9717, 249.9699, 249.9699, 249.9697, 
    249.9699, 249.9696, 249.9697, 249.9698, 249.9701, 249.9702, 249.9703, 
    249.9704, 249.9706, 249.9709, 249.9711, 249.9713, 249.9713, 249.9713, 
    249.9714, 249.9713, 249.9714, 249.9714, 249.9714, 249.9717, 249.9716, 
    249.9717, 249.9717, 249.9699, 249.97, 249.97, 249.97, 249.97, 249.9702, 
    249.9703, 249.9707, 249.9706, 249.9708, 249.9706, 249.9706, 249.9708, 
    249.9706, 249.9711, 249.9707, 249.9714, 249.971, 249.9714, 249.9713, 
    249.9715, 249.9715, 249.9717, 249.9719, 249.9718, 249.972, 249.9701, 
    249.9702, 249.9702, 249.9704, 249.9704, 249.9706, 249.9709, 249.9708, 
    249.971, 249.9711, 249.9707, 249.9709, 249.9703, 249.9704, 249.9704, 
    249.9701, 249.9708, 249.9705, 249.9711, 249.9709, 249.9715, 249.9712, 
    249.9718, 249.972, 249.9723, 249.9725, 249.9703, 249.9702, 249.9704, 
    249.9706, 249.9707, 249.971, 249.971, 249.971, 249.9711, 249.9712, 
    249.971, 249.9713, 249.9704, 249.9709, 249.9702, 249.9704, 249.9705, 
    249.9705, 249.9708, 249.9709, 249.9712, 249.971, 249.972, 249.9716, 
    249.9727, 249.9724, 249.9702, 249.9703, 249.9707, 249.9705, 249.971, 
    249.9711, 249.9712, 249.9713, 249.9713, 249.9714, 249.9713, 249.9714, 
    249.971, 249.9712, 249.9706, 249.9707, 249.9707, 249.9706, 249.9708, 
    249.971, 249.9711, 249.9711, 249.9713, 249.971, 249.972, 249.9714, 
    249.9704, 249.9706, 249.9706, 249.9706, 249.9711, 249.9709, 249.9714, 
    249.9713, 249.9715, 249.9714, 249.9714, 249.9712, 249.9711, 249.9709, 
    249.9707, 249.9706, 249.9706, 249.9708, 249.9711, 249.9713, 249.9713, 
    249.9715, 249.9709, 249.9712, 249.9711, 249.9713, 249.9708, 249.9712, 
    249.9707, 249.9707, 249.9709, 249.9712, 249.9713, 249.9713, 249.9713, 
    249.9711, 249.971, 249.9709, 249.9709, 249.9707, 249.9707, 249.9707, 
    249.9708, 249.9711, 249.9713, 249.9715, 249.9716, 249.9719, 249.9716, 
    249.972, 249.9717, 249.9723, 249.9713, 249.9717, 249.9709, 249.971, 
    249.9711, 249.9715, 249.9713, 249.9715, 249.971, 249.9708, 249.9707, 
    249.9706, 249.9707, 249.9707, 249.9708, 249.9708, 249.9711, 249.9709, 
    249.9714, 249.9715, 249.972, 249.9723, 249.9726, 249.9727, 249.9727, 
    249.9727 ;

 TREFMNAV_R =
  249.9696, 249.9699, 249.9698, 249.9701, 249.9699, 249.9701, 249.9697, 
    249.9699, 249.9698, 249.9697, 249.9704, 249.9701, 249.9709, 249.9706, 
    249.9713, 249.9708, 249.9713, 249.9713, 249.9715, 249.9715, 249.9718, 
    249.9716, 249.972, 249.9718, 249.9718, 249.9716, 249.9702, 249.9704, 
    249.9701, 249.9702, 249.9702, 249.9699, 249.9698, 249.9696, 249.9697, 
    249.9698, 249.9702, 249.9701, 249.9704, 249.9704, 249.9707, 249.9706, 
    249.9711, 249.971, 249.9715, 249.9713, 249.9715, 249.9714, 249.9715, 
    249.9713, 249.9714, 249.9712, 249.9706, 249.9708, 249.9702, 249.9699, 
    249.9697, 249.9696, 249.9696, 249.9696, 249.9698, 249.97, 249.9702, 
    249.9703, 249.9704, 249.9707, 249.9708, 249.9712, 249.9711, 249.9712, 
    249.9713, 249.9715, 249.9715, 249.9716, 249.9712, 249.9714, 249.9711, 
    249.9712, 249.9704, 249.9701, 249.97, 249.9699, 249.9696, 249.9698, 
    249.9697, 249.9699, 249.97, 249.9699, 249.9703, 249.9701, 249.9708, 
    249.9705, 249.9713, 249.9711, 249.9714, 249.9713, 249.9715, 249.9713, 
    249.9716, 249.9716, 249.9716, 249.9718, 249.9713, 249.9715, 249.9699, 
    249.9699, 249.97, 249.9698, 249.9698, 249.9696, 249.9698, 249.9698, 
    249.97, 249.9701, 249.9702, 249.9704, 249.9706, 249.9709, 249.9711, 
    249.9713, 249.9712, 249.9713, 249.9712, 249.9711, 249.9716, 249.9714, 
    249.9718, 249.9717, 249.9716, 249.9717, 249.9699, 249.9699, 249.9697, 
    249.9699, 249.9696, 249.9697, 249.9698, 249.9701, 249.9702, 249.9703, 
    249.9704, 249.9706, 249.9709, 249.9711, 249.9713, 249.9713, 249.9713, 
    249.9714, 249.9713, 249.9714, 249.9714, 249.9714, 249.9717, 249.9716, 
    249.9717, 249.9717, 249.9699, 249.97, 249.97, 249.97, 249.97, 249.9702, 
    249.9703, 249.9707, 249.9706, 249.9708, 249.9706, 249.9706, 249.9708, 
    249.9706, 249.9711, 249.9707, 249.9714, 249.971, 249.9714, 249.9713, 
    249.9715, 249.9715, 249.9717, 249.9719, 249.9718, 249.972, 249.9701, 
    249.9702, 249.9702, 249.9704, 249.9704, 249.9706, 249.9709, 249.9708, 
    249.971, 249.9711, 249.9707, 249.9709, 249.9703, 249.9704, 249.9704, 
    249.9701, 249.9708, 249.9705, 249.9711, 249.9709, 249.9715, 249.9712, 
    249.9718, 249.972, 249.9723, 249.9725, 249.9703, 249.9702, 249.9704, 
    249.9706, 249.9707, 249.971, 249.971, 249.971, 249.9711, 249.9712, 
    249.971, 249.9713, 249.9704, 249.9709, 249.9702, 249.9704, 249.9705, 
    249.9705, 249.9708, 249.9709, 249.9712, 249.971, 249.972, 249.9716, 
    249.9727, 249.9724, 249.9702, 249.9703, 249.9707, 249.9705, 249.971, 
    249.9711, 249.9712, 249.9713, 249.9713, 249.9714, 249.9713, 249.9714, 
    249.971, 249.9712, 249.9706, 249.9707, 249.9707, 249.9706, 249.9708, 
    249.971, 249.9711, 249.9711, 249.9713, 249.971, 249.972, 249.9714, 
    249.9704, 249.9706, 249.9706, 249.9706, 249.9711, 249.9709, 249.9714, 
    249.9713, 249.9715, 249.9714, 249.9714, 249.9712, 249.9711, 249.9709, 
    249.9707, 249.9706, 249.9706, 249.9708, 249.9711, 249.9713, 249.9713, 
    249.9715, 249.9709, 249.9712, 249.9711, 249.9713, 249.9708, 249.9712, 
    249.9707, 249.9707, 249.9709, 249.9712, 249.9713, 249.9713, 249.9713, 
    249.9711, 249.971, 249.9709, 249.9709, 249.9707, 249.9707, 249.9707, 
    249.9708, 249.9711, 249.9713, 249.9715, 249.9716, 249.9719, 249.9716, 
    249.972, 249.9717, 249.9723, 249.9713, 249.9717, 249.9709, 249.971, 
    249.9711, 249.9715, 249.9713, 249.9715, 249.971, 249.9708, 249.9707, 
    249.9706, 249.9707, 249.9707, 249.9708, 249.9708, 249.9711, 249.9709, 
    249.9714, 249.9715, 249.972, 249.9723, 249.9726, 249.9727, 249.9727, 
    249.9727 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  258.5157, 258.5161, 258.516, 258.5164, 258.5162, 258.5164, 258.5158, 
    258.5161, 258.5159, 258.5157, 258.517, 258.5164, 258.5176, 258.5172, 
    258.5182, 258.5175, 258.5184, 258.5182, 258.5187, 258.5186, 258.5191, 
    258.5187, 258.5194, 258.519, 258.5191, 258.5187, 258.5165, 258.5169, 
    258.5165, 258.5165, 258.5165, 258.5162, 258.516, 258.5157, 258.5157, 
    258.516, 258.5165, 258.5164, 258.5168, 258.5168, 258.5174, 258.5172, 
    258.5181, 258.5178, 258.5186, 258.5184, 258.5186, 258.5185, 258.5186, 
    258.5182, 258.5184, 258.5181, 258.5172, 258.5175, 258.5166, 258.5161, 
    258.5158, 258.5156, 258.5156, 258.5157, 258.516, 258.5163, 258.5165, 
    258.5167, 258.5168, 258.5173, 258.5175, 258.5181, 258.518, 258.5182, 
    258.5183, 258.5186, 258.5186, 258.5187, 258.5182, 258.5185, 258.5179, 
    258.5181, 258.5168, 258.5164, 258.5162, 258.5161, 258.5156, 258.5159, 
    258.5158, 258.5161, 258.5162, 258.5162, 258.5167, 258.5165, 258.5175, 
    258.5171, 258.5183, 258.518, 258.5184, 258.5182, 258.5185, 258.5182, 
    258.5187, 258.5188, 258.5188, 258.519, 258.5182, 258.5185, 258.5161, 
    258.5162, 258.5162, 258.516, 258.5159, 258.5157, 258.5159, 258.516, 
    258.5163, 258.5164, 258.5165, 258.5168, 258.5172, 258.5177, 258.518, 
    258.5183, 258.5181, 258.5183, 258.5181, 258.5181, 258.5188, 258.5184, 
    258.519, 258.519, 258.5187, 258.519, 258.5162, 258.5161, 258.5158, 
    258.5161, 258.5157, 258.5159, 258.516, 258.5165, 258.5166, 258.5167, 
    258.5169, 258.5172, 258.5176, 258.518, 258.5183, 258.5183, 258.5183, 
    258.5184, 258.5182, 258.5184, 258.5185, 258.5184, 258.519, 258.5188, 
    258.519, 258.5189, 258.5161, 258.5163, 258.5162, 258.5163, 258.5162, 
    258.5167, 258.5168, 258.5174, 258.5172, 258.5175, 258.5172, 258.5172, 
    258.5175, 258.5172, 258.518, 258.5175, 258.5184, 258.5179, 258.5185, 
    258.5183, 258.5185, 258.5187, 258.5189, 258.5192, 258.5191, 258.5194, 
    258.5165, 258.5166, 258.5166, 258.5168, 258.5169, 258.5172, 258.5177, 
    258.5175, 258.5179, 258.5179, 258.5174, 258.5177, 258.5168, 258.5169, 
    258.5168, 258.5165, 258.5176, 258.517, 258.5181, 258.5178, 258.5186, 
    258.5182, 258.5191, 258.5194, 258.5198, 258.5202, 258.5167, 258.5166, 
    258.5168, 258.5171, 258.5174, 258.5178, 258.5178, 258.5179, 258.5181, 
    258.5182, 258.5179, 258.5182, 258.5169, 258.5176, 258.5166, 258.5169, 
    258.5171, 258.517, 258.5175, 258.5176, 258.5181, 258.5179, 258.5193, 
    258.5187, 258.5205, 258.52, 258.5166, 258.5167, 258.5173, 258.517, 
    258.5178, 258.518, 258.5181, 258.5183, 258.5183, 258.5185, 258.5183, 
    258.5185, 258.5178, 258.5181, 258.5172, 258.5174, 258.5173, 258.5172, 
    258.5175, 258.5179, 258.5179, 258.518, 258.5183, 258.5178, 258.5194, 
    258.5184, 258.5169, 258.5172, 258.5173, 258.5172, 258.5179, 258.5177, 
    258.5185, 258.5182, 258.5186, 258.5184, 258.5184, 258.5182, 258.518, 
    258.5177, 258.5174, 258.5172, 258.5172, 258.5175, 258.5179, 258.5183, 
    258.5182, 258.5186, 258.5177, 258.5181, 258.5179, 258.5183, 258.5175, 
    258.5182, 258.5174, 258.5174, 258.5177, 258.5181, 258.5182, 258.5183, 
    258.5182, 258.5179, 258.5179, 258.5176, 258.5176, 258.5174, 258.5173, 
    258.5174, 258.5175, 258.5179, 258.5183, 258.5187, 258.5188, 258.5192, 
    258.5188, 258.5194, 258.5189, 258.5198, 258.5182, 258.5189, 258.5177, 
    258.5178, 258.518, 258.5186, 258.5183, 258.5186, 258.5179, 258.5175, 
    258.5174, 258.5172, 258.5174, 258.5174, 258.5175, 258.5175, 258.5179, 
    258.5177, 258.5184, 258.5186, 258.5194, 258.5198, 258.5203, 258.5205, 
    258.5205, 258.5205 ;

 TREFMXAV_R =
  258.5157, 258.5161, 258.516, 258.5164, 258.5162, 258.5164, 258.5158, 
    258.5161, 258.5159, 258.5157, 258.517, 258.5164, 258.5176, 258.5172, 
    258.5182, 258.5175, 258.5184, 258.5182, 258.5187, 258.5186, 258.5191, 
    258.5187, 258.5194, 258.519, 258.5191, 258.5187, 258.5165, 258.5169, 
    258.5165, 258.5165, 258.5165, 258.5162, 258.516, 258.5157, 258.5157, 
    258.516, 258.5165, 258.5164, 258.5168, 258.5168, 258.5174, 258.5172, 
    258.5181, 258.5178, 258.5186, 258.5184, 258.5186, 258.5185, 258.5186, 
    258.5182, 258.5184, 258.5181, 258.5172, 258.5175, 258.5166, 258.5161, 
    258.5158, 258.5156, 258.5156, 258.5157, 258.516, 258.5163, 258.5165, 
    258.5167, 258.5168, 258.5173, 258.5175, 258.5181, 258.518, 258.5182, 
    258.5183, 258.5186, 258.5186, 258.5187, 258.5182, 258.5185, 258.5179, 
    258.5181, 258.5168, 258.5164, 258.5162, 258.5161, 258.5156, 258.5159, 
    258.5158, 258.5161, 258.5162, 258.5162, 258.5167, 258.5165, 258.5175, 
    258.5171, 258.5183, 258.518, 258.5184, 258.5182, 258.5185, 258.5182, 
    258.5187, 258.5188, 258.5188, 258.519, 258.5182, 258.5185, 258.5161, 
    258.5162, 258.5162, 258.516, 258.5159, 258.5157, 258.5159, 258.516, 
    258.5163, 258.5164, 258.5165, 258.5168, 258.5172, 258.5177, 258.518, 
    258.5183, 258.5181, 258.5183, 258.5181, 258.5181, 258.5188, 258.5184, 
    258.519, 258.519, 258.5187, 258.519, 258.5162, 258.5161, 258.5158, 
    258.5161, 258.5157, 258.5159, 258.516, 258.5165, 258.5166, 258.5167, 
    258.5169, 258.5172, 258.5176, 258.518, 258.5183, 258.5183, 258.5183, 
    258.5184, 258.5182, 258.5184, 258.5185, 258.5184, 258.519, 258.5188, 
    258.519, 258.5189, 258.5161, 258.5163, 258.5162, 258.5163, 258.5162, 
    258.5167, 258.5168, 258.5174, 258.5172, 258.5175, 258.5172, 258.5172, 
    258.5175, 258.5172, 258.518, 258.5175, 258.5184, 258.5179, 258.5185, 
    258.5183, 258.5185, 258.5187, 258.5189, 258.5192, 258.5191, 258.5194, 
    258.5165, 258.5166, 258.5166, 258.5168, 258.5169, 258.5172, 258.5177, 
    258.5175, 258.5179, 258.5179, 258.5174, 258.5177, 258.5168, 258.5169, 
    258.5168, 258.5165, 258.5176, 258.517, 258.5181, 258.5178, 258.5186, 
    258.5182, 258.5191, 258.5194, 258.5198, 258.5202, 258.5167, 258.5166, 
    258.5168, 258.5171, 258.5174, 258.5178, 258.5178, 258.5179, 258.5181, 
    258.5182, 258.5179, 258.5182, 258.5169, 258.5176, 258.5166, 258.5169, 
    258.5171, 258.517, 258.5175, 258.5176, 258.5181, 258.5179, 258.5193, 
    258.5187, 258.5205, 258.52, 258.5166, 258.5167, 258.5173, 258.517, 
    258.5178, 258.518, 258.5181, 258.5183, 258.5183, 258.5185, 258.5183, 
    258.5185, 258.5178, 258.5181, 258.5172, 258.5174, 258.5173, 258.5172, 
    258.5175, 258.5179, 258.5179, 258.518, 258.5183, 258.5178, 258.5194, 
    258.5184, 258.5169, 258.5172, 258.5173, 258.5172, 258.5179, 258.5177, 
    258.5185, 258.5182, 258.5186, 258.5184, 258.5184, 258.5182, 258.518, 
    258.5177, 258.5174, 258.5172, 258.5172, 258.5175, 258.5179, 258.5183, 
    258.5182, 258.5186, 258.5177, 258.5181, 258.5179, 258.5183, 258.5175, 
    258.5182, 258.5174, 258.5174, 258.5177, 258.5181, 258.5182, 258.5183, 
    258.5182, 258.5179, 258.5179, 258.5176, 258.5176, 258.5174, 258.5173, 
    258.5174, 258.5175, 258.5179, 258.5183, 258.5187, 258.5188, 258.5192, 
    258.5188, 258.5194, 258.5189, 258.5198, 258.5182, 258.5189, 258.5177, 
    258.5178, 258.518, 258.5186, 258.5183, 258.5186, 258.5179, 258.5175, 
    258.5174, 258.5172, 258.5174, 258.5174, 258.5175, 258.5175, 258.5179, 
    258.5177, 258.5184, 258.5186, 258.5194, 258.5198, 258.5203, 258.5205, 
    258.5205, 258.5205 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  253.9562, 253.9564, 253.9564, 253.9565, 253.9565, 253.9565, 253.9563, 
    253.9564, 253.9563, 253.9563, 253.9568, 253.9565, 253.9571, 253.9569, 
    253.9573, 253.957, 253.9574, 253.9573, 253.9575, 253.9575, 253.9577, 
    253.9576, 253.9579, 253.9577, 253.9577, 253.9576, 253.9566, 253.9568, 
    253.9566, 253.9566, 253.9566, 253.9565, 253.9564, 253.9562, 253.9563, 
    253.9564, 253.9566, 253.9565, 253.9567, 253.9567, 253.957, 253.9569, 
    253.9573, 253.9571, 253.9575, 253.9574, 253.9575, 253.9574, 253.9575, 
    253.9574, 253.9574, 253.9573, 253.9569, 253.957, 253.9566, 253.9564, 
    253.9563, 253.9562, 253.9562, 253.9562, 253.9564, 253.9565, 253.9566, 
    253.9567, 253.9567, 253.9569, 253.957, 253.9573, 253.9572, 253.9573, 
    253.9574, 253.9575, 253.9575, 253.9575, 253.9573, 253.9575, 253.9572, 
    253.9573, 253.9567, 253.9565, 253.9565, 253.9564, 253.9562, 253.9563, 
    253.9563, 253.9564, 253.9565, 253.9564, 253.9567, 253.9566, 253.957, 
    253.9568, 253.9574, 253.9572, 253.9574, 253.9573, 253.9575, 253.9573, 
    253.9576, 253.9576, 253.9576, 253.9577, 253.9573, 253.9575, 253.9564, 
    253.9565, 253.9565, 253.9563, 253.9563, 253.9562, 253.9563, 253.9564, 
    253.9565, 253.9565, 253.9566, 253.9567, 253.9569, 253.9571, 253.9572, 
    253.9574, 253.9573, 253.9574, 253.9573, 253.9573, 253.9576, 253.9574, 
    253.9577, 253.9577, 253.9575, 253.9577, 253.9565, 253.9564, 253.9563, 
    253.9564, 253.9562, 253.9563, 253.9564, 253.9566, 253.9566, 253.9567, 
    253.9568, 253.9569, 253.9571, 253.9572, 253.9574, 253.9574, 253.9574, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9577, 253.9576, 
    253.9577, 253.9576, 253.9564, 253.9565, 253.9565, 253.9565, 253.9565, 
    253.9566, 253.9567, 253.957, 253.9569, 253.957, 253.9569, 253.9569, 
    253.957, 253.9569, 253.9572, 253.957, 253.9574, 253.9572, 253.9574, 
    253.9574, 253.9575, 253.9575, 253.9576, 253.9577, 253.9577, 253.9578, 
    253.9566, 253.9566, 253.9566, 253.9567, 253.9568, 253.9569, 253.9571, 
    253.957, 253.9572, 253.9572, 253.957, 253.9571, 253.9567, 253.9568, 
    253.9567, 253.9566, 253.957, 253.9568, 253.9573, 253.9571, 253.9575, 
    253.9573, 253.9577, 253.9579, 253.958, 253.9582, 253.9567, 253.9566, 
    253.9567, 253.9568, 253.957, 253.9571, 253.9572, 253.9572, 253.9573, 
    253.9573, 253.9572, 253.9573, 253.9568, 253.9571, 253.9566, 253.9568, 
    253.9568, 253.9568, 253.957, 253.9571, 253.9573, 253.9572, 253.9578, 
    253.9575, 253.9583, 253.9581, 253.9566, 253.9567, 253.9569, 253.9568, 
    253.9571, 253.9572, 253.9573, 253.9574, 253.9574, 253.9574, 253.9574, 
    253.9574, 253.9571, 253.9573, 253.9569, 253.957, 253.957, 253.9569, 
    253.957, 253.9572, 253.9572, 253.9572, 253.9574, 253.9571, 253.9578, 
    253.9574, 253.9568, 253.9569, 253.9569, 253.9569, 253.9572, 253.9571, 
    253.9574, 253.9573, 253.9575, 253.9574, 253.9574, 253.9573, 253.9572, 
    253.9571, 253.957, 253.9569, 253.9569, 253.957, 253.9572, 253.9574, 
    253.9573, 253.9575, 253.9571, 253.9573, 253.9572, 253.9574, 253.957, 
    253.9573, 253.957, 253.957, 253.9571, 253.9573, 253.9573, 253.9574, 
    253.9573, 253.9572, 253.9572, 253.9571, 253.9571, 253.957, 253.9569, 
    253.957, 253.957, 253.9572, 253.9574, 253.9575, 253.9576, 253.9577, 
    253.9576, 253.9578, 253.9576, 253.958, 253.9573, 253.9576, 253.9571, 
    253.9572, 253.9572, 253.9575, 253.9574, 253.9575, 253.9572, 253.957, 
    253.957, 253.9569, 253.957, 253.957, 253.957, 253.957, 253.9572, 
    253.9571, 253.9574, 253.9575, 253.9578, 253.958, 253.9582, 253.9583, 
    253.9583, 253.9583 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  253.9562, 253.9564, 253.9564, 253.9565, 253.9565, 253.9565, 253.9563, 
    253.9564, 253.9563, 253.9563, 253.9568, 253.9565, 253.9571, 253.9569, 
    253.9573, 253.957, 253.9574, 253.9573, 253.9575, 253.9575, 253.9577, 
    253.9576, 253.9579, 253.9577, 253.9577, 253.9576, 253.9566, 253.9568, 
    253.9566, 253.9566, 253.9566, 253.9565, 253.9564, 253.9562, 253.9563, 
    253.9564, 253.9566, 253.9565, 253.9567, 253.9567, 253.957, 253.9569, 
    253.9573, 253.9571, 253.9575, 253.9574, 253.9575, 253.9574, 253.9575, 
    253.9574, 253.9574, 253.9573, 253.9569, 253.957, 253.9566, 253.9564, 
    253.9563, 253.9562, 253.9562, 253.9562, 253.9564, 253.9565, 253.9566, 
    253.9567, 253.9567, 253.9569, 253.957, 253.9573, 253.9572, 253.9573, 
    253.9574, 253.9575, 253.9575, 253.9575, 253.9573, 253.9575, 253.9572, 
    253.9573, 253.9567, 253.9565, 253.9565, 253.9564, 253.9562, 253.9563, 
    253.9563, 253.9564, 253.9565, 253.9564, 253.9567, 253.9566, 253.957, 
    253.9568, 253.9574, 253.9572, 253.9574, 253.9573, 253.9575, 253.9573, 
    253.9576, 253.9576, 253.9576, 253.9577, 253.9573, 253.9575, 253.9564, 
    253.9565, 253.9565, 253.9563, 253.9563, 253.9562, 253.9563, 253.9564, 
    253.9565, 253.9565, 253.9566, 253.9567, 253.9569, 253.9571, 253.9572, 
    253.9574, 253.9573, 253.9574, 253.9573, 253.9573, 253.9576, 253.9574, 
    253.9577, 253.9577, 253.9575, 253.9577, 253.9565, 253.9564, 253.9563, 
    253.9564, 253.9562, 253.9563, 253.9564, 253.9566, 253.9566, 253.9567, 
    253.9568, 253.9569, 253.9571, 253.9572, 253.9574, 253.9574, 253.9574, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9577, 253.9576, 
    253.9577, 253.9576, 253.9564, 253.9565, 253.9565, 253.9565, 253.9565, 
    253.9566, 253.9567, 253.957, 253.9569, 253.957, 253.9569, 253.9569, 
    253.957, 253.9569, 253.9572, 253.957, 253.9574, 253.9572, 253.9574, 
    253.9574, 253.9575, 253.9575, 253.9576, 253.9577, 253.9577, 253.9578, 
    253.9566, 253.9566, 253.9566, 253.9567, 253.9568, 253.9569, 253.9571, 
    253.957, 253.9572, 253.9572, 253.957, 253.9571, 253.9567, 253.9568, 
    253.9567, 253.9566, 253.957, 253.9568, 253.9573, 253.9571, 253.9575, 
    253.9573, 253.9577, 253.9579, 253.958, 253.9582, 253.9567, 253.9566, 
    253.9567, 253.9568, 253.957, 253.9571, 253.9572, 253.9572, 253.9573, 
    253.9573, 253.9572, 253.9573, 253.9568, 253.9571, 253.9566, 253.9568, 
    253.9568, 253.9568, 253.957, 253.9571, 253.9573, 253.9572, 253.9578, 
    253.9575, 253.9583, 253.9581, 253.9566, 253.9567, 253.9569, 253.9568, 
    253.9571, 253.9572, 253.9573, 253.9574, 253.9574, 253.9574, 253.9574, 
    253.9574, 253.9571, 253.9573, 253.9569, 253.957, 253.957, 253.9569, 
    253.957, 253.9572, 253.9572, 253.9572, 253.9574, 253.9571, 253.9578, 
    253.9574, 253.9568, 253.9569, 253.9569, 253.9569, 253.9572, 253.9571, 
    253.9574, 253.9573, 253.9575, 253.9574, 253.9574, 253.9573, 253.9572, 
    253.9571, 253.957, 253.9569, 253.9569, 253.957, 253.9572, 253.9574, 
    253.9573, 253.9575, 253.9571, 253.9573, 253.9572, 253.9574, 253.957, 
    253.9573, 253.957, 253.957, 253.9571, 253.9573, 253.9573, 253.9574, 
    253.9573, 253.9572, 253.9572, 253.9571, 253.9571, 253.957, 253.9569, 
    253.957, 253.957, 253.9572, 253.9574, 253.9575, 253.9576, 253.9577, 
    253.9576, 253.9578, 253.9576, 253.958, 253.9573, 253.9576, 253.9571, 
    253.9572, 253.9572, 253.9575, 253.9574, 253.9575, 253.9572, 253.957, 
    253.957, 253.9569, 253.957, 253.957, 253.957, 253.957, 253.9572, 
    253.9571, 253.9574, 253.9575, 253.9578, 253.958, 253.9582, 253.9583, 
    253.9583, 253.9583 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  254.3913, 254.3927, 254.3925, 254.3936, 254.393, 254.3937, 254.3916, 
    254.3928, 254.392, 254.3914, 254.3958, 254.3937, 254.3982, 254.3968, 
    254.4003, 254.3979, 254.4008, 254.4003, 254.4019, 254.4014, 254.4035, 
    254.4021, 254.4046, 254.4032, 254.4034, 254.4021, 254.3941, 254.3955, 
    254.394, 254.3942, 254.3941, 254.393, 254.3924, 254.3912, 254.3914, 
    254.3923, 254.3943, 254.3937, 254.3954, 254.3954, 254.3973, 254.3964, 
    254.3997, 254.3988, 254.4015, 254.4008, 254.4014, 254.4012, 254.4014, 
    254.4004, 254.4009, 254.4, 254.3966, 254.3976, 254.3946, 254.3928, 
    254.3916, 254.3908, 254.3909, 254.3912, 254.3923, 254.3934, 254.3943, 
    254.3948, 254.3954, 254.397, 254.3979, 254.3999, 254.3995, 254.4001, 
    254.4007, 254.4017, 254.4015, 254.402, 254.4001, 254.4013, 254.3993, 
    254.3999, 254.3954, 254.3938, 254.3931, 254.3925, 254.391, 254.3921, 
    254.3916, 254.3926, 254.3932, 254.3929, 254.3948, 254.3941, 254.3979, 
    254.3963, 254.4007, 254.3996, 254.4009, 254.4002, 254.4014, 254.4004, 
    254.4021, 254.4025, 254.4022, 254.4033, 254.4003, 254.4014, 254.3929, 
    254.393, 254.3932, 254.3922, 254.3921, 254.3912, 254.392, 254.3924, 
    254.3933, 254.3938, 254.3943, 254.3954, 254.3967, 254.3984, 254.3997, 
    254.4005, 254.4, 254.4005, 254.3999, 254.3997, 254.4023, 254.4008, 
    254.4031, 254.403, 254.402, 254.403, 254.393, 254.3927, 254.3917, 
    254.3925, 254.3911, 254.3919, 254.3923, 254.3941, 254.3945, 254.3948, 
    254.3956, 254.3965, 254.3981, 254.3995, 254.4008, 254.4007, 254.4007, 
    254.401, 254.4003, 254.4011, 254.4012, 254.4009, 254.403, 254.4024, 
    254.403, 254.4026, 254.3928, 254.3933, 254.3931, 254.3935, 254.3932, 
    254.3947, 254.3951, 254.3973, 254.3964, 254.3978, 254.3966, 254.3968, 
    254.3978, 254.3967, 254.3994, 254.3975, 254.401, 254.3991, 254.4011, 
    254.4007, 254.4013, 254.4019, 254.4025, 254.4038, 254.4035, 254.4045, 
    254.394, 254.3946, 254.3946, 254.3952, 254.3957, 254.3968, 254.3985, 
    254.3978, 254.399, 254.3992, 254.3975, 254.3985, 254.3951, 254.3956, 
    254.3953, 254.3941, 254.3979, 254.3959, 254.3997, 254.3986, 254.4018, 
    254.4002, 254.4033, 254.4046, 254.4059, 254.4074, 254.395, 254.3946, 
    254.3953, 254.3963, 254.3974, 254.3987, 254.3988, 254.399, 254.3997, 
    254.4002, 254.3991, 254.4003, 254.3957, 254.3981, 254.3944, 254.3955, 
    254.3963, 254.396, 254.3978, 254.3982, 254.3999, 254.399, 254.4043, 
    254.4019, 254.4086, 254.4067, 254.3944, 254.395, 254.397, 254.396, 
    254.3988, 254.3994, 254.4, 254.4007, 254.4007, 254.4012, 254.4005, 
    254.4011, 254.3987, 254.3998, 254.3968, 254.3975, 254.3972, 254.3968, 
    254.3979, 254.3991, 254.3992, 254.3995, 254.4005, 254.3988, 254.4045, 
    254.4009, 254.3956, 254.3967, 254.3969, 254.3965, 254.3994, 254.3983, 
    254.4012, 254.4004, 254.4016, 254.401, 254.4009, 254.4001, 254.3996, 
    254.3983, 254.3973, 254.3965, 254.3967, 254.3976, 254.3992, 254.4007, 
    254.4004, 254.4016, 254.3986, 254.3998, 254.3993, 254.4006, 254.3978, 
    254.4001, 254.3972, 254.3975, 254.3983, 254.3999, 254.4003, 254.4006, 
    254.4004, 254.3992, 254.3991, 254.3983, 254.398, 254.3974, 254.3969, 
    254.3974, 254.3978, 254.3992, 254.4005, 254.4019, 254.4022, 254.4037, 
    254.4025, 254.4046, 254.4027, 254.4059, 254.4003, 254.4027, 254.3983, 
    254.3988, 254.3996, 254.4016, 254.4006, 254.4018, 254.399, 254.3976, 
    254.3972, 254.3966, 254.3973, 254.3972, 254.3979, 254.3977, 254.3993, 
    254.3984, 254.4009, 254.4018, 254.4044, 254.406, 254.4076, 254.4084, 
    254.4086, 254.4087,
  255.5014, 255.5029, 255.5026, 255.5038, 255.5031, 255.5039, 255.5017, 
    255.5029, 255.5021, 255.5015, 255.506, 255.5038, 255.5084, 255.507, 
    255.5107, 255.5082, 255.5112, 255.5106, 255.5123, 255.5118, 255.514, 
    255.5126, 255.5152, 255.5137, 255.5139, 255.5125, 255.5043, 255.5057, 
    255.5042, 255.5044, 255.5043, 255.5031, 255.5025, 255.5013, 255.5015, 
    255.5024, 255.5045, 255.5038, 255.5056, 255.5056, 255.5076, 255.5067, 
    255.51, 255.5091, 255.5119, 255.5112, 255.5118, 255.5116, 255.5118, 
    255.5108, 255.5112, 255.5103, 255.5068, 255.5078, 255.5048, 255.5029, 
    255.5017, 255.5009, 255.501, 255.5012, 255.5024, 255.5036, 255.5044, 
    255.505, 255.5056, 255.5072, 255.5081, 255.5102, 255.5099, 255.5105, 
    255.5111, 255.5121, 255.5119, 255.5124, 255.5105, 255.5117, 255.5097, 
    255.5102, 255.5056, 255.504, 255.5032, 255.5026, 255.5011, 255.5022, 
    255.5017, 255.5027, 255.5034, 255.5031, 255.505, 255.5042, 255.5082, 
    255.5065, 255.511, 255.5099, 255.5113, 255.5106, 255.5118, 255.5107, 
    255.5125, 255.5129, 255.5127, 255.5137, 255.5107, 255.5118, 255.5031, 
    255.5031, 255.5033, 255.5023, 255.5022, 255.5013, 255.5021, 255.5025, 
    255.5034, 255.504, 255.5045, 255.5056, 255.5069, 255.5087, 255.51, 
    255.5109, 255.5103, 255.5108, 255.5103, 255.51, 255.5128, 255.5112, 
    255.5136, 255.5134, 255.5124, 255.5135, 255.5031, 255.5029, 255.5018, 
    255.5026, 255.5012, 255.502, 255.5024, 255.5042, 255.5047, 255.505, 
    255.5058, 255.5067, 255.5083, 255.5098, 255.5111, 255.511, 255.5111, 
    255.5114, 255.5106, 255.5115, 255.5116, 255.5112, 255.5134, 255.5128, 
    255.5134, 255.513, 255.5029, 255.5034, 255.5032, 255.5037, 255.5033, 
    255.5049, 255.5053, 255.5076, 255.5067, 255.5081, 255.5068, 255.507, 
    255.5081, 255.5069, 255.5097, 255.5078, 255.5114, 255.5094, 255.5115, 
    255.5111, 255.5117, 255.5123, 255.513, 255.5143, 255.514, 255.515, 
    255.5042, 255.5048, 255.5048, 255.5054, 255.5059, 255.507, 255.5088, 
    255.5081, 255.5093, 255.5096, 255.5077, 255.5088, 255.5052, 255.5058, 
    255.5055, 255.5042, 255.5082, 255.5061, 255.51, 255.5089, 255.5122, 
    255.5105, 255.5138, 255.5152, 255.5165, 255.518, 255.5052, 255.5047, 
    255.5055, 255.5066, 255.5076, 255.509, 255.5091, 255.5094, 255.51, 
    255.5106, 255.5094, 255.5107, 255.5059, 255.5084, 255.5046, 255.5057, 
    255.5065, 255.5062, 255.508, 255.5085, 255.5102, 255.5093, 255.5148, 
    255.5124, 255.5192, 255.5173, 255.5046, 255.5052, 255.5072, 255.5062, 
    255.509, 255.5098, 255.5103, 255.511, 255.5111, 255.5115, 255.5108, 
    255.5115, 255.509, 255.5101, 255.507, 255.5077, 255.5074, 255.507, 
    255.5082, 255.5094, 255.5095, 255.5099, 255.5109, 255.5091, 255.5151, 
    255.5113, 255.5058, 255.5069, 255.5071, 255.5067, 255.5097, 255.5086, 
    255.5115, 255.5107, 255.5121, 255.5114, 255.5113, 255.5105, 255.5099, 
    255.5086, 255.5076, 255.5067, 255.5069, 255.5078, 255.5095, 255.5111, 
    255.5108, 255.5119, 255.5089, 255.5101, 255.5096, 255.511, 255.5081, 
    255.5104, 255.5075, 255.5077, 255.5086, 255.5102, 255.5106, 255.511, 
    255.5108, 255.5096, 255.5094, 255.5085, 255.5083, 255.5077, 255.5072, 
    255.5076, 255.5081, 255.5096, 255.5109, 255.5123, 255.5126, 255.5143, 
    255.5129, 255.5151, 255.5132, 255.5165, 255.5106, 255.5132, 255.5086, 
    255.5091, 255.51, 255.512, 255.5109, 255.5122, 255.5094, 255.5079, 
    255.5075, 255.5068, 255.5075, 255.5075, 255.5082, 255.5079, 255.5096, 
    255.5087, 255.5113, 255.5122, 255.5149, 255.5166, 255.5183, 255.519, 
    255.5193, 255.5194,
  257.1078, 257.1091, 257.1089, 257.1099, 257.1093, 257.11, 257.1081, 
    257.1091, 257.1085, 257.1079, 257.112, 257.11, 257.1142, 257.1129, 
    257.1162, 257.114, 257.1167, 257.1162, 257.1177, 257.1173, 257.1193, 
    257.118, 257.1203, 257.119, 257.1192, 257.1179, 257.1104, 257.1117, 
    257.1103, 257.1105, 257.1104, 257.1093, 257.1088, 257.1077, 257.1079, 
    257.1087, 257.1106, 257.11, 257.1116, 257.1115, 257.1134, 257.1125, 
    257.1156, 257.1147, 257.1173, 257.1167, 257.1173, 257.1171, 257.1173, 
    257.1163, 257.1167, 257.1159, 257.1127, 257.1136, 257.1108, 257.1092, 
    257.1081, 257.1073, 257.1074, 257.1076, 257.1087, 257.1097, 257.1105, 
    257.111, 257.1115, 257.113, 257.1139, 257.1158, 257.1155, 257.116, 
    257.1166, 257.1175, 257.1174, 257.1178, 257.116, 257.1172, 257.1153, 
    257.1158, 257.1116, 257.1101, 257.1094, 257.1089, 257.1075, 257.1085, 
    257.1081, 257.109, 257.1096, 257.1093, 257.1111, 257.1104, 257.114, 
    257.1124, 257.1165, 257.1155, 257.1168, 257.1161, 257.1172, 257.1162, 
    257.1179, 257.1183, 257.118, 257.119, 257.1162, 257.1173, 257.1093, 
    257.1093, 257.1095, 257.1086, 257.1085, 257.1077, 257.1084, 257.1088, 
    257.1096, 257.1101, 257.1106, 257.1116, 257.1128, 257.1144, 257.1156, 
    257.1164, 257.1159, 257.1163, 257.1159, 257.1156, 257.1182, 257.1167, 
    257.1189, 257.1188, 257.1178, 257.1188, 257.1093, 257.1091, 257.1082, 
    257.1089, 257.1076, 257.1083, 257.1087, 257.1104, 257.1107, 257.1111, 
    257.1117, 257.1126, 257.1141, 257.1154, 257.1166, 257.1165, 257.1166, 
    257.1169, 257.1162, 257.1169, 257.1171, 257.1167, 257.1187, 257.1182, 
    257.1188, 257.1184, 257.1092, 257.1096, 257.1094, 257.1098, 257.1095, 
    257.1109, 257.1114, 257.1134, 257.1125, 257.1139, 257.1127, 257.1129, 
    257.1139, 257.1128, 257.1153, 257.1136, 257.1169, 257.1151, 257.117, 
    257.1166, 257.1172, 257.1177, 257.1183, 257.1195, 257.1192, 257.1202, 
    257.1103, 257.1109, 257.1108, 257.1115, 257.1119, 257.1129, 257.1145, 
    257.1139, 257.115, 257.1152, 257.1135, 257.1145, 257.1113, 257.1118, 
    257.1115, 257.1103, 257.114, 257.1121, 257.1156, 257.1146, 257.1176, 
    257.1161, 257.1191, 257.1203, 257.1216, 257.123, 257.1112, 257.1108, 
    257.1115, 257.1125, 257.1134, 257.1147, 257.1148, 257.115, 257.1156, 
    257.1161, 257.1151, 257.1162, 257.1118, 257.1142, 257.1106, 257.1117, 
    257.1124, 257.1121, 257.1138, 257.1142, 257.1158, 257.115, 257.12, 
    257.1178, 257.1241, 257.1223, 257.1107, 257.1112, 257.113, 257.1122, 
    257.1147, 257.1154, 257.1159, 257.1165, 257.1166, 257.117, 257.1164, 
    257.117, 257.1147, 257.1157, 257.1129, 257.1135, 257.1132, 257.1129, 
    257.114, 257.1151, 257.1151, 257.1155, 257.1165, 257.1147, 257.1203, 
    257.1168, 257.1118, 257.1128, 257.1129, 257.1125, 257.1153, 257.1143, 
    257.117, 257.1163, 257.1175, 257.1169, 257.1168, 257.116, 257.1155, 
    257.1143, 257.1134, 257.1126, 257.1128, 257.1136, 257.1151, 257.1166, 
    257.1163, 257.1174, 257.1145, 257.1157, 257.1153, 257.1165, 257.1139, 
    257.116, 257.1133, 257.1135, 257.1143, 257.1158, 257.1161, 257.1165, 
    257.1163, 257.1152, 257.115, 257.1143, 257.114, 257.1135, 257.113, 
    257.1134, 257.1139, 257.1152, 257.1164, 257.1177, 257.118, 257.1195, 
    257.1183, 257.1203, 257.1185, 257.1216, 257.1162, 257.1185, 257.1143, 
    257.1148, 257.1156, 257.1175, 257.1165, 257.1176, 257.115, 257.1136, 
    257.1133, 257.1127, 257.1133, 257.1133, 257.1139, 257.1137, 257.1152, 
    257.1144, 257.1168, 257.1176, 257.1201, 257.1216, 257.1232, 257.1239, 
    257.1241, 257.1242,
  259.2219, 259.2228, 259.2226, 259.2234, 259.223, 259.2235, 259.222, 
    259.2228, 259.2224, 259.222, 259.2249, 259.2234, 259.2265, 259.2256, 
    259.228, 259.2263, 259.2284, 259.228, 259.2292, 259.2288, 259.2303, 
    259.2293, 259.2311, 259.23, 259.2302, 259.2292, 259.2238, 259.2247, 
    259.2237, 259.2238, 259.2238, 259.223, 259.2226, 259.2218, 259.2219, 
    259.2225, 259.2239, 259.2234, 259.2246, 259.2246, 259.2259, 259.2253, 
    259.2276, 259.2269, 259.2288, 259.2283, 259.2288, 259.2287, 259.2288, 
    259.2281, 259.2284, 259.2278, 259.2254, 259.2261, 259.2241, 259.2228, 
    259.2221, 259.2215, 259.2216, 259.2218, 259.2225, 259.2233, 259.2238, 
    259.2242, 259.2246, 259.2257, 259.2263, 259.2277, 259.2274, 259.2279, 
    259.2283, 259.229, 259.2289, 259.2292, 259.2279, 259.2287, 259.2273, 
    259.2277, 259.2246, 259.2236, 259.2231, 259.2227, 259.2217, 259.2224, 
    259.2221, 259.2227, 259.2231, 259.223, 259.2242, 259.2237, 259.2263, 
    259.2252, 259.2282, 259.2275, 259.2284, 259.228, 259.2288, 259.228, 
    259.2293, 259.2296, 259.2294, 259.2301, 259.228, 259.2288, 259.2229, 
    259.223, 259.2231, 259.2224, 259.2224, 259.2218, 259.2224, 259.2226, 
    259.2232, 259.2235, 259.2239, 259.2246, 259.2255, 259.2267, 259.2276, 
    259.2281, 259.2278, 259.2281, 259.2278, 259.2276, 259.2295, 259.2284, 
    259.23, 259.2299, 259.2292, 259.2299, 259.223, 259.2228, 259.2221, 
    259.2227, 259.2217, 259.2222, 259.2225, 259.2237, 259.224, 259.2242, 
    259.2247, 259.2253, 259.2264, 259.2274, 259.2283, 259.2282, 259.2283, 
    259.2285, 259.228, 259.2285, 259.2286, 259.2284, 259.2299, 259.2295, 
    259.2299, 259.2296, 259.2229, 259.2232, 259.223, 259.2233, 259.2231, 
    259.2241, 259.2245, 259.2259, 259.2253, 259.2263, 259.2254, 259.2256, 
    259.2263, 259.2255, 259.2274, 259.226, 259.2285, 259.2271, 259.2286, 
    259.2283, 259.2287, 259.2291, 259.2296, 259.2305, 259.2303, 259.231, 
    259.2237, 259.2241, 259.2241, 259.2245, 259.2248, 259.2256, 259.2267, 
    259.2263, 259.2271, 259.2273, 259.226, 259.2268, 259.2244, 259.2248, 
    259.2245, 259.2237, 259.2264, 259.225, 259.2276, 259.2268, 259.229, 
    259.2279, 259.2301, 259.2311, 259.232, 259.2331, 259.2243, 259.2241, 
    259.2246, 259.2253, 259.226, 259.2269, 259.227, 259.2271, 259.2276, 
    259.2279, 259.2272, 259.228, 259.2248, 259.2265, 259.2239, 259.2247, 
    259.2252, 259.225, 259.2262, 259.2265, 259.2277, 259.2271, 259.2308, 
    259.2292, 259.2339, 259.2326, 259.2239, 259.2243, 259.2257, 259.225, 
    259.2269, 259.2274, 259.2278, 259.2282, 259.2283, 259.2286, 259.2281, 
    259.2286, 259.2269, 259.2276, 259.2256, 259.226, 259.2258, 259.2256, 
    259.2263, 259.2272, 259.2272, 259.2275, 259.2282, 259.2269, 259.231, 
    259.2285, 259.2248, 259.2255, 259.2256, 259.2253, 259.2273, 259.2266, 
    259.2286, 259.2281, 259.2289, 259.2285, 259.2284, 259.2279, 259.2275, 
    259.2266, 259.2259, 259.2254, 259.2255, 259.2261, 259.2272, 259.2283, 
    259.2281, 259.2289, 259.2268, 259.2277, 259.2273, 259.2282, 259.2263, 
    259.2278, 259.2259, 259.226, 259.2266, 259.2277, 259.228, 259.2282, 
    259.2281, 259.2273, 259.2271, 259.2266, 259.2264, 259.226, 259.2256, 
    259.226, 259.2263, 259.2273, 259.2281, 259.2291, 259.2293, 259.2304, 
    259.2295, 259.231, 259.2297, 259.232, 259.228, 259.2297, 259.2266, 
    259.227, 259.2275, 259.2289, 259.2282, 259.2291, 259.2271, 259.2261, 
    259.2259, 259.2254, 259.2259, 259.2259, 259.2263, 259.2262, 259.2273, 
    259.2267, 259.2284, 259.2291, 259.2309, 259.2321, 259.2332, 259.2338, 
    259.2339, 259.234,
  261.4064, 261.4069, 261.4068, 261.4071, 261.407, 261.4072, 261.4065, 
    261.4069, 261.4066, 261.4065, 261.4078, 261.4072, 261.4086, 261.4081, 
    261.4094, 261.4085, 261.4095, 261.4093, 261.4099, 261.4097, 261.4105, 
    261.41, 261.4109, 261.4104, 261.4104, 261.41, 261.4073, 261.4077, 
    261.4073, 261.4073, 261.4073, 261.407, 261.4067, 261.4064, 261.4065, 
    261.4067, 261.4073, 261.4071, 261.4077, 261.4077, 261.4083, 261.4081, 
    261.4091, 261.4088, 261.4098, 261.4095, 261.4097, 261.4097, 261.4097, 
    261.4094, 261.4095, 261.4092, 261.4081, 261.4084, 261.4074, 261.4069, 
    261.4065, 261.4063, 261.4063, 261.4064, 261.4067, 261.4071, 261.4073, 
    261.4075, 261.4077, 261.4082, 261.4085, 261.4092, 261.4091, 261.4093, 
    261.4095, 261.4098, 261.4098, 261.4099, 261.4093, 261.4097, 261.409, 
    261.4092, 261.4077, 261.4072, 261.407, 261.4068, 261.4063, 261.4066, 
    261.4065, 261.4068, 261.407, 261.4069, 261.4075, 261.4073, 261.4085, 
    261.408, 261.4095, 261.4091, 261.4095, 261.4093, 261.4097, 261.4094, 
    261.41, 261.4101, 261.41, 261.4104, 261.4093, 261.4097, 261.4069, 
    261.4069, 261.407, 261.4067, 261.4067, 261.4064, 261.4066, 261.4067, 
    261.407, 261.4072, 261.4073, 261.4077, 261.4081, 261.4087, 261.4091, 
    261.4094, 261.4092, 261.4094, 261.4092, 261.4091, 261.4101, 261.4095, 
    261.4103, 261.4103, 261.4099, 261.4103, 261.407, 261.4069, 261.4066, 
    261.4068, 261.4063, 261.4066, 261.4067, 261.4073, 261.4074, 261.4075, 
    261.4077, 261.4081, 261.4086, 261.4091, 261.4095, 261.4095, 261.4095, 
    261.4096, 261.4093, 261.4096, 261.4097, 261.4095, 261.4103, 261.4101, 
    261.4103, 261.4102, 261.4069, 261.407, 261.407, 261.4071, 261.407, 
    261.4075, 261.4076, 261.4083, 261.4081, 261.4085, 261.4081, 261.4082, 
    261.4085, 261.4081, 261.409, 261.4084, 261.4096, 261.4089, 261.4096, 
    261.4095, 261.4097, 261.4099, 261.4101, 261.4106, 261.4105, 261.4108, 
    261.4073, 261.4075, 261.4074, 261.4077, 261.4078, 261.4082, 261.4087, 
    261.4085, 261.4089, 261.409, 261.4084, 261.4088, 261.4076, 261.4078, 
    261.4077, 261.4073, 261.4085, 261.4079, 261.4091, 261.4088, 261.4099, 
    261.4093, 261.4104, 261.4109, 261.4113, 261.4119, 261.4076, 261.4074, 
    261.4077, 261.408, 261.4084, 261.4088, 261.4088, 261.4089, 261.4091, 
    261.4093, 261.4089, 261.4094, 261.4078, 261.4086, 261.4074, 261.4077, 
    261.408, 261.4079, 261.4085, 261.4086, 261.4092, 261.4089, 261.4108, 
    261.4099, 261.4123, 261.4116, 261.4074, 261.4076, 261.4082, 261.4079, 
    261.4088, 261.4091, 261.4092, 261.4095, 261.4095, 261.4096, 261.4094, 
    261.4096, 261.4088, 261.4091, 261.4081, 261.4084, 261.4083, 261.4082, 
    261.4085, 261.4089, 261.409, 261.4091, 261.4094, 261.4088, 261.4109, 
    261.4096, 261.4078, 261.4081, 261.4082, 261.4081, 261.409, 261.4087, 
    261.4096, 261.4094, 261.4098, 261.4096, 261.4095, 261.4093, 261.4091, 
    261.4087, 261.4083, 261.4081, 261.4081, 261.4084, 261.409, 261.4095, 
    261.4094, 261.4098, 261.4088, 261.4092, 261.409, 261.4095, 261.4085, 
    261.4093, 261.4083, 261.4084, 261.4087, 261.4092, 261.4093, 261.4095, 
    261.4094, 261.409, 261.4089, 261.4087, 261.4086, 261.4084, 261.4082, 
    261.4084, 261.4085, 261.409, 261.4094, 261.4099, 261.41, 261.4106, 
    261.4101, 261.4109, 261.4102, 261.4113, 261.4093, 261.4102, 261.4087, 
    261.4088, 261.4091, 261.4098, 261.4095, 261.4099, 261.4089, 261.4084, 
    261.4083, 261.4081, 261.4083, 261.4083, 261.4085, 261.4084, 261.409, 
    261.4087, 261.4095, 261.4099, 261.4108, 261.4114, 261.412, 261.4122, 
    261.4123, 261.4124,
  262.7626, 262.7627, 262.7627, 262.7628, 262.7627, 262.7628, 262.7626, 
    262.7627, 262.7627, 262.7626, 262.7629, 262.7628, 262.7631, 262.763, 
    262.7633, 262.7631, 262.7633, 262.7633, 262.7635, 262.7634, 262.7636, 
    262.7635, 262.7637, 262.7635, 262.7636, 262.7635, 262.7628, 262.7629, 
    262.7628, 262.7628, 262.7628, 262.7627, 262.7627, 262.7626, 262.7626, 
    262.7627, 262.7628, 262.7628, 262.7629, 262.7629, 262.7631, 262.763, 
    262.7632, 262.7632, 262.7634, 262.7633, 262.7634, 262.7634, 262.7634, 
    262.7633, 262.7634, 262.7633, 262.763, 262.7631, 262.7628, 262.7627, 
    262.7626, 262.7626, 262.7626, 262.7626, 262.7627, 262.7628, 262.7628, 
    262.7629, 262.7629, 262.763, 262.7631, 262.7633, 262.7632, 262.7633, 
    262.7633, 262.7634, 262.7634, 262.7635, 262.7633, 262.7634, 262.7632, 
    262.7633, 262.7629, 262.7628, 262.7628, 262.7627, 262.7626, 262.7627, 
    262.7626, 262.7627, 262.7628, 262.7627, 262.7629, 262.7628, 262.7631, 
    262.763, 262.7633, 262.7632, 262.7634, 262.7633, 262.7634, 262.7633, 
    262.7635, 262.7635, 262.7635, 262.7635, 262.7633, 262.7634, 262.7627, 
    262.7627, 262.7628, 262.7627, 262.7627, 262.7626, 262.7627, 262.7627, 
    262.7628, 262.7628, 262.7628, 262.7629, 262.763, 262.7632, 262.7632, 
    262.7633, 262.7633, 262.7633, 262.7633, 262.7632, 262.7635, 262.7634, 
    262.7635, 262.7635, 262.7635, 262.7635, 262.7627, 262.7627, 262.7626, 
    262.7627, 262.7626, 262.7627, 262.7627, 262.7628, 262.7628, 262.7629, 
    262.7629, 262.763, 262.7631, 262.7632, 262.7633, 262.7633, 262.7633, 
    262.7634, 262.7633, 262.7634, 262.7634, 262.7634, 262.7635, 262.7635, 
    262.7635, 262.7635, 262.7627, 262.7628, 262.7627, 262.7628, 262.7628, 
    262.7628, 262.7629, 262.7631, 262.763, 262.7631, 262.763, 262.763, 
    262.7631, 262.763, 262.7632, 262.7631, 262.7634, 262.7632, 262.7634, 
    262.7633, 262.7634, 262.7634, 262.7635, 262.7636, 262.7636, 262.7637, 
    262.7628, 262.7628, 262.7628, 262.7629, 262.7629, 262.763, 262.7632, 
    262.7631, 262.7632, 262.7632, 262.7631, 262.7632, 262.7629, 262.7629, 
    262.7629, 262.7628, 262.7631, 262.763, 262.7632, 262.7632, 262.7634, 
    262.7633, 262.7636, 262.7637, 262.7638, 262.7639, 262.7629, 262.7628, 
    262.7629, 262.763, 262.7631, 262.7632, 262.7632, 262.7632, 262.7632, 
    262.7633, 262.7632, 262.7633, 262.7629, 262.7631, 262.7628, 262.7629, 
    262.763, 262.763, 262.7631, 262.7631, 262.7633, 262.7632, 262.7637, 
    262.7635, 262.7641, 262.7639, 262.7628, 262.7629, 262.763, 262.763, 
    262.7632, 262.7632, 262.7633, 262.7633, 262.7633, 262.7634, 262.7633, 
    262.7634, 262.7632, 262.7633, 262.763, 262.7631, 262.7631, 262.763, 
    262.7631, 262.7632, 262.7632, 262.7632, 262.7633, 262.7632, 262.7637, 
    262.7634, 262.7629, 262.763, 262.763, 262.763, 262.7632, 262.7632, 
    262.7634, 262.7633, 262.7634, 262.7634, 262.7634, 262.7633, 262.7632, 
    262.7632, 262.7631, 262.763, 262.763, 262.7631, 262.7632, 262.7633, 
    262.7633, 262.7634, 262.7632, 262.7633, 262.7632, 262.7633, 262.7631, 
    262.7633, 262.7631, 262.7631, 262.7632, 262.7633, 262.7633, 262.7633, 
    262.7633, 262.7632, 262.7632, 262.7631, 262.7631, 262.7631, 262.763, 
    262.7631, 262.7631, 262.7632, 262.7633, 262.7634, 262.7635, 262.7636, 
    262.7635, 262.7637, 262.7635, 262.7638, 262.7633, 262.7635, 262.7632, 
    262.7632, 262.7632, 262.7634, 262.7633, 262.7634, 262.7632, 262.7631, 
    262.7631, 262.763, 262.7631, 262.7631, 262.7631, 262.7631, 262.7632, 
    262.7632, 262.7634, 262.7634, 262.7637, 262.7638, 262.764, 262.764, 
    262.7641, 262.7641,
  263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1177, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 
    263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1179, 263.1179, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1177, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1179, 263.1179, 263.1177, 263.1177, 263.1178, 263.1177, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1177, 263.1178, 263.1178, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1179, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1179, 263.1179, 263.1179, 
    263.1179, 263.1179,
  263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.1117, 263.1257, 263.123, 263.1342, 263.128, 263.1353, 263.1145, 
    263.1263, 263.1188, 263.113, 263.1557, 263.1347, 263.1775, 263.1642, 
    263.1977, 263.1754, 263.2021, 263.197, 263.2124, 263.208, 263.2276, 
    263.2145, 263.2378, 263.2245, 263.2266, 263.214, 263.1389, 263.1531, 
    263.1381, 263.1401, 263.1392, 263.1281, 263.1225, 263.1106, 263.1128, 
    263.1215, 263.141, 263.1345, 263.151, 263.1507, 263.1691, 263.1608, 
    263.1917, 263.1829, 263.2082, 263.2018, 263.2079, 263.2061, 263.2079, 
    263.1986, 263.2026, 263.1944, 263.1623, 263.1718, 263.1436, 263.1265, 
    263.1151, 263.1069, 263.1081, 263.1103, 263.1216, 263.1321, 263.1401, 
    263.1454, 263.1506, 263.1664, 263.1747, 263.1934, 263.1901, 263.1958, 
    263.2012, 263.2104, 263.2088, 263.2129, 263.1956, 263.2071, 263.1882, 
    263.1933, 263.152, 263.1362, 263.1295, 263.1235, 263.1089, 263.119, 
    263.1151, 263.1245, 263.1305, 263.1275, 263.1455, 263.1385, 263.1752, 
    263.1595, 263.2006, 263.1908, 263.2029, 263.1967, 263.2074, 263.1978, 
    263.2144, 263.218, 263.2155, 263.2249, 263.1973, 263.2079, 263.1274, 
    263.1279, 263.1302, 263.1203, 263.1197, 263.1106, 263.1187, 263.1221, 
    263.1308, 263.1359, 263.1407, 263.1513, 263.1631, 263.1796, 263.1914, 
    263.1993, 263.1945, 263.1988, 263.194, 263.1917, 263.2166, 263.2026, 
    263.2236, 263.2224, 263.213, 263.2226, 263.1283, 263.1255, 263.1158, 
    263.1234, 263.1096, 263.1173, 263.1217, 263.1387, 263.1424, 263.1458, 
    263.1526, 263.1612, 263.1764, 263.1895, 263.2015, 263.2007, 263.201, 
    263.2036, 263.197, 263.2047, 263.206, 263.2026, 263.2223, 263.2167, 
    263.2224, 263.2188, 263.1264, 263.131, 263.1285, 263.1332, 263.1299, 
    263.1446, 263.1489, 263.1694, 263.161, 263.1744, 263.1624, 263.1645, 
    263.1748, 263.1631, 263.1888, 263.1713, 263.2037, 263.1863, 263.2048, 
    263.2015, 263.207, 263.212, 263.2183, 263.2297, 263.2271, 263.2367, 
    263.1379, 263.1439, 263.1433, 263.1496, 263.1542, 263.1642, 263.1801, 
    263.1741, 263.1852, 263.1873, 263.1706, 263.1809, 263.1478, 263.1532, 
    263.15, 263.1384, 263.1755, 263.1565, 263.1916, 263.1813, 263.2113, 
    263.1964, 263.2256, 263.238, 263.2497, 263.2633, 263.1471, 263.1431, 
    263.1503, 263.1603, 263.1696, 263.1819, 263.1832, 263.1855, 263.1915, 
    263.1965, 263.1862, 263.1978, 263.1544, 263.1772, 263.1415, 263.1523, 
    263.1597, 263.1565, 263.1734, 263.1774, 263.1936, 263.1853, 263.2349, 
    263.213, 263.2737, 263.2568, 263.1417, 263.1471, 263.166, 263.157, 
    263.1828, 263.1891, 263.1942, 263.2008, 263.2015, 263.2054, 263.199, 
    263.2051, 263.1819, 263.1923, 263.1639, 263.1708, 263.1676, 263.1641, 
    263.1749, 263.1864, 263.1866, 263.1903, 263.2006, 263.1829, 263.2377, 
    263.2039, 263.153, 263.1635, 263.165, 263.1609, 263.1884, 263.1785, 
    263.2053, 263.198, 263.2099, 263.204, 263.2031, 263.1956, 263.1909, 
    263.179, 263.1693, 263.1616, 263.1633, 263.1718, 263.1871, 263.2015, 
    263.1984, 263.209, 263.1809, 263.1927, 263.1881, 263.2, 263.174, 
    263.1961, 263.1683, 263.1707, 263.1783, 263.1935, 263.1968, 263.2004, 
    263.1982, 263.1875, 263.1857, 263.1781, 263.176, 263.1702, 263.1654, 
    263.1698, 263.1744, 263.1875, 263.1992, 263.2121, 263.2152, 263.2301, 
    263.218, 263.2379, 263.2209, 263.2503, 263.1974, 263.2204, 263.1786, 
    263.1832, 263.1913, 263.21, 263.2, 263.2117, 263.1856, 263.1721, 
    263.1686, 263.162, 263.1687, 263.1682, 263.1746, 263.1725, 263.1879, 
    263.1797, 263.2031, 263.2116, 263.2357, 263.2503, 263.2652, 263.2718, 
    263.2738, 263.2747 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9051, 253.9059, 253.9058, 253.9064, 253.9061, 253.9065, 253.9053, 
    253.906, 253.9055, 253.9052, 253.9077, 253.9065, 253.9091, 253.9083, 
    253.9104, 253.909, 253.9107, 253.9104, 253.9113, 253.911, 253.9122, 
    253.9115, 253.9129, 253.9121, 253.9122, 253.9114, 253.9067, 253.9076, 
    253.9067, 253.9068, 253.9068, 253.9061, 253.9057, 253.905, 253.9052, 
    253.9057, 253.9069, 253.9065, 253.9075, 253.9075, 253.9086, 253.9081, 
    253.91, 253.9095, 253.9111, 253.9107, 253.911, 253.9109, 253.911, 
    253.9104, 253.9107, 253.9102, 253.9082, 253.9088, 253.907, 253.906, 
    253.9053, 253.9048, 253.9049, 253.905, 253.9057, 253.9063, 253.9068, 
    253.9072, 253.9075, 253.9084, 253.909, 253.9101, 253.9099, 253.9103, 
    253.9106, 253.9112, 253.9111, 253.9113, 253.9103, 253.911, 253.9098, 
    253.9101, 253.9075, 253.9066, 253.9061, 253.9058, 253.9049, 253.9055, 
    253.9053, 253.9059, 253.9062, 253.9061, 253.9072, 253.9067, 253.909, 
    253.908, 253.9106, 253.91, 253.9107, 253.9103, 253.911, 253.9104, 
    253.9114, 253.9117, 253.9115, 253.9121, 253.9104, 253.911, 253.906, 
    253.9061, 253.9062, 253.9056, 253.9056, 253.905, 253.9055, 253.9057, 
    253.9062, 253.9066, 253.9069, 253.9075, 253.9082, 253.9093, 253.91, 
    253.9105, 253.9102, 253.9105, 253.9102, 253.91, 253.9116, 253.9107, 
    253.912, 253.9119, 253.9113, 253.912, 253.9061, 253.9059, 253.9053, 
    253.9058, 253.905, 253.9054, 253.9057, 253.9067, 253.907, 253.9072, 
    253.9076, 253.9081, 253.9091, 253.9099, 253.9106, 253.9106, 253.9106, 
    253.9108, 253.9104, 253.9108, 253.9109, 253.9107, 253.9119, 253.9116, 
    253.9119, 253.9117, 253.906, 253.9063, 253.9061, 253.9064, 253.9062, 
    253.9071, 253.9073, 253.9086, 253.9081, 253.9089, 253.9082, 253.9083, 
    253.9089, 253.9082, 253.9098, 253.9087, 253.9108, 253.9097, 253.9108, 
    253.9106, 253.911, 253.9113, 253.9117, 253.9124, 253.9122, 253.9128, 
    253.9067, 253.907, 253.907, 253.9074, 253.9077, 253.9083, 253.9093, 
    253.9089, 253.9096, 253.9097, 253.9087, 253.9093, 253.9073, 253.9076, 
    253.9074, 253.9067, 253.909, 253.9078, 253.91, 253.9094, 253.9112, 
    253.9103, 253.9121, 253.9129, 253.9137, 253.9145, 253.9072, 253.907, 
    253.9075, 253.9081, 253.9086, 253.9094, 253.9095, 253.9096, 253.91, 
    253.9103, 253.9097, 253.9104, 253.9077, 253.9091, 253.9069, 253.9075, 
    253.908, 253.9078, 253.9089, 253.9091, 253.9101, 253.9096, 253.9127, 
    253.9113, 253.9152, 253.9141, 253.9069, 253.9073, 253.9084, 253.9079, 
    253.9095, 253.9099, 253.9102, 253.9106, 253.9106, 253.9109, 253.9105, 
    253.9109, 253.9094, 253.9101, 253.9083, 253.9087, 253.9085, 253.9083, 
    253.909, 253.9097, 253.9097, 253.9099, 253.9105, 253.9095, 253.9129, 
    253.9107, 253.9076, 253.9082, 253.9084, 253.9081, 253.9098, 253.9092, 
    253.9109, 253.9104, 253.9112, 253.9108, 253.9107, 253.9103, 253.91, 
    253.9092, 253.9086, 253.9081, 253.9083, 253.9088, 253.9097, 253.9106, 
    253.9104, 253.9111, 253.9093, 253.9101, 253.9098, 253.9105, 253.9089, 
    253.9102, 253.9086, 253.9087, 253.9092, 253.9101, 253.9103, 253.9106, 
    253.9104, 253.9097, 253.9096, 253.9092, 253.909, 253.9087, 253.9084, 
    253.9087, 253.9089, 253.9098, 253.9105, 253.9113, 253.9115, 253.9124, 
    253.9116, 253.9129, 253.9118, 253.9137, 253.9103, 253.9118, 253.9092, 
    253.9095, 253.91, 253.9111, 253.9105, 253.9113, 253.9096, 253.9088, 
    253.9086, 253.9082, 253.9086, 253.9086, 253.909, 253.9088, 253.9098, 
    253.9093, 253.9107, 253.9113, 253.9128, 253.9137, 253.9147, 253.9151, 
    253.9152, 253.9153 ;

 TWS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 T_SCALAR =
  0.1400014, 0.1400093, 0.1400078, 0.1400141, 0.1400107, 0.1400147, 
    0.1400031, 0.1400096, 0.1400055, 0.1400022, 0.1400261, 0.1400144, 
    0.140039, 0.1400314, 0.1400508, 0.1400377, 0.1400534, 0.1400505, 
    0.1400596, 0.140057, 0.1400684, 0.1400608, 0.1400745, 0.1400666, 
    0.1400678, 0.1400606, 0.1400169, 0.1400246, 0.1400164, 0.1400175, 
    0.140017, 0.1400107, 0.1400074, 0.1400009, 0.1400021, 0.1400069, 
    0.140018, 0.1400143, 0.1400239, 0.1400237, 0.1400342, 0.1400295, 
    0.1400474, 0.1400423, 0.1400571, 0.1400534, 0.1400569, 0.1400559, 
    0.140057, 0.1400515, 0.1400538, 0.140049, 0.1400303, 0.1400357, 
    0.1400195, 0.1400095, 0.1400033, 0.1399988, 0.1399995, 0.1400006, 
    0.1400069, 0.140013, 0.1400176, 0.1400206, 0.1400236, 0.1400324, 
    0.1400374, 0.1400483, 0.1400465, 0.1400497, 0.140053, 0.1400584, 
    0.1400575, 0.1400598, 0.1400497, 0.1400564, 0.1400454, 0.1400484, 
    0.1400239, 0.1400153, 0.1400112, 0.1400081, 0.1399999, 0.1400055, 
    0.1400033, 0.1400087, 0.140012, 0.1400104, 0.1400207, 0.1400167, 
    0.1400377, 0.1400286, 0.1400526, 0.1400469, 0.140054, 0.1400504, 
    0.1400566, 0.140051, 0.1400607, 0.1400628, 0.1400614, 0.140067, 
    0.1400507, 0.1400569, 0.1400103, 0.1400106, 0.1400119, 0.1400062, 
    0.1400059, 0.1400009, 0.1400054, 0.1400073, 0.1400123, 0.1400151, 
    0.1400179, 0.140024, 0.1400307, 0.1400403, 0.1400473, 0.1400519, 
    0.1400491, 0.1400516, 0.1400488, 0.1400475, 0.140062, 0.1400538, 
    0.1400662, 0.1400655, 0.1400599, 0.1400656, 0.1400108, 0.1400093, 
    0.1400038, 0.1400081, 0.1400003, 0.1400046, 0.140007, 0.1400166, 
    0.1400189, 0.1400208, 0.1400247, 0.1400297, 0.1400384, 0.1400461, 
    0.1400532, 0.1400527, 0.1400529, 0.1400544, 0.1400505, 0.1400551, 
    0.1400558, 0.1400539, 0.1400654, 0.1400621, 0.1400655, 0.1400634, 
    0.1400098, 0.1400124, 0.140011, 0.1400136, 0.1400117, 0.14002, 0.1400225, 
    0.1400343, 0.1400296, 0.1400373, 0.1400304, 0.1400316, 0.1400373, 
    0.1400308, 0.1400456, 0.1400353, 0.1400545, 0.140044, 0.1400551, 
    0.1400532, 0.1400565, 0.1400593, 0.140063, 0.1400697, 0.1400682, 
    0.1400739, 0.1400163, 0.1400196, 0.1400194, 0.140023, 0.1400256, 
    0.1400314, 0.1400407, 0.1400372, 0.1400436, 0.1400449, 0.1400352, 
    0.1400411, 0.140022, 0.1400249, 0.1400232, 0.1400165, 0.1400379, 
    0.1400268, 0.1400474, 0.1400414, 0.1400589, 0.1400501, 0.1400673, 
    0.1400745, 0.1400817, 0.1400897, 0.1400216, 0.1400193, 0.1400235, 
    0.1400291, 0.1400346, 0.1400417, 0.1400425, 0.1400438, 0.1400473, 
    0.1400503, 0.1400441, 0.140051, 0.1400254, 0.1400389, 0.1400183, 
    0.1400244, 0.1400288, 0.1400269, 0.1400369, 0.1400391, 0.1400485, 
    0.1400437, 0.1400726, 0.1400598, 0.1400961, 0.1400858, 0.1400185, 
    0.1400216, 0.1400324, 0.1400273, 0.1400422, 0.1400459, 0.140049, 
    0.1400527, 0.1400532, 0.1400554, 0.1400517, 0.1400553, 0.1400417, 
    0.1400478, 0.1400313, 0.1400352, 0.1400335, 0.1400314, 0.1400377, 
    0.1400442, 0.1400445, 0.1400466, 0.1400521, 0.1400423, 0.140074, 
    0.1400541, 0.140025, 0.1400309, 0.1400319, 0.1400296, 0.1400455, 
    0.1400397, 0.1400554, 0.1400512, 0.1400581, 0.1400547, 0.1400541, 
    0.1400497, 0.1400469, 0.14004, 0.1400343, 0.14003, 0.140031, 0.1400358, 
    0.1400446, 0.1400532, 0.1400513, 0.1400576, 0.1400411, 0.1400479, 
    0.1400453, 0.1400523, 0.1400371, 0.1400495, 0.1400339, 0.1400353, 
    0.1400396, 0.1400483, 0.1400505, 0.1400525, 0.1400513, 0.1400449, 
    0.1400439, 0.1400395, 0.1400383, 0.140035, 0.1400322, 0.1400347, 
    0.1400373, 0.140045, 0.1400518, 0.1400593, 0.1400613, 0.1400697, 
    0.1400626, 0.1400741, 0.140064, 0.1400817, 0.1400505, 0.140064, 
    0.1400399, 0.1400425, 0.1400471, 0.140058, 0.1400523, 0.140059, 
    0.1400439, 0.1400359, 0.140034, 0.1400302, 0.1400341, 0.1400338, 
    0.1400375, 0.1400363, 0.1400452, 0.1400404, 0.1400541, 0.140059, 
    0.1400733, 0.1400819, 0.140091, 0.140095, 0.1400962, 0.1400967,
  0.1463853, 0.146394, 0.1463923, 0.1463993, 0.1463955, 0.1464, 0.1463871, 
    0.1463943, 0.1463897, 0.1463861, 0.1464126, 0.1463996, 0.1464269, 
    0.1464184, 0.14644, 0.1464255, 0.146443, 0.1464398, 0.1464499, 0.146447, 
    0.1464596, 0.1464512, 0.1464665, 0.1464577, 0.146459, 0.1464509, 
    0.1464024, 0.1464109, 0.1464018, 0.1464031, 0.1464025, 0.1463955, 
    0.1463918, 0.1463847, 0.146386, 0.1463913, 0.1464036, 0.1463995, 
    0.1464101, 0.1464099, 0.1464216, 0.1464163, 0.1464363, 0.1464306, 
    0.1464471, 0.1464429, 0.1464469, 0.1464457, 0.1464469, 0.1464408, 
    0.1464434, 0.146438, 0.1464173, 0.1464233, 0.1464053, 0.1463943, 
    0.1463874, 0.1463824, 0.1463831, 0.1463844, 0.1463914, 0.1463981, 
    0.1464031, 0.1464065, 0.1464099, 0.1464196, 0.1464251, 0.1464373, 
    0.1464353, 0.1464389, 0.1464425, 0.1464485, 0.1464475, 0.1464501, 
    0.1464389, 0.1464463, 0.1464341, 0.1464374, 0.1464102, 0.1464007, 
    0.1463961, 0.1463926, 0.1463836, 0.1463898, 0.1463874, 0.1463933, 
    0.146397, 0.1463952, 0.1464066, 0.1464021, 0.1464255, 0.1464154, 
    0.1464421, 0.1464357, 0.1464436, 0.1464396, 0.1464465, 0.1464403, 
    0.1464511, 0.1464534, 0.1464518, 0.1464581, 0.1464399, 0.1464468, 
    0.1463951, 0.1463954, 0.1463968, 0.1463906, 0.1463902, 0.1463846, 
    0.1463896, 0.1463917, 0.1463973, 0.1464004, 0.1464035, 0.1464102, 
    0.1464177, 0.1464283, 0.1464361, 0.1464413, 0.1464381, 0.1464409, 
    0.1464378, 0.1464364, 0.1464525, 0.1464434, 0.1464572, 0.1464564, 
    0.1464501, 0.1464565, 0.1463956, 0.1463939, 0.1463879, 0.1463926, 
    0.146384, 0.1463888, 0.1463914, 0.1464021, 0.1464046, 0.1464067, 
    0.1464111, 0.1464166, 0.1464263, 0.1464348, 0.1464427, 0.1464422, 
    0.1464424, 0.1464441, 0.1464398, 0.1464448, 0.1464456, 0.1464434, 
    0.1464563, 0.1464527, 0.1464564, 0.146454, 0.1463945, 0.1463974, 
    0.1463958, 0.1463987, 0.1463966, 0.1464058, 0.1464086, 0.1464217, 
    0.1464165, 0.146425, 0.1464174, 0.1464187, 0.146425, 0.1464178, 
    0.1464342, 0.1464229, 0.1464442, 0.1464325, 0.1464449, 0.1464427, 
    0.1464463, 0.1464495, 0.1464537, 0.1464612, 0.1464594, 0.1464658, 
    0.1464017, 0.1464054, 0.1464052, 0.1464092, 0.1464121, 0.1464185, 
    0.1464288, 0.1464249, 0.1464321, 0.1464335, 0.1464227, 0.1464292, 
    0.146408, 0.1464113, 0.1464094, 0.146402, 0.1464257, 0.1464134, 
    0.1464362, 0.1464295, 0.1464491, 0.1464392, 0.1464585, 0.1464665, 
    0.1464746, 0.1464834, 0.1464076, 0.146405, 0.1464097, 0.1464159, 
    0.146422, 0.1464299, 0.1464308, 0.1464323, 0.1464362, 0.1464394, 
    0.1464326, 0.1464403, 0.1464119, 0.1464268, 0.146404, 0.1464107, 
    0.1464156, 0.1464135, 0.1464245, 0.1464271, 0.1464375, 0.1464322, 
    0.1464644, 0.1464501, 0.1464906, 0.1464791, 0.1464041, 0.1464076, 
    0.1464196, 0.1464139, 0.1464305, 0.1464346, 0.146438, 0.1464422, 
    0.1464427, 0.1464452, 0.1464411, 0.1464451, 0.1464299, 0.1464367, 
    0.1464184, 0.1464227, 0.1464208, 0.1464185, 0.1464255, 0.1464327, 
    0.146433, 0.1464353, 0.1464415, 0.1464306, 0.146466, 0.1464438, 
    0.1464114, 0.1464179, 0.146419, 0.1464165, 0.1464342, 0.1464277, 
    0.1464451, 0.1464405, 0.1464482, 0.1464443, 0.1464438, 0.1464389, 
    0.1464358, 0.146428, 0.1464217, 0.1464169, 0.146418, 0.1464234, 
    0.1464332, 0.1464427, 0.1464406, 0.1464476, 0.1464293, 0.1464369, 
    0.1464339, 0.1464417, 0.1464248, 0.1464387, 0.1464212, 0.1464228, 
    0.1464276, 0.1464373, 0.1464397, 0.1464419, 0.1464406, 0.1464335, 
    0.1464324, 0.1464275, 0.1464261, 0.1464224, 0.1464193, 0.1464221, 
    0.146425, 0.1464335, 0.1464412, 0.1464496, 0.1464517, 0.1464611, 
    0.1464532, 0.1464661, 0.1464548, 0.1464745, 0.1464397, 0.1464548, 
    0.1464279, 0.1464308, 0.1464359, 0.1464481, 0.1464417, 0.1464492, 
    0.1464324, 0.1464235, 0.1464214, 0.1464171, 0.1464215, 0.1464211, 
    0.1464253, 0.1464239, 0.1464338, 0.1464285, 0.1464437, 0.1464492, 
    0.1464651, 0.1464748, 0.146485, 0.1464894, 0.1464907, 0.1464913,
  0.1561714, 0.1561798, 0.1561782, 0.1561849, 0.1561813, 0.1561856, 
    0.1561732, 0.1561801, 0.1561757, 0.1561723, 0.1561978, 0.1561852, 
    0.1562117, 0.1562034, 0.1562244, 0.1562103, 0.1562273, 0.1562242, 
    0.156234, 0.1562312, 0.1562436, 0.1562353, 0.1562503, 0.1562417, 
    0.156243, 0.1562351, 0.1561879, 0.1561962, 0.1561874, 0.1561886, 
    0.1561881, 0.1561813, 0.1561778, 0.1561709, 0.1561722, 0.1561773, 
    0.1561891, 0.1561852, 0.1561954, 0.1561952, 0.1562065, 0.1562014, 
    0.1562207, 0.1562153, 0.1562313, 0.1562272, 0.1562311, 0.15623, 
    0.1562311, 0.1562252, 0.1562277, 0.1562225, 0.1562023, 0.1562082, 
    0.1561907, 0.1561801, 0.1561735, 0.1561687, 0.1561694, 0.1561706, 
    0.1561773, 0.1561837, 0.1561886, 0.1561919, 0.1561951, 0.1562046, 
    0.15621, 0.1562218, 0.1562198, 0.1562233, 0.1562268, 0.1562327, 
    0.1562317, 0.1562342, 0.1562233, 0.1562305, 0.1562186, 0.1562218, 
    0.1561955, 0.1561863, 0.1561819, 0.1561785, 0.1561699, 0.1561758, 
    0.1561734, 0.1561792, 0.1561827, 0.156181, 0.156192, 0.1561877, 
    0.1562103, 0.1562005, 0.1562264, 0.1562202, 0.1562279, 0.156224, 
    0.1562307, 0.1562247, 0.1562352, 0.1562375, 0.1562359, 0.1562421, 
    0.1562243, 0.1562311, 0.1561809, 0.1561812, 0.1561826, 0.1561765, 
    0.1561762, 0.1561708, 0.1561756, 0.1561777, 0.156183, 0.156186, 0.156189, 
    0.1561955, 0.1562027, 0.156213, 0.1562206, 0.1562257, 0.1562226, 
    0.1562253, 0.1562223, 0.1562209, 0.1562366, 0.1562277, 0.1562412, 
    0.1562405, 0.1562343, 0.1562405, 0.1561814, 0.1561798, 0.1561739, 
    0.1561785, 0.1561703, 0.1561748, 0.1561774, 0.1561877, 0.1561901, 
    0.1561921, 0.1561963, 0.1562017, 0.156211, 0.1562194, 0.1562271, 
    0.1562265, 0.1562267, 0.1562284, 0.1562242, 0.1562291, 0.1562299, 
    0.1562278, 0.1562404, 0.1562368, 0.1562404, 0.1562381, 0.1561803, 
    0.1561831, 0.1561816, 0.1561844, 0.1561824, 0.1561912, 0.1561939, 
    0.1562066, 0.1562015, 0.1562098, 0.1562024, 0.1562037, 0.1562098, 
    0.1562028, 0.1562188, 0.1562078, 0.1562285, 0.1562171, 0.1562292, 
    0.156227, 0.1562306, 0.1562337, 0.1562378, 0.1562451, 0.1562434, 
    0.1562496, 0.1561873, 0.1561909, 0.1561906, 0.1561945, 0.1561973, 
    0.1562035, 0.1562135, 0.1562097, 0.1562167, 0.1562181, 0.1562076, 
    0.1562139, 0.1561933, 0.1561965, 0.1561947, 0.1561875, 0.1562105, 
    0.1561986, 0.1562207, 0.1562142, 0.1562333, 0.1562237, 0.1562425, 
    0.1562503, 0.1562582, 0.156267, 0.1561929, 0.1561905, 0.156195, 0.156201, 
    0.1562069, 0.1562146, 0.1562154, 0.1562169, 0.1562207, 0.1562239, 
    0.1562172, 0.1562247, 0.1561971, 0.1562115, 0.1561895, 0.1561959, 
    0.1562007, 0.1561987, 0.1562093, 0.1562118, 0.156222, 0.1562168, 
    0.1562483, 0.1562342, 0.156274, 0.1562627, 0.1561896, 0.156193, 
    0.1562046, 0.1561991, 0.1562152, 0.1562191, 0.1562224, 0.1562265, 
    0.156227, 0.1562295, 0.1562255, 0.1562293, 0.1562146, 0.1562212, 
    0.1562034, 0.1562076, 0.1562057, 0.1562035, 0.1562103, 0.1562173, 
    0.1562176, 0.1562199, 0.1562259, 0.1562152, 0.1562498, 0.1562281, 
    0.1561966, 0.1562029, 0.156204, 0.1562015, 0.1562187, 0.1562124, 
    0.1562294, 0.1562248, 0.1562324, 0.1562286, 0.1562281, 0.1562233, 
    0.1562203, 0.1562127, 0.1562066, 0.1562019, 0.156203, 0.1562082, 
    0.1562178, 0.156227, 0.156225, 0.1562318, 0.156214, 0.1562214, 0.1562185, 
    0.1562261, 0.1562096, 0.1562231, 0.1562061, 0.1562076, 0.1562123, 
    0.1562217, 0.1562241, 0.1562263, 0.156225, 0.1562181, 0.156217, 
    0.1562123, 0.1562109, 0.1562073, 0.1562043, 0.156207, 0.1562098, 
    0.1562181, 0.1562255, 0.1562337, 0.1562358, 0.1562451, 0.1562373, 
    0.1562499, 0.1562389, 0.1562582, 0.1562242, 0.1562389, 0.1562126, 
    0.1562154, 0.1562204, 0.1562323, 0.156226, 0.1562334, 0.156217, 
    0.1562083, 0.1562063, 0.1562022, 0.1562064, 0.156206, 0.1562101, 
    0.1562088, 0.1562184, 0.1562132, 0.156228, 0.1562334, 0.1562489, 
    0.1562584, 0.1562685, 0.1562728, 0.1562742, 0.1562747,
  0.1699164, 0.1699228, 0.1699216, 0.1699268, 0.1699239, 0.1699273, 
    0.1699177, 0.169923, 0.1699197, 0.169917, 0.1699368, 0.169927, 0.1699477, 
    0.1699412, 0.1699577, 0.1699466, 0.16996, 0.1699575, 0.1699654, 
    0.1699631, 0.169973, 0.1699664, 0.1699784, 0.1699715, 0.1699725, 
    0.1699662, 0.1699291, 0.1699356, 0.1699287, 0.1699296, 0.1699292, 
    0.169924, 0.1699212, 0.169916, 0.1699169, 0.1699209, 0.16993, 0.169927, 
    0.1699349, 0.1699348, 0.1699436, 0.1699396, 0.1699549, 0.1699505, 
    0.1699632, 0.16996, 0.1699631, 0.1699621, 0.1699631, 0.1699583, 
    0.1699603, 0.1699562, 0.1699404, 0.1699449, 0.1699313, 0.1699231, 
    0.1699179, 0.1699142, 0.1699148, 0.1699157, 0.1699209, 0.1699259, 
    0.1699297, 0.1699322, 0.1699347, 0.1699421, 0.1699463, 0.1699557, 
    0.1699541, 0.1699569, 0.1699597, 0.1699643, 0.1699635, 0.1699656, 
    0.1699569, 0.1699626, 0.1699532, 0.1699557, 0.169935, 0.1699278, 
    0.1699245, 0.1699218, 0.1699152, 0.1699197, 0.1699179, 0.1699223, 
    0.1699251, 0.1699237, 0.1699323, 0.1699289, 0.1699466, 0.1699389, 
    0.1699593, 0.1699544, 0.1699605, 0.1699574, 0.1699627, 0.169958, 
    0.1699663, 0.1699681, 0.1699669, 0.1699718, 0.1699577, 0.169963, 
    0.1699237, 0.1699239, 0.169925, 0.1699203, 0.16992, 0.1699159, 0.1699196, 
    0.1699212, 0.1699253, 0.1699277, 0.16993, 0.169935, 0.1699407, 0.1699488, 
    0.1699547, 0.1699587, 0.1699563, 0.1699584, 0.169956, 0.1699549, 
    0.1699674, 0.1699603, 0.1699711, 0.1699705, 0.1699656, 0.1699706, 
    0.1699241, 0.1699228, 0.1699183, 0.1699218, 0.1699155, 0.169919, 
    0.169921, 0.1699289, 0.1699308, 0.1699324, 0.1699356, 0.1699398, 
    0.1699472, 0.1699537, 0.1699599, 0.1699594, 0.1699596, 0.1699609, 
    0.1699575, 0.1699614, 0.1699621, 0.1699604, 0.1699704, 0.1699675, 
    0.1699705, 0.1699686, 0.1699232, 0.1699254, 0.1699242, 0.1699264, 
    0.1699248, 0.1699317, 0.1699338, 0.1699437, 0.1699397, 0.1699462, 
    0.1699404, 0.1699414, 0.1699463, 0.1699408, 0.1699533, 0.1699446, 
    0.1699609, 0.169952, 0.1699615, 0.1699598, 0.1699626, 0.1699651, 
    0.1699684, 0.1699742, 0.1699729, 0.1699778, 0.1699286, 0.1699314, 
    0.1699312, 0.1699342, 0.1699364, 0.1699413, 0.1699491, 0.1699462, 
    0.1699516, 0.1699527, 0.1699445, 0.1699494, 0.1699333, 0.1699358, 
    0.1699344, 0.1699288, 0.1699467, 0.1699374, 0.1699548, 0.1699497, 
    0.1699648, 0.1699571, 0.1699721, 0.1699784, 0.1699847, 0.1699918, 
    0.169933, 0.1699311, 0.1699346, 0.1699393, 0.1699439, 0.16995, 0.1699507, 
    0.1699518, 0.1699548, 0.1699573, 0.1699521, 0.1699579, 0.1699363, 
    0.1699476, 0.1699303, 0.1699354, 0.1699391, 0.1699375, 0.1699459, 
    0.1699478, 0.1699558, 0.1699517, 0.1699768, 0.1699656, 0.1699975, 
    0.1699884, 0.1699304, 0.169933, 0.1699421, 0.1699378, 0.1699504, 
    0.1699536, 0.1699562, 0.1699594, 0.1699598, 0.1699618, 0.1699586, 
    0.1699616, 0.16995, 0.1699552, 0.1699412, 0.1699445, 0.169943, 0.1699413, 
    0.1699466, 0.1699521, 0.1699524, 0.1699542, 0.1699589, 0.1699505, 
    0.169978, 0.1699607, 0.1699359, 0.1699408, 0.1699417, 0.1699397, 
    0.1699532, 0.1699483, 0.1699617, 0.1699581, 0.1699641, 0.1699611, 
    0.1699606, 0.1699568, 0.1699545, 0.1699485, 0.1699437, 0.16994, 
    0.1699409, 0.169945, 0.1699525, 0.1699598, 0.1699582, 0.1699636, 
    0.1699495, 0.1699553, 0.169953, 0.1699591, 0.1699461, 0.1699567, 
    0.1699433, 0.1699445, 0.1699482, 0.1699556, 0.1699575, 0.1699592, 
    0.1699582, 0.1699527, 0.1699519, 0.1699481, 0.1699471, 0.1699443, 
    0.1699419, 0.169944, 0.1699463, 0.1699528, 0.1699586, 0.1699651, 
    0.1699668, 0.1699742, 0.169968, 0.1699781, 0.1699693, 0.1699847, 
    0.1699575, 0.1699692, 0.1699484, 0.1699506, 0.1699546, 0.169964, 
    0.169959, 0.1699649, 0.1699519, 0.1699451, 0.1699435, 0.1699402, 
    0.1699435, 0.1699433, 0.1699464, 0.1699454, 0.169953, 0.1699489, 
    0.1699606, 0.1699649, 0.1699773, 0.1699849, 0.169993, 0.1699965, 
    0.1699976, 0.169998,
  0.1852159, 0.1852192, 0.1852185, 0.1852212, 0.1852197, 0.1852214, 
    0.1852166, 0.1852193, 0.1852176, 0.1852162, 0.1852263, 0.1852213, 
    0.185232, 0.1852286, 0.1852373, 0.1852314, 0.1852386, 0.1852372, 
    0.1852414, 0.1852402, 0.1852455, 0.185242, 0.1852484, 0.1852447, 
    0.1852453, 0.1852418, 0.1852224, 0.1852257, 0.1852222, 0.1852226, 
    0.1852224, 0.1852197, 0.1852183, 0.1852157, 0.1852162, 0.1852182, 
    0.1852228, 0.1852213, 0.1852254, 0.1852253, 0.1852299, 0.1852278, 
    0.1852358, 0.1852335, 0.1852403, 0.1852385, 0.1852402, 0.1852397, 
    0.1852402, 0.1852376, 0.1852387, 0.1852365, 0.1852282, 0.1852306, 
    0.1852235, 0.1852193, 0.1852167, 0.1852148, 0.1852151, 0.1852156, 
    0.1852182, 0.1852207, 0.1852227, 0.185224, 0.1852253, 0.1852291, 
    0.1852313, 0.1852362, 0.1852354, 0.1852369, 0.1852384, 0.1852408, 
    0.1852404, 0.1852415, 0.1852369, 0.1852399, 0.1852349, 0.1852362, 
    0.1852254, 0.1852217, 0.18522, 0.1852186, 0.1852153, 0.1852176, 
    0.1852167, 0.1852189, 0.1852203, 0.1852196, 0.185224, 0.1852223, 
    0.1852314, 0.1852274, 0.1852382, 0.1852356, 0.1852388, 0.1852372, 
    0.18524, 0.1852375, 0.1852419, 0.1852429, 0.1852422, 0.1852449, 
    0.1852373, 0.1852401, 0.1852196, 0.1852197, 0.1852202, 0.1852179, 
    0.1852177, 0.1852157, 0.1852175, 0.1852183, 0.1852204, 0.1852216, 
    0.1852228, 0.1852254, 0.1852283, 0.1852326, 0.1852357, 0.1852379, 
    0.1852366, 0.1852377, 0.1852364, 0.1852358, 0.1852425, 0.1852387, 
    0.1852445, 0.1852442, 0.1852415, 0.1852442, 0.1852198, 0.1852192, 
    0.1852169, 0.1852186, 0.1852154, 0.1852172, 0.1852182, 0.1852223, 
    0.1852232, 0.185224, 0.1852257, 0.1852279, 0.1852318, 0.1852352, 
    0.1852385, 0.1852382, 0.1852383, 0.185239, 0.1852372, 0.1852393, 
    0.1852396, 0.1852387, 0.1852441, 0.1852426, 0.1852442, 0.1852432, 
    0.1852194, 0.1852205, 0.1852199, 0.185221, 0.1852202, 0.1852237, 
    0.1852248, 0.1852299, 0.1852279, 0.1852312, 0.1852282, 0.1852287, 
    0.1852313, 0.1852284, 0.185235, 0.1852304, 0.185239, 0.1852343, 
    0.1852393, 0.1852384, 0.1852399, 0.1852413, 0.185243, 0.1852462, 
    0.1852455, 0.1852482, 0.1852221, 0.1852235, 0.1852235, 0.185225, 
    0.1852261, 0.1852287, 0.1852328, 0.1852312, 0.1852341, 0.1852347, 
    0.1852303, 0.1852329, 0.1852245, 0.1852258, 0.1852251, 0.1852222, 
    0.1852315, 0.1852267, 0.1852358, 0.1852331, 0.1852411, 0.185237, 
    0.185245, 0.1852485, 0.1852519, 0.1852558, 0.1852244, 0.1852234, 
    0.1852252, 0.1852276, 0.18523, 0.1852332, 0.1852336, 0.1852342, 
    0.1852358, 0.1852371, 0.1852343, 0.1852374, 0.1852261, 0.185232, 
    0.185223, 0.1852256, 0.1852275, 0.1852267, 0.1852311, 0.1852321, 
    0.1852363, 0.1852341, 0.1852476, 0.1852415, 0.185259, 0.1852539, 
    0.185223, 0.1852244, 0.1852291, 0.1852268, 0.1852335, 0.1852351, 
    0.1852365, 0.1852382, 0.1852384, 0.1852395, 0.1852378, 0.1852394, 
    0.1852332, 0.185236, 0.1852286, 0.1852303, 0.1852296, 0.1852287, 
    0.1852314, 0.1852344, 0.1852345, 0.1852354, 0.185238, 0.1852335, 
    0.1852482, 0.1852389, 0.1852259, 0.1852284, 0.1852289, 0.1852279, 
    0.1852349, 0.1852323, 0.1852394, 0.1852375, 0.1852407, 0.1852391, 
    0.1852389, 0.1852369, 0.1852356, 0.1852324, 0.1852299, 0.185228, 
    0.1852285, 0.1852306, 0.1852345, 0.1852384, 0.1852376, 0.1852405, 
    0.185233, 0.1852361, 0.1852348, 0.185238, 0.1852312, 0.1852368, 
    0.1852297, 0.1852303, 0.1852323, 0.1852362, 0.1852372, 0.1852381, 
    0.1852376, 0.1852347, 0.1852342, 0.1852323, 0.1852317, 0.1852302, 
    0.185229, 0.1852301, 0.1852313, 0.1852347, 0.1852378, 0.1852413, 
    0.1852422, 0.1852462, 0.1852428, 0.1852483, 0.1852435, 0.1852519, 
    0.1852372, 0.1852435, 0.1852324, 0.1852336, 0.1852357, 0.1852407, 
    0.185238, 0.1852411, 0.1852342, 0.1852306, 0.1852298, 0.1852281, 
    0.1852298, 0.1852297, 0.1852313, 0.1852308, 0.1852348, 0.1852327, 
    0.1852389, 0.1852411, 0.1852479, 0.185252, 0.1852565, 0.1852584, 
    0.185259, 0.1852593,
  0.1954502, 0.1954509, 0.1954508, 0.1954514, 0.1954511, 0.1954515, 
    0.1954503, 0.195451, 0.1954506, 0.1954502, 0.1954527, 0.1954515, 
    0.1954542, 0.1954533, 0.1954556, 0.195454, 0.1954559, 0.1954555, 
    0.1954566, 0.1954563, 0.1954578, 0.1954568, 0.1954586, 0.1954575, 
    0.1954577, 0.1954568, 0.1954517, 0.1954526, 0.1954517, 0.1954518, 
    0.1954518, 0.1954511, 0.1954508, 0.1954501, 0.1954502, 0.1954507, 
    0.1954519, 0.1954515, 0.1954525, 0.1954525, 0.1954536, 0.1954531, 
    0.1954551, 0.1954546, 0.1954563, 0.1954559, 0.1954563, 0.1954562, 
    0.1954563, 0.1954556, 0.1954559, 0.1954553, 0.1954532, 0.1954538, 
    0.195452, 0.195451, 0.1954504, 0.1954499, 0.19545, 0.1954501, 0.1954507, 
    0.1954513, 0.1954518, 0.1954521, 0.1954525, 0.1954534, 0.195454, 
    0.1954553, 0.195455, 0.1954554, 0.1954558, 0.1954565, 0.1954564, 
    0.1954567, 0.1954554, 0.1954562, 0.1954549, 0.1954553, 0.1954525, 
    0.1954516, 0.1954512, 0.1954508, 0.19545, 0.1954506, 0.1954504, 
    0.1954509, 0.1954512, 0.1954511, 0.1954521, 0.1954517, 0.195454, 
    0.195453, 0.1954558, 0.1954551, 0.195456, 0.1954555, 0.1954563, 
    0.1954556, 0.1954568, 0.195457, 0.1954569, 0.1954576, 0.1954556, 
    0.1954563, 0.1954511, 0.1954511, 0.1954512, 0.1954506, 0.1954506, 
    0.1954501, 0.1954506, 0.1954508, 0.1954513, 0.1954516, 0.1954518, 
    0.1954525, 0.1954532, 0.1954543, 0.1954551, 0.1954557, 0.1954554, 
    0.1954557, 0.1954553, 0.1954552, 0.1954569, 0.1954559, 0.1954575, 
    0.1954574, 0.1954567, 0.1954574, 0.1954511, 0.1954509, 0.1954504, 
    0.1954508, 0.1954501, 0.1954505, 0.1954507, 0.1954517, 0.1954519, 
    0.1954522, 0.1954526, 0.1954531, 0.1954541, 0.195455, 0.1954558, 
    0.1954558, 0.1954558, 0.195456, 0.1954555, 0.1954561, 0.1954562, 
    0.1954559, 0.1954574, 0.195457, 0.1954574, 0.1954571, 0.195451, 
    0.1954513, 0.1954511, 0.1954514, 0.1954512, 0.1954521, 0.1954523, 
    0.1954536, 0.1954531, 0.195454, 0.1954532, 0.1954533, 0.195454, 
    0.1954532, 0.1954549, 0.1954537, 0.195456, 0.1954547, 0.1954561, 
    0.1954558, 0.1954563, 0.1954566, 0.1954571, 0.1954579, 0.1954577, 
    0.1954585, 0.1954517, 0.195452, 0.195452, 0.1954524, 0.1954527, 
    0.1954533, 0.1954544, 0.195454, 0.1954547, 0.1954549, 0.1954537, 
    0.1954544, 0.1954523, 0.1954526, 0.1954524, 0.1954517, 0.195454, 
    0.1954528, 0.1954551, 0.1954544, 0.1954565, 0.1954555, 0.1954576, 
    0.1954586, 0.1954595, 0.1954606, 0.1954522, 0.195452, 0.1954524, 
    0.195453, 0.1954537, 0.1954545, 0.1954546, 0.1954547, 0.1954551, 
    0.1954555, 0.1954548, 0.1954556, 0.1954526, 0.1954542, 0.1954519, 
    0.1954525, 0.195453, 0.1954528, 0.1954539, 0.1954542, 0.1954553, 
    0.1954547, 0.1954583, 0.1954567, 0.1954615, 0.1954601, 0.1954519, 
    0.1954522, 0.1954534, 0.1954529, 0.1954545, 0.195455, 0.1954553, 
    0.1954558, 0.1954558, 0.1954561, 0.1954557, 0.1954561, 0.1954545, 
    0.1954552, 0.1954533, 0.1954537, 0.1954535, 0.1954533, 0.195454, 
    0.1954548, 0.1954548, 0.195455, 0.1954557, 0.1954546, 0.1954585, 
    0.195456, 0.1954526, 0.1954532, 0.1954534, 0.1954531, 0.1954549, 
    0.1954543, 0.1954561, 0.1954556, 0.1954564, 0.195456, 0.195456, 
    0.1954554, 0.1954551, 0.1954543, 0.1954536, 0.1954531, 0.1954533, 
    0.1954538, 0.1954548, 0.1954558, 0.1954556, 0.1954564, 0.1954544, 
    0.1954552, 0.1954549, 0.1954557, 0.1954539, 0.1954554, 0.1954536, 
    0.1954537, 0.1954542, 0.1954553, 0.1954555, 0.1954558, 0.1954556, 
    0.1954549, 0.1954547, 0.1954542, 0.1954541, 0.1954537, 0.1954534, 
    0.1954537, 0.195454, 0.1954549, 0.1954557, 0.1954566, 0.1954568, 
    0.1954579, 0.195457, 0.1954585, 0.1954572, 0.1954595, 0.1954555, 
    0.1954572, 0.1954543, 0.1954546, 0.1954551, 0.1954564, 0.1954557, 
    0.1954566, 0.1954547, 0.1954538, 0.1954536, 0.1954532, 0.1954536, 
    0.1954536, 0.195454, 0.1954539, 0.1954549, 0.1954543, 0.195456, 
    0.1954566, 0.1954584, 0.1954596, 0.1954608, 0.1954614, 0.1954615, 
    0.1954616,
  0.1982628, 0.1982629, 0.1982629, 0.198263, 0.1982629, 0.198263, 0.1982629, 
    0.1982629, 0.1982629, 0.1982629, 0.1982631, 0.198263, 0.1982633, 
    0.1982632, 0.1982635, 0.1982633, 0.1982635, 0.1982635, 0.1982636, 
    0.1982636, 0.1982638, 0.1982637, 0.1982639, 0.1982637, 0.1982638, 
    0.1982637, 0.198263, 0.1982631, 0.198263, 0.198263, 0.198263, 0.1982629, 
    0.1982629, 0.1982628, 0.1982629, 0.1982629, 0.198263, 0.198263, 
    0.1982631, 0.1982631, 0.1982633, 0.1982632, 0.1982635, 0.1982634, 
    0.1982636, 0.1982635, 0.1982636, 0.1982636, 0.1982636, 0.1982635, 
    0.1982635, 0.1982635, 0.1982632, 0.1982633, 0.1982631, 0.1982629, 
    0.1982629, 0.1982628, 0.1982628, 0.1982628, 0.1982629, 0.198263, 
    0.198263, 0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982635, 
    0.1982634, 0.1982635, 0.1982635, 0.1982636, 0.1982636, 0.1982636, 
    0.1982635, 0.1982636, 0.1982634, 0.1982635, 0.1982631, 0.198263, 
    0.198263, 0.1982629, 0.1982628, 0.1982629, 0.1982629, 0.1982629, 
    0.198263, 0.1982629, 0.1982631, 0.198263, 0.1982633, 0.1982632, 
    0.1982635, 0.1982634, 0.1982635, 0.1982635, 0.1982636, 0.1982635, 
    0.1982637, 0.1982637, 0.1982637, 0.1982638, 0.1982635, 0.1982636, 
    0.1982629, 0.1982629, 0.198263, 0.1982629, 0.1982629, 0.1982628, 
    0.1982629, 0.1982629, 0.198263, 0.198263, 0.198263, 0.1982631, 0.1982632, 
    0.1982633, 0.1982634, 0.1982635, 0.1982635, 0.1982635, 0.1982635, 
    0.1982635, 0.1982637, 0.1982635, 0.1982637, 0.1982637, 0.1982636, 
    0.1982637, 0.198263, 0.1982629, 0.1982629, 0.1982629, 0.1982628, 
    0.1982629, 0.1982629, 0.198263, 0.198263, 0.1982631, 0.1982631, 
    0.1982632, 0.1982633, 0.1982634, 0.1982635, 0.1982635, 0.1982635, 
    0.1982636, 0.1982635, 0.1982636, 0.1982636, 0.1982635, 0.1982637, 
    0.1982637, 0.1982637, 0.1982637, 0.1982629, 0.198263, 0.198263, 0.198263, 
    0.198263, 0.1982631, 0.1982631, 0.1982633, 0.1982632, 0.1982633, 
    0.1982632, 0.1982632, 0.1982633, 0.1982632, 0.1982634, 0.1982633, 
    0.1982636, 0.1982634, 0.1982636, 0.1982635, 0.1982636, 0.1982636, 
    0.1982637, 0.1982638, 0.1982638, 0.1982639, 0.198263, 0.1982631, 
    0.1982631, 0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982633, 
    0.1982634, 0.1982634, 0.1982633, 0.1982633, 0.1982631, 0.1982631, 
    0.1982631, 0.198263, 0.1982633, 0.1982632, 0.1982635, 0.1982634, 
    0.1982636, 0.1982635, 0.1982638, 0.1982639, 0.198264, 0.1982642, 
    0.1982631, 0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982634, 
    0.1982634, 0.1982634, 0.1982635, 0.1982635, 0.1982634, 0.1982635, 
    0.1982631, 0.1982633, 0.198263, 0.1982631, 0.1982632, 0.1982632, 
    0.1982633, 0.1982633, 0.1982635, 0.1982634, 0.1982639, 0.1982636, 
    0.1982643, 0.1982641, 0.198263, 0.1982631, 0.1982632, 0.1982632, 
    0.1982634, 0.1982634, 0.1982635, 0.1982635, 0.1982635, 0.1982636, 
    0.1982635, 0.1982636, 0.1982634, 0.1982635, 0.1982632, 0.1982633, 
    0.1982632, 0.1982632, 0.1982633, 0.1982634, 0.1982634, 0.1982634, 
    0.1982635, 0.1982634, 0.1982639, 0.1982636, 0.1982631, 0.1982632, 
    0.1982632, 0.1982632, 0.1982634, 0.1982633, 0.1982636, 0.1982635, 
    0.1982636, 0.1982636, 0.1982636, 0.1982635, 0.1982634, 0.1982633, 
    0.1982633, 0.1982632, 0.1982632, 0.1982633, 0.1982634, 0.1982635, 
    0.1982635, 0.1982636, 0.1982633, 0.1982635, 0.1982634, 0.1982635, 
    0.1982633, 0.1982635, 0.1982632, 0.1982633, 0.1982633, 0.1982635, 
    0.1982635, 0.1982635, 0.1982635, 0.1982634, 0.1982634, 0.1982633, 
    0.1982633, 0.1982633, 0.1982632, 0.1982633, 0.1982633, 0.1982634, 
    0.1982635, 0.1982636, 0.1982637, 0.1982638, 0.1982637, 0.1982639, 
    0.1982637, 0.198264, 0.1982635, 0.1982637, 0.1982633, 0.1982634, 
    0.1982634, 0.1982636, 0.1982635, 0.1982636, 0.1982634, 0.1982633, 
    0.1982633, 0.1982632, 0.1982633, 0.1982632, 0.1982633, 0.1982633, 
    0.1982634, 0.1982633, 0.1982636, 0.1982636, 0.1982639, 0.198264, 
    0.1982642, 0.1982643, 0.1982643, 0.1982643,
  0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  8.601481, 8.601533, 8.601523, 8.601563, 8.601542, 8.601567, 8.601493, 
    8.601534, 8.601508, 8.601487, 8.601641, 8.601565, 8.601724, 8.601675, 
    8.601799, 8.601716, 8.601816, 8.601798, 8.601856, 8.601839, 8.601912, 
    8.601864, 8.601951, 8.601901, 8.601908, 8.601862, 8.601582, 8.601631, 
    8.601579, 8.601585, 8.601583, 8.601542, 8.601521, 8.601479, 8.601486, 
    8.601517, 8.601589, 8.601565, 8.601627, 8.601625, 8.601693, 8.601663, 
    8.601778, 8.601746, 8.60184, 8.601816, 8.601839, 8.601832, 8.601839, 
    8.601804, 8.601819, 8.601789, 8.601668, 8.601704, 8.601599, 8.601534, 
    8.601494, 8.601465, 8.601469, 8.601477, 8.601518, 8.601557, 8.601586, 
    8.601605, 8.601625, 8.601682, 8.601714, 8.601784, 8.601772, 8.601793, 
    8.601814, 8.601848, 8.601843, 8.601857, 8.601793, 8.601835, 8.601766, 
    8.601785, 8.601627, 8.601572, 8.601545, 8.601524, 8.601472, 8.601508, 
    8.601494, 8.601529, 8.60155, 8.60154, 8.601606, 8.601581, 8.601716, 
    8.601657, 8.601811, 8.601774, 8.60182, 8.601797, 8.601836, 8.601801, 
    8.601863, 8.601876, 8.601867, 8.601903, 8.601799, 8.601838, 8.60154, 
    8.601542, 8.601549, 8.601513, 8.601511, 8.601478, 8.601507, 8.60152, 
    8.601552, 8.60157, 8.601588, 8.601627, 8.60167, 8.601732, 8.601777, 
    8.601807, 8.601789, 8.601805, 8.601787, 8.601779, 8.601871, 8.601819, 
    8.601898, 8.601893, 8.601857, 8.601894, 8.601542, 8.601532, 8.601497, 
    8.601524, 8.601475, 8.601502, 8.601518, 8.60158, 8.601595, 8.601607, 
    8.601632, 8.601665, 8.60172, 8.601769, 8.601815, 8.601812, 8.601813, 
    8.601823, 8.601798, 8.601827, 8.601831, 8.601819, 8.601893, 8.601872, 
    8.601893, 8.60188, 8.601536, 8.601553, 8.601543, 8.601561, 8.601548, 
    8.601602, 8.601618, 8.601694, 8.601664, 8.601713, 8.601668, 8.601676, 
    8.601713, 8.601671, 8.601767, 8.601701, 8.601823, 8.601756, 8.601828, 
    8.601815, 8.601836, 8.601854, 8.601878, 8.60192, 8.601911, 8.601947, 
    8.601578, 8.6016, 8.601599, 8.601622, 8.601638, 8.601675, 8.601735, 
    8.601712, 8.601754, 8.601762, 8.6017, 8.601737, 8.601614, 8.601633, 
    8.601623, 8.60158, 8.601717, 8.601645, 8.601778, 8.601739, 8.601851, 
    8.601795, 8.601905, 8.601951, 8.601996, 8.602047, 8.601612, 8.601597, 
    8.601624, 8.60166, 8.601695, 8.601742, 8.601747, 8.601755, 8.601778, 
    8.601796, 8.601757, 8.601801, 8.601637, 8.601724, 8.601591, 8.60163, 
    8.601659, 8.601646, 8.60171, 8.601725, 8.601785, 8.601754, 8.601939, 
    8.601857, 8.602088, 8.602022, 8.601592, 8.601612, 8.601682, 8.601648, 
    8.601745, 8.601768, 8.601788, 8.601811, 8.601815, 8.60183, 8.601806, 
    8.601829, 8.601742, 8.601781, 8.601675, 8.6017, 8.601688, 8.601676, 
    8.601716, 8.601757, 8.601759, 8.601772, 8.601808, 8.601746, 8.601948, 
    8.601821, 8.601634, 8.601672, 8.601679, 8.601664, 8.601766, 8.601728, 
    8.601829, 8.601802, 8.601847, 8.601825, 8.601821, 8.601793, 8.601775, 
    8.60173, 8.601694, 8.601666, 8.601672, 8.601704, 8.60176, 8.601814, 
    8.601803, 8.601843, 8.601738, 8.601782, 8.601765, 8.60181, 8.601712, 
    8.601791, 8.601691, 8.6017, 8.601728, 8.601784, 8.601797, 8.60181, 
    8.601803, 8.601762, 8.601756, 8.601727, 8.601719, 8.601698, 8.601681, 
    8.601696, 8.601713, 8.601763, 8.601806, 8.601854, 8.601867, 8.60192, 
    8.601875, 8.601948, 8.601884, 8.601996, 8.601798, 8.601884, 8.601729, 
    8.601747, 8.601776, 8.601846, 8.60181, 8.601852, 8.601755, 8.601704, 
    8.601692, 8.601667, 8.601692, 8.60169, 8.601714, 8.601707, 8.601764, 
    8.601733, 8.601821, 8.601852, 8.601943, 8.601998, 8.602056, 8.602081, 
    8.602089, 8.602092 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  3.955521e-15, 3.955926e-15, 3.955849e-15, 3.956172e-15, 3.955995e-15, 
    3.956205e-15, 3.955607e-15, 3.955939e-15, 3.955729e-15, 3.955563e-15, 
    3.956788e-15, 3.956187e-15, 3.957447e-15, 3.957057e-15, 3.958049e-15, 
    3.957382e-15, 3.958185e-15, 3.958037e-15, 3.9585e-15, 3.958368e-15, 
    3.958945e-15, 3.958562e-15, 3.959258e-15, 3.958858e-15, 3.958917e-15, 
    3.958548e-15, 3.956315e-15, 3.956711e-15, 3.95629e-15, 3.956347e-15, 
    3.956323e-15, 3.955996e-15, 3.955827e-15, 3.955496e-15, 3.955557e-15, 
    3.955803e-15, 3.956372e-15, 3.956184e-15, 3.956674e-15, 3.956663e-15, 
    3.957204e-15, 3.95696e-15, 3.957877e-15, 3.957618e-15, 3.958374e-15, 
    3.958182e-15, 3.958364e-15, 3.958309e-15, 3.958364e-15, 3.958084e-15, 
    3.958204e-15, 3.957959e-15, 3.957004e-15, 3.957282e-15, 3.95645e-15, 
    3.955939e-15, 3.95562e-15, 3.955388e-15, 3.95542e-15, 3.955481e-15, 
    3.955805e-15, 3.956116e-15, 3.956351e-15, 3.956507e-15, 3.956662e-15, 
    3.957111e-15, 3.957366e-15, 3.957925e-15, 3.957831e-15, 3.957996e-15, 
    3.958164e-15, 3.958436e-15, 3.958392e-15, 3.958511e-15, 3.957996e-15, 
    3.958336e-15, 3.957776e-15, 3.957928e-15, 3.956677e-15, 3.956236e-15, 
    3.956026e-15, 3.955863e-15, 3.955445e-15, 3.955732e-15, 3.955618e-15, 
    3.955895e-15, 3.956067e-15, 3.955983e-15, 3.956511e-15, 3.956305e-15, 
    3.957381e-15, 3.956917e-15, 3.958144e-15, 3.957851e-15, 3.958215e-15, 
    3.958031e-15, 3.958345e-15, 3.958062e-15, 3.958557e-15, 3.958661e-15, 
    3.958589e-15, 3.958876e-15, 3.958046e-15, 3.958361e-15, 3.955979e-15, 
    3.955992e-15, 3.956059e-15, 3.955768e-15, 3.955751e-15, 3.955493e-15, 
    3.955725e-15, 3.955822e-15, 3.956079e-15, 3.956226e-15, 3.956367e-15, 
    3.956679e-15, 3.957023e-15, 3.957513e-15, 3.957869e-15, 3.958108e-15, 
    3.957963e-15, 3.958091e-15, 3.957947e-15, 3.957882e-15, 3.95862e-15, 
    3.958203e-15, 3.958835e-15, 3.9588e-15, 3.958512e-15, 3.958805e-15, 
    3.956003e-15, 3.955924e-15, 3.955642e-15, 3.955863e-15, 3.955465e-15, 
    3.955684e-15, 3.955808e-15, 3.956303e-15, 3.956418e-15, 3.956517e-15, 
    3.956717e-15, 3.956972e-15, 3.957418e-15, 3.957811e-15, 3.958174e-15, 
    3.958149e-15, 3.958157e-15, 3.958236e-15, 3.958038e-15, 3.958268e-15, 
    3.958305e-15, 3.958206e-15, 3.958796e-15, 3.958628e-15, 3.9588e-15, 
    3.958691e-15, 3.95595e-15, 3.956084e-15, 3.956011e-15, 3.956146e-15, 
    3.956049e-15, 3.956474e-15, 3.956602e-15, 3.957208e-15, 3.956966e-15, 
    3.957359e-15, 3.957008e-15, 3.957069e-15, 3.95736e-15, 3.957028e-15, 
    3.957784e-15, 3.957262e-15, 3.958239e-15, 3.957705e-15, 3.958272e-15, 
    3.958173e-15, 3.958339e-15, 3.958485e-15, 3.958675e-15, 3.959015e-15, 
    3.958938e-15, 3.959228e-15, 3.956285e-15, 3.956457e-15, 3.956447e-15, 
    3.956629e-15, 3.956764e-15, 3.957061e-15, 3.957532e-15, 3.957357e-15, 
    3.957685e-15, 3.95775e-15, 3.957253e-15, 3.957553e-15, 3.956575e-15, 
    3.956728e-15, 3.95664e-15, 3.956296e-15, 3.95739e-15, 3.956825e-15, 
    3.957875e-15, 3.957569e-15, 3.958464e-15, 3.958013e-15, 3.958894e-15, 
    3.959258e-15, 3.959625e-15, 3.960027e-15, 3.956556e-15, 3.956439e-15, 
    3.956653e-15, 3.956939e-15, 3.957221e-15, 3.957587e-15, 3.957627e-15, 
    3.957694e-15, 3.957874e-15, 3.958023e-15, 3.95771e-15, 3.958061e-15, 
    3.956753e-15, 3.957442e-15, 3.95639e-15, 3.956699e-15, 3.956925e-15, 
    3.956831e-15, 3.957338e-15, 3.957456e-15, 3.957933e-15, 3.957689e-15, 
    3.959163e-15, 3.958509e-15, 3.960351e-15, 3.959831e-15, 3.956397e-15, 
    3.956558e-15, 3.957111e-15, 3.956848e-15, 3.957614e-15, 3.9578e-15, 
    3.957956e-15, 3.958147e-15, 3.958172e-15, 3.958286e-15, 3.958099e-15, 
    3.958281e-15, 3.957587e-15, 3.957897e-15, 3.957054e-15, 3.957256e-15, 
    3.957165e-15, 3.957061e-15, 3.957381e-15, 3.957714e-15, 3.957729e-15, 
    3.957834e-15, 3.958117e-15, 3.957617e-15, 3.959233e-15, 3.958219e-15, 
    3.956733e-15, 3.957032e-15, 3.957085e-15, 3.956967e-15, 3.957781e-15, 
    3.957485e-15, 3.958284e-15, 3.95807e-15, 3.958424e-15, 3.958247e-15, 
    3.958221e-15, 3.957996e-15, 3.957854e-15, 3.957497e-15, 3.957209e-15, 
    3.956985e-15, 3.957038e-15, 3.957284e-15, 3.957736e-15, 3.958171e-15, 
    3.958074e-15, 3.958397e-15, 3.957558e-15, 3.957905e-15, 3.957768e-15, 
    3.958127e-15, 3.95735e-15, 3.957987e-15, 3.957185e-15, 3.957257e-15, 
    3.957479e-15, 3.957923e-15, 3.958034e-15, 3.958137e-15, 3.958075e-15, 
    3.957749e-15, 3.957699e-15, 3.957476e-15, 3.95741e-15, 3.957242e-15, 
    3.957099e-15, 3.957227e-15, 3.957361e-15, 3.957753e-15, 3.958102e-15, 
    3.958486e-15, 3.958583e-15, 3.959013e-15, 3.958652e-15, 3.959237e-15, 
    3.958723e-15, 3.959622e-15, 3.958035e-15, 3.958724e-15, 3.957492e-15, 
    3.957626e-15, 3.957861e-15, 3.958417e-15, 3.958125e-15, 3.958471e-15, 
    3.957698e-15, 3.957288e-15, 3.957193e-15, 3.956997e-15, 3.957197e-15, 
    3.957181e-15, 3.957372e-15, 3.957311e-15, 3.957766e-15, 3.957522e-15, 
    3.958218e-15, 3.95847e-15, 3.959195e-15, 3.959635e-15, 3.960097e-15, 
    3.960297e-15, 3.960358e-15, 3.960384e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  9.872261, 9.920599, 9.911189, 9.950092, 9.928573, 9.953949, 9.882047, 
    9.922523, 9.89667, 9.876603, 10.02506, 9.951811, 10.10145, 10.05449, 
    10.1727, 10.09414, 10.18858, 10.17042, 10.22512, 10.20943, 10.2796, 
    10.23237, 10.31608, 10.26831, 10.27577, 10.23081, 9.966517, 10.01592, 
    9.963596, 9.970631, 9.967472, 9.929023, 9.909469, 9.868567, 9.875984, 
    9.906026, 9.973795, 9.95092, 10.00862, 10.00731, 10.07178, 10.04268, 
    10.15141, 10.12043, 10.21008, 10.1875, 10.20902, 10.20249, 10.20911, 
    10.17599, 10.19017, 10.16106, 10.04813, 10.08124, 9.982681, 9.923481, 
    9.883821, 9.855742, 9.859709, 9.867274, 9.906201, 9.94282, 9.970409, 
    9.988893, 10.00712, 10.06245, 10.09179, 10.15768, 10.14576, 10.16595, 
    10.18525, 10.21771, 10.21236, 10.22668, 10.16541, 10.20611, 10.13898, 
    10.15731, 10.01211, 9.957087, 9.933701, 9.912998, 9.86276, 9.897438, 
    9.883759, 9.916315, 9.937039, 9.926785, 9.989398, 9.965098, 10.09353, 
    10.03809, 10.183, 10.14821, 10.19135, 10.16932, 10.20708, 10.17309, 
    10.23201, 10.24487, 10.23608, 10.26985, 10.17121, 10.20903, 9.926499, 
    9.928171, 9.93596, 9.90175, 9.899658, 9.868366, 9.896204, 9.908075, 
    9.938239, 9.955855, 9.972608, 10.0095, 10.05081, 10.10873, 10.15046, 
    10.17849, 10.1613, 10.17648, 10.15951, 10.15156, 10.24005, 10.19031, 
    10.26499, 10.26085, 10.22702, 10.26131, 9.929345, 9.919725, 9.886379, 
    9.91247, 9.864962, 9.891541, 9.906845, 9.965612, 9.97844, 9.990353, 
    10.0139, 10.04417, 10.09741, 10.14386, 10.18637, 10.18325, 10.18435, 
    10.19386, 10.17031, 10.19773, 10.20234, 10.1903, 10.26029, 10.24027, 
    10.26076, 10.24771, 9.922852, 9.93904, 9.930292, 9.946635, 9.935156, 
    9.986075, 10.00136, 10.07304, 10.04357, 10.09048, 10.04833, 10.05579, 
    10.09202, 10.0506, 10.1413, 10.07977, 10.19423, 10.13261, 10.1981, 
    10.18619, 10.20592, 10.22361, 10.24589, 10.28708, 10.27754, 10.31204, 
    9.962845, 9.983588, 9.981756, 10.00349, 10.01958, 10.0545, 10.11067, 
    10.08952, 10.12836, 10.13617, 10.07717, 10.11337, 9.997482, 10.01616, 
    10.00503, 9.964483, 10.0944, 10.0276, 10.15115, 10.11481, 10.22109, 
    10.16816, 10.27228, 10.317, 10.35916, 10.40859, 9.994915, 9.980808, 
    10.00607, 10.0411, 10.07365, 10.11703, 10.12147, 10.12961, 10.15071, 
    10.16848, 10.13219, 10.17294, 10.0205, 10.10021, 9.975483, 10.01295, 
    10.03903, 10.02758, 10.08711, 10.10117, 10.15844, 10.12881, 10.30596, 
    10.22736, 10.4463, 10.38485, 9.975883, 9.994864, 10.0611, 10.02955, 
    10.11992, 10.14224, 10.16041, 10.18366, 10.18617, 10.19996, 10.17737, 
    10.19907, 10.11712, 10.15369, 10.05351, 10.07784, 10.06664, 10.05437, 
    10.09228, 10.13276, 10.13362, 10.14662, 10.18334, 10.12029, 10.31614, 
    10.19494, 10.01559, 10.05227, 10.0575, 10.04328, 10.14, 10.10489, 
    10.19963, 10.17397, 10.21602, 10.19511, 10.19204, 10.16523, 10.14855, 
    10.1065, 10.07237, 10.04534, 10.05162, 10.08132, 10.13524, 10.1864, 
    10.17518, 10.21282, 10.11335, 10.155, 10.13889, 10.18091, 10.08896, 
    10.16726, 10.06901, 10.0776, 10.1042, 10.15783, 10.16971, 10.18241, 
    10.17457, 10.13661, 10.13039, 10.10355, 10.09615, 10.07573, 10.05885, 
    10.07427, 10.09049, 10.13662, 10.17831, 10.22386, 10.23503, 10.28847, 
    10.24497, 10.31682, 10.25573, 10.36161, 10.1718, 10.25392, 10.10541, 
    10.12134, 10.15021, 10.2166, 10.18072, 10.22268, 10.13015, 10.08235, 
    10.06999, 10.04698, 10.07052, 10.06861, 10.09116, 10.08391, 10.13815, 
    10.10899, 10.19197, 10.22235, 10.30842, 10.3614, 10.41548, 10.43941, 
    10.4467, 10.44975 ;

 WIND =
  8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  1.701001e-09, 1.681535e-09, 1.685283e-09, 1.669849e-09, 1.678374e-09, 
    1.668321e-09, 1.697016e-09, 1.680772e-09, 1.691104e-09, 1.69923e-09, 
    1.640732e-09, 1.669168e-09, 1.612257e-09, 1.629618e-09, 1.586731e-09, 
    1.614933e-09, 1.581169e-09, 1.587531e-09, 1.568544e-09, 1.573935e-09, 
    1.550158e-09, 1.566069e-09, 1.538125e-09, 1.553927e-09, 1.551433e-09, 
    1.566599e-09, 1.663363e-09, 1.644217e-09, 1.664512e-09, 1.661749e-09, 
    1.662988e-09, 1.678197e-09, 1.685972e-09, 1.702509e-09, 1.699481e-09, 
    1.687348e-09, 1.66051e-09, 1.66952e-09, 1.64701e-09, 1.647511e-09, 
    1.623175e-09, 1.634054e-09, 1.594258e-09, 1.605361e-09, 1.573709e-09, 
    1.581546e-09, 1.574075e-09, 1.576333e-09, 1.574046e-09, 1.585573e-09, 
    1.580613e-09, 1.590835e-09, 1.632004e-09, 1.619675e-09, 1.65704e-09, 
    1.680394e-09, 1.696297e-09, 1.707776e-09, 1.706143e-09, 1.703039e-09, 
    1.687278e-09, 1.672739e-09, 1.661835e-09, 1.654624e-09, 1.647584e-09, 
    1.626649e-09, 1.615795e-09, 1.592032e-09, 1.596267e-09, 1.589107e-09, 
    1.58233e-09, 1.571086e-09, 1.572925e-09, 1.568012e-09, 1.589296e-09, 
    1.575084e-09, 1.59869e-09, 1.59216e-09, 1.645677e-09, 1.667079e-09, 
    1.676352e-09, 1.684561e-09, 1.70489e-09, 1.690796e-09, 1.696322e-09, 
    1.683238e-09, 1.675033e-09, 1.679081e-09, 1.654428e-09, 1.663921e-09, 
    1.615156e-09, 1.635788e-09, 1.583118e-09, 1.595396e-09, 1.580204e-09, 
    1.587918e-09, 1.574747e-09, 1.586591e-09, 1.566192e-09, 1.561822e-09, 
    1.564805e-09, 1.55341e-09, 1.587253e-09, 1.574075e-09, 1.679194e-09, 
    1.678533e-09, 1.675458e-09, 1.689063e-09, 1.689903e-09, 1.702592e-09, 
    1.691292e-09, 1.686527e-09, 1.674561e-09, 1.667566e-09, 1.660974e-09, 
    1.646671e-09, 1.631e-09, 1.609605e-09, 1.594594e-09, 1.584694e-09, 
    1.59075e-09, 1.585401e-09, 1.591383e-09, 1.594203e-09, 1.563456e-09, 
    1.580566e-09, 1.555038e-09, 1.556428e-09, 1.567895e-09, 1.556272e-09, 
    1.678068e-09, 1.681881e-09, 1.69526e-09, 1.684771e-09, 1.703986e-09, 
    1.693173e-09, 1.687021e-09, 1.66372e-09, 1.658693e-09, 1.654058e-09, 
    1.644985e-09, 1.633493e-09, 1.613735e-09, 1.596947e-09, 1.581938e-09, 
    1.583028e-09, 1.582644e-09, 1.579328e-09, 1.587569e-09, 1.577983e-09, 
    1.576386e-09, 1.580569e-09, 1.556615e-09, 1.563381e-09, 1.556458e-09, 
    1.560856e-09, 1.68064e-09, 1.674245e-09, 1.677694e-09, 1.671221e-09, 
    1.675776e-09, 1.65572e-09, 1.649806e-09, 1.62271e-09, 1.633717e-09, 
    1.616274e-09, 1.631928e-09, 1.629131e-09, 1.61571e-09, 1.631074e-09, 
    1.597863e-09, 1.620221e-09, 1.579199e-09, 1.600978e-09, 1.577855e-09, 
    1.582002e-09, 1.575148e-09, 1.569061e-09, 1.561473e-09, 1.54767e-09, 
    1.550844e-09, 1.539446e-09, 1.664808e-09, 1.656687e-09, 1.657399e-09, 
    1.648983e-09, 1.642815e-09, 1.629614e-09, 1.608899e-09, 1.616624e-09, 
    1.602502e-09, 1.599698e-09, 1.621177e-09, 1.607917e-09, 1.651299e-09, 
    1.644123e-09, 1.648388e-09, 1.664164e-09, 1.614836e-09, 1.639761e-09, 
    1.594349e-09, 1.607396e-09, 1.569926e-09, 1.588329e-09, 1.552597e-09, 
    1.537825e-09, 1.524189e-09, 1.508565e-09, 1.652291e-09, 1.657769e-09, 
    1.647988e-09, 1.634653e-09, 1.622483e-09, 1.606594e-09, 1.604987e-09, 
    1.602052e-09, 1.594504e-09, 1.588214e-09, 1.601126e-09, 1.586645e-09, 
    1.642467e-09, 1.61271e-09, 1.659849e-09, 1.645351e-09, 1.635433e-09, 
    1.639769e-09, 1.617512e-09, 1.612358e-09, 1.591763e-09, 1.602341e-09, 
    1.541443e-09, 1.567781e-09, 1.49689e-09, 1.516024e-09, 1.659691e-09, 
    1.65231e-09, 1.627148e-09, 1.639019e-09, 1.605545e-09, 1.597524e-09, 
    1.591065e-09, 1.582886e-09, 1.582009e-09, 1.57721e-09, 1.58509e-09, 
    1.57752e-09, 1.60656e-09, 1.593446e-09, 1.629984e-09, 1.62093e-09, 
    1.625082e-09, 1.629662e-09, 1.615613e-09, 1.600921e-09, 1.600611e-09, 
    1.595961e-09, 1.583005e-09, 1.605412e-09, 1.538108e-09, 1.578958e-09, 
    1.644339e-09, 1.630453e-09, 1.628492e-09, 1.633827e-09, 1.598324e-09, 
    1.611e-09, 1.577327e-09, 1.586282e-09, 1.571664e-09, 1.578893e-09, 
    1.579962e-09, 1.589362e-09, 1.595273e-09, 1.610414e-09, 1.622957e-09, 
    1.633051e-09, 1.630692e-09, 1.619645e-09, 1.600032e-09, 1.581929e-09, 
    1.585858e-09, 1.572765e-09, 1.607924e-09, 1.592983e-09, 1.598723e-09, 
    1.583846e-09, 1.61683e-09, 1.58865e-09, 1.624202e-09, 1.621018e-09, 
    1.611253e-09, 1.591979e-09, 1.587781e-09, 1.583323e-09, 1.586071e-09, 
    1.59954e-09, 1.60177e-09, 1.61149e-09, 1.614194e-09, 1.62171e-09, 
    1.627988e-09, 1.62225e-09, 1.616269e-09, 1.599535e-09, 1.584761e-09, 
    1.568974e-09, 1.565161e-09, 1.547214e-09, 1.56179e-09, 1.537887e-09, 
    1.558157e-09, 1.523412e-09, 1.58705e-09, 1.558764e-09, 1.610812e-09, 
    1.605032e-09, 1.594684e-09, 1.57147e-09, 1.583915e-09, 1.569382e-09, 
    1.601858e-09, 1.619266e-09, 1.623836e-09, 1.632434e-09, 1.623641e-09, 
    1.624352e-09, 1.616023e-09, 1.61869e-09, 1.598986e-09, 1.609507e-09, 
    1.579989e-09, 1.569496e-09, 1.540632e-09, 1.523476e-09, 1.506416e-09, 
    1.499008e-09, 1.496769e-09, 1.495834e-09 ;

 W_SCALAR =
  0.6251647, 0.6268236, 0.6265013, 0.6278382, 0.6270967, 0.6279719, 
    0.6255011, 0.6268895, 0.6260033, 0.625314, 0.6304291, 0.6278978, 
    0.6330526, 0.6314422, 0.6354835, 0.6328022, 0.6360235, 0.6354061, 
    0.6372628, 0.6367311, 0.6391034, 0.6375081, 0.6403309, 0.6387225, 
    0.6389743, 0.6374555, 0.6284074, 0.6301143, 0.6283063, 0.6285498, 
    0.6284405, 0.627112, 0.6264422, 0.6250377, 0.6252927, 0.6263242, 
    0.6286593, 0.627867, 0.6298626, 0.6298175, 0.6320359, 0.6310362, 
    0.6347587, 0.6337017, 0.6367534, 0.6359866, 0.6367174, 0.6364958, 
    0.6367203, 0.6355956, 0.6360776, 0.6350874, 0.6312234, 0.6323603, 
    0.6289667, 0.6269222, 0.6255621, 0.6245962, 0.6247327, 0.6249931, 
    0.6263303, 0.627586, 0.6285422, 0.6291815, 0.6298111, 0.6317154, 
    0.6327217, 0.6349724, 0.6345664, 0.635254, 0.6359103, 0.6370117, 
    0.6368305, 0.6373155, 0.6352357, 0.6366184, 0.634335, 0.63496, 0.6299828, 
    0.6280808, 0.627272, 0.6265633, 0.6248378, 0.6260296, 0.6255599, 
    0.626677, 0.6273863, 0.6270355, 0.629199, 0.6283583, 0.6327813, 0.630878, 
    0.6358338, 0.6346497, 0.6361175, 0.6353686, 0.6366514, 0.635497, 
    0.6374959, 0.6379308, 0.6376337, 0.6387746, 0.635433, 0.6367174, 
    0.6270257, 0.6270829, 0.6273494, 0.6261775, 0.6261058, 0.6250307, 
    0.6259873, 0.6263945, 0.6274274, 0.628038, 0.6286183, 0.6298931, 
    0.6313155, 0.6333016, 0.6347265, 0.6356807, 0.6350957, 0.6356122, 
    0.6350347, 0.634764, 0.637768, 0.6360821, 0.6386105, 0.6384708, 
    0.6373271, 0.6384865, 0.6271231, 0.6267938, 0.6256499, 0.6265452, 
    0.6249136, 0.6258272, 0.6263523, 0.6283761, 0.6288201, 0.6292319, 
    0.6300448, 0.6310873, 0.6329141, 0.6345014, 0.6359485, 0.6358425, 
    0.6358798, 0.6362029, 0.6354025, 0.6363343, 0.6364907, 0.6360819, 
    0.6384521, 0.6377754, 0.6384678, 0.6380273, 0.6269008, 0.6274548, 
    0.6271555, 0.6277183, 0.6273219, 0.6290841, 0.6296119, 0.6320789, 
    0.6310669, 0.632677, 0.6312305, 0.6314869, 0.6327297, 0.6313086, 
    0.634414, 0.6323097, 0.6362155, 0.6341174, 0.6363469, 0.6359422, 
    0.6366121, 0.6372117, 0.6379656, 0.6393555, 0.6390338, 0.6401951, 
    0.6282803, 0.6289981, 0.6289348, 0.6296856, 0.6302406, 0.6314425, 
    0.633368, 0.6326442, 0.6339725, 0.634239, 0.6322209, 0.6334605, 
    0.6294782, 0.6301226, 0.6297389, 0.628337, 0.6328112, 0.630517, 0.63475, 
    0.6335096, 0.6371263, 0.6353291, 0.6388566, 0.6403618, 0.6417761, 
    0.6434274, 0.6293896, 0.628902, 0.6297748, 0.6309816, 0.6320999, 
    0.6335853, 0.6337371, 0.6340152, 0.6347351, 0.6353402, 0.6341032, 
    0.6354917, 0.6302722, 0.6330101, 0.6287178, 0.6300119, 0.6309104, 
    0.6305162, 0.6325614, 0.6330431, 0.6349983, 0.6339878, 0.6399906, 
    0.6373385, 0.6446828, 0.642635, 0.6287317, 0.6293879, 0.6316692, 
    0.6305842, 0.6336843, 0.6344463, 0.6350653, 0.6358563, 0.6359416, 
    0.6364099, 0.6356423, 0.6363796, 0.6335885, 0.6348366, 0.6314085, 
    0.6322438, 0.6318595, 0.6314381, 0.6327385, 0.6341228, 0.6341521, 
    0.6345957, 0.6358451, 0.6336969, 0.6403329, 0.6362392, 0.6301031, 
    0.6313656, 0.6315456, 0.6310568, 0.63437, 0.6331705, 0.6363985, 
    0.6355269, 0.6369547, 0.6362454, 0.6361411, 0.6352293, 0.6346615, 
    0.6332256, 0.632056, 0.6311277, 0.6313435, 0.6323631, 0.6342074, 
    0.6359494, 0.635568, 0.6368462, 0.6334598, 0.634881, 0.634332, 0.635763, 
    0.632625, 0.6352983, 0.6319409, 0.6322356, 0.6331467, 0.6349775, 
    0.6353819, 0.6358139, 0.6355473, 0.6342541, 0.634042, 0.6331245, 
    0.6328712, 0.6321714, 0.6315919, 0.6321214, 0.6326774, 0.6342546, 
    0.6356743, 0.6372203, 0.6375982, 0.639402, 0.6379341, 0.6403556, 
    0.6382976, 0.6418577, 0.6354527, 0.6382366, 0.6331881, 0.6337329, 
    0.634718, 0.6369739, 0.6357563, 0.6371801, 0.6340337, 0.6323984, 
    0.6319746, 0.6311842, 0.6319927, 0.631927, 0.6327003, 0.6324518, 
    0.6343069, 0.6333107, 0.6361384, 0.6371688, 0.6400735, 0.6418509, 
    0.643657, 0.6444536, 0.6446959, 0.6447972,
  0.546157, 0.5482014, 0.5478041, 0.5494519, 0.5485379, 0.5496167, 0.5465716, 
    0.5482826, 0.5471904, 0.546341, 0.5526459, 0.5495253, 0.555881, 
    0.5538949, 0.5588794, 0.5555722, 0.5595455, 0.5587839, 0.5610747, 
    0.5604187, 0.563346, 0.5613773, 0.5648611, 0.5628759, 0.5631867, 
    0.5613124, 0.5501536, 0.5522578, 0.5500289, 0.550329, 0.5501943, 
    0.5485569, 0.5477313, 0.5460005, 0.5463148, 0.5475859, 0.550464, 
    0.5494874, 0.5519474, 0.5518919, 0.554627, 0.5533943, 0.5579852, 
    0.5566816, 0.5604461, 0.5595002, 0.5604017, 0.5601283, 0.5604053, 
    0.5590177, 0.5596123, 0.5583908, 0.5536253, 0.5550272, 0.550843, 
    0.5483229, 0.5466467, 0.5454565, 0.5456248, 0.5459456, 0.5475933, 
    0.549141, 0.5503197, 0.5511078, 0.5518839, 0.5542318, 0.5554729, 
    0.5582489, 0.557748, 0.5585963, 0.559406, 0.5607648, 0.5605412, 
    0.5611397, 0.5585737, 0.5602796, 0.5574627, 0.5582336, 0.5520956, 
    0.5497509, 0.548754, 0.5478805, 0.5457542, 0.5472229, 0.546644, 
    0.5480206, 0.5488949, 0.5484625, 0.5511293, 0.550093, 0.5555463, 
    0.5531994, 0.5593116, 0.5578508, 0.5596615, 0.5587378, 0.5603203, 
    0.5588961, 0.5613623, 0.561899, 0.5615323, 0.5629402, 0.5588171, 
    0.5604017, 0.5484505, 0.548521, 0.5488495, 0.5474051, 0.5473167, 
    0.5459919, 0.5471707, 0.5476725, 0.5489455, 0.5496982, 0.5504134, 
    0.551985, 0.5537388, 0.556188, 0.5579455, 0.5591227, 0.5584009, 
    0.5590382, 0.5583258, 0.5579918, 0.561698, 0.5596179, 0.5627378, 
    0.5625653, 0.5611539, 0.5625847, 0.5485705, 0.5481646, 0.546755, 
    0.5478582, 0.5458476, 0.5469734, 0.5476205, 0.5501148, 0.5506622, 
    0.5511699, 0.5521721, 0.5534574, 0.5557102, 0.5576679, 0.5594531, 
    0.5593223, 0.5593683, 0.559767, 0.5587795, 0.5599291, 0.560122, 
    0.5596176, 0.5625422, 0.5617071, 0.5625616, 0.5620179, 0.5482965, 
    0.5489793, 0.5486104, 0.5493042, 0.5488155, 0.5509876, 0.5516384, 
    0.5546801, 0.5534322, 0.5554177, 0.5536339, 0.5539501, 0.5554827, 
    0.5537303, 0.5575601, 0.5549648, 0.5597825, 0.5571942, 0.5599446, 
    0.5594453, 0.5602717, 0.5610116, 0.5619419, 0.5636572, 0.5632601, 
    0.5646935, 0.5499968, 0.5508817, 0.5508036, 0.5517291, 0.5524134, 
    0.5538954, 0.5562699, 0.5553773, 0.5570155, 0.5573443, 0.5548552, 
    0.556384, 0.5514736, 0.5522679, 0.5517949, 0.5500666, 0.5555832, 
    0.5527542, 0.5579746, 0.5564446, 0.5609062, 0.5586889, 0.5630415, 
    0.5648993, 0.5666452, 0.568684, 0.5513642, 0.5507632, 0.5518392, 
    0.553327, 0.554706, 0.556538, 0.5567252, 0.5570682, 0.5579562, 0.5587025, 
    0.5571768, 0.5588896, 0.5524524, 0.5558285, 0.5505361, 0.5521315, 
    0.5532393, 0.5527533, 0.5552752, 0.5558692, 0.5582808, 0.5570344, 
    0.5644411, 0.5611681, 0.5702342, 0.5677056, 0.5505532, 0.5513622, 
    0.554175, 0.5528371, 0.5566601, 0.5576, 0.5583635, 0.5593393, 0.5594445, 
    0.5600224, 0.5590754, 0.5599849, 0.5565419, 0.5580813, 0.5538535, 
    0.5548835, 0.5544097, 0.5538899, 0.5554936, 0.5572008, 0.5572371, 
    0.5577842, 0.5593255, 0.5566756, 0.5648635, 0.5598118, 0.5522438, 
    0.5538005, 0.5540225, 0.5534198, 0.5575058, 0.5560263, 0.5600083, 
    0.558933, 0.5606945, 0.5598193, 0.5596906, 0.5585659, 0.5578654, 
    0.5560943, 0.5546519, 0.5535071, 0.5537734, 0.5550306, 0.5573052, 
    0.5594542, 0.5589837, 0.5605606, 0.5563832, 0.5581362, 0.5574589, 
    0.5592243, 0.5553536, 0.558651, 0.5545099, 0.5548733, 0.555997, 
    0.5582552, 0.5587541, 0.559287, 0.5589581, 0.5573629, 0.5571012, 
    0.5559696, 0.5556571, 0.5547942, 0.5540795, 0.5547326, 0.5554181, 
    0.5573635, 0.5591148, 0.5610222, 0.5614886, 0.5637145, 0.5619031, 
    0.5648916, 0.5623516, 0.5667459, 0.5588415, 0.5622764, 0.556048, 0.55672, 
    0.5579351, 0.5607182, 0.559216, 0.5609726, 0.557091, 0.5550741, 
    0.5545516, 0.5535768, 0.5545738, 0.5544928, 0.5554464, 0.55514, 0.557428, 
    0.5561993, 0.5596874, 0.5609587, 0.5645434, 0.5667375, 0.5689675, 
    0.5699512, 0.5702505, 0.5703756,
  0.5139313, 0.5161815, 0.5157441, 0.5175582, 0.516552, 0.5177397, 0.5143875, 
    0.5162709, 0.5150687, 0.5141338, 0.5210757, 0.5176391, 0.5246401, 
    0.5224517, 0.5279453, 0.5242998, 0.5286797, 0.52784, 0.5303661, 
    0.5296426, 0.5328715, 0.5306999, 0.5345433, 0.5323529, 0.5326958, 
    0.5306283, 0.5183308, 0.5206482, 0.5181935, 0.5185241, 0.5183757, 
    0.5165728, 0.515664, 0.5137591, 0.514105, 0.515504, 0.5186727, 0.5175973, 
    0.5203063, 0.5202452, 0.5232583, 0.5219002, 0.5269595, 0.5255224, 
    0.5296728, 0.5286297, 0.5296239, 0.5293224, 0.5296278, 0.5280977, 
    0.5287534, 0.5274066, 0.5221546, 0.5236993, 0.51909, 0.5163153, 
    0.5144702, 0.5131604, 0.5133456, 0.5136987, 0.5155122, 0.517216, 
    0.5185137, 0.5193816, 0.5202364, 0.5228229, 0.5241903, 0.5272501, 
    0.5266979, 0.5276331, 0.5285259, 0.5300243, 0.5297777, 0.5304378, 
    0.5276083, 0.5294892, 0.5263835, 0.5272333, 0.5204695, 0.5178874, 
    0.5167899, 0.5158283, 0.513488, 0.5151044, 0.5144673, 0.5159825, 
    0.516945, 0.516469, 0.5194053, 0.5182641, 0.5242713, 0.5216854, 
    0.5284218, 0.5268112, 0.5288076, 0.5277891, 0.529534, 0.5279636, 
    0.5306833, 0.5312753, 0.5308708, 0.5324239, 0.5278766, 0.5296239, 
    0.5164557, 0.5165333, 0.5168949, 0.515305, 0.5152077, 0.5137497, 
    0.515047, 0.5155994, 0.5170007, 0.5178295, 0.518617, 0.5203478, 
    0.5222796, 0.5249785, 0.5269157, 0.5282135, 0.5274177, 0.5281203, 
    0.5273349, 0.5269667, 0.5310535, 0.5287595, 0.5322006, 0.5320103, 
    0.5304535, 0.5320317, 0.5165879, 0.516141, 0.5145894, 0.5158038, 
    0.5135908, 0.5148298, 0.515542, 0.5182882, 0.518891, 0.5194501, 
    0.5205538, 0.5219697, 0.5244519, 0.5266096, 0.5285777, 0.5284336, 
    0.5284843, 0.5289239, 0.5278351, 0.5291026, 0.5293154, 0.5287592, 
    0.5319847, 0.5310636, 0.5320062, 0.5314065, 0.5162863, 0.517038, 
    0.5166318, 0.5173956, 0.5168576, 0.5192493, 0.5199659, 0.5233168, 
    0.5219419, 0.5241295, 0.5221641, 0.5225125, 0.5242012, 0.5222703, 
    0.5264909, 0.5236305, 0.528941, 0.5260875, 0.5291197, 0.5285692, 
    0.5294805, 0.5302965, 0.5313225, 0.5332149, 0.5327768, 0.5343584, 
    0.5181582, 0.5191326, 0.5190467, 0.520066, 0.5208196, 0.5224522, 
    0.5250688, 0.524085, 0.5258905, 0.5262529, 0.5235097, 0.5251945, 
    0.5197845, 0.5206594, 0.5201384, 0.5182351, 0.524312, 0.5211951, 
    0.5269477, 0.5252612, 0.5301802, 0.5277352, 0.5325356, 0.5345855, 
    0.5365125, 0.5387634, 0.5196641, 0.5190022, 0.5201871, 0.521826, 
    0.5233454, 0.5253642, 0.5255706, 0.5259486, 0.5269275, 0.5277503, 
    0.5260683, 0.5279564, 0.5208626, 0.5245823, 0.518752, 0.5205091, 
    0.5217294, 0.521194, 0.5239726, 0.5246271, 0.5272853, 0.5259114, 
    0.5340798, 0.5304691, 0.5404754, 0.5376831, 0.5187709, 0.5196617, 
    0.5227602, 0.5212864, 0.5254988, 0.5265348, 0.5273765, 0.5284523, 
    0.5285684, 0.5292056, 0.5281613, 0.5291643, 0.5253685, 0.5270654, 
    0.522406, 0.5235409, 0.5230188, 0.5224462, 0.5242132, 0.5260948, 
    0.5261347, 0.5267379, 0.5284371, 0.5255159, 0.534546, 0.5289733, 
    0.5206329, 0.5223477, 0.5225922, 0.5219282, 0.5264309, 0.5248003, 
    0.52919, 0.5280043, 0.5299467, 0.5289817, 0.5288397, 0.5275996, 
    0.5268273, 0.5248752, 0.5232857, 0.5220245, 0.5223178, 0.523703, 
    0.5262098, 0.528579, 0.5280603, 0.5297992, 0.5251936, 0.5271259, 
    0.5263793, 0.5283255, 0.5240589, 0.5276934, 0.5231293, 0.5235297, 
    0.5247679, 0.5272571, 0.5278071, 0.5283946, 0.5280321, 0.5262734, 
    0.525985, 0.5247378, 0.5243934, 0.5234425, 0.5226551, 0.5233746, 0.52413, 
    0.526274, 0.5282048, 0.5303082, 0.5308225, 0.5332782, 0.5312797, 
    0.5345771, 0.5317745, 0.5366237, 0.5279034, 0.5316915, 0.5248242, 
    0.5255648, 0.5269042, 0.5299729, 0.5283164, 0.5302535, 0.5259737, 
    0.5237509, 0.5231752, 0.5221012, 0.5231997, 0.5231104, 0.5241612, 
    0.5238235, 0.5263452, 0.5249909, 0.5288362, 0.5302381, 0.5341928, 
    0.5366143, 0.5390764, 0.5401628, 0.5404934, 0.5406315,
  0.5071235, 0.5095142, 0.5090494, 0.5109773, 0.5099078, 0.5111702, 
    0.5076081, 0.5096092, 0.5083317, 0.5073386, 0.5147178, 0.5110633, 
    0.5185111, 0.5161818, 0.5220314, 0.5181488, 0.522814, 0.5219192, 
    0.5246115, 0.5238402, 0.5272833, 0.5249674, 0.529067, 0.5267302, 
    0.5270959, 0.524891, 0.5117986, 0.514263, 0.5116526, 0.5120041, 
    0.5118464, 0.50993, 0.5089643, 0.5069406, 0.507308, 0.5087942, 0.5121621, 
    0.5110189, 0.5138994, 0.5138344, 0.5170403, 0.515595, 0.5209812, 
    0.5194507, 0.5238724, 0.5227607, 0.5238203, 0.523499, 0.5238245, 
    0.5221938, 0.5228925, 0.5214575, 0.5158657, 0.5175096, 0.5126059, 
    0.5096563, 0.507696, 0.5063048, 0.5065015, 0.5068765, 0.5088029, 
    0.5106135, 0.5119932, 0.5129159, 0.513825, 0.5165768, 0.5180323, 
    0.5212908, 0.5207026, 0.5216988, 0.5226501, 0.5242472, 0.5239843, 
    0.5246879, 0.5216724, 0.5236768, 0.5203676, 0.5212729, 0.514073, 
    0.5113273, 0.5101607, 0.5091388, 0.5066527, 0.5083697, 0.5076929, 
    0.5093027, 0.5103256, 0.5098196, 0.5129412, 0.5117278, 0.5181186, 
    0.5153664, 0.5225391, 0.5208233, 0.5229503, 0.521865, 0.5237246, 
    0.522051, 0.5249497, 0.5255808, 0.5251496, 0.5268058, 0.5219582, 
    0.5238203, 0.5098055, 0.5098881, 0.5102723, 0.5085828, 0.5084794, 
    0.5069306, 0.5083087, 0.5088955, 0.5103848, 0.5112657, 0.512103, 
    0.5139435, 0.5159987, 0.5188715, 0.5209346, 0.5223172, 0.5214694, 
    0.5222179, 0.5213811, 0.5209889, 0.5253444, 0.5228991, 0.5265676, 
    0.5263647, 0.5247047, 0.5263875, 0.5099459, 0.5094711, 0.5078226, 
    0.5091127, 0.5067619, 0.508078, 0.5088347, 0.5117533, 0.5123942, 
    0.5129887, 0.5141626, 0.5156689, 0.5183108, 0.5206085, 0.5227054, 
    0.5225518, 0.5226058, 0.5230743, 0.521914, 0.5232648, 0.5234915, 
    0.5228987, 0.5263375, 0.5253552, 0.5263603, 0.5257208, 0.5096254, 
    0.5104244, 0.5099927, 0.5108045, 0.5102326, 0.5127752, 0.5135373, 
    0.5171025, 0.5156393, 0.5179676, 0.5158758, 0.5162466, 0.5180439, 
    0.5159888, 0.520482, 0.5174364, 0.5230925, 0.5200525, 0.5232829, 
    0.5226963, 0.5236675, 0.5245373, 0.5256313, 0.5276496, 0.5271823, 
    0.5288697, 0.5116151, 0.5126511, 0.5125598, 0.5136437, 0.5144454, 
    0.5161823, 0.5189676, 0.5179203, 0.5198427, 0.5202286, 0.5173079, 
    0.5191014, 0.5133443, 0.514275, 0.5137208, 0.5116969, 0.5181618, 
    0.5148448, 0.5209687, 0.5191725, 0.5244133, 0.5218076, 0.526925, 
    0.529112, 0.5311689, 0.5335729, 0.5132164, 0.5125125, 0.5137726, 
    0.515516, 0.5171329, 0.5192821, 0.5195019, 0.5199045, 0.5209471, 
    0.5218236, 0.520032, 0.5220433, 0.5144911, 0.5184496, 0.5122465, 
    0.5141151, 0.5154132, 0.5148436, 0.5178005, 0.5184973, 0.5213283, 
    0.5198649, 0.5285724, 0.5247213, 0.5354021, 0.532419, 0.5122666, 
    0.5132139, 0.5165101, 0.5149419, 0.5194255, 0.5205288, 0.5214254, 
    0.5225717, 0.5226954, 0.5233744, 0.5222617, 0.5233305, 0.5192867, 
    0.521094, 0.5161332, 0.517341, 0.5167854, 0.5161759, 0.5180567, 
    0.5200602, 0.5201027, 0.5207451, 0.5225555, 0.5194436, 0.5290699, 
    0.5231269, 0.5142467, 0.5160711, 0.5163314, 0.5156248, 0.5204182, 
    0.5186818, 0.5233579, 0.5220943, 0.5241644, 0.5231358, 0.5229845, 
    0.5216631, 0.5208404, 0.5187615, 0.5170694, 0.5157272, 0.5160393, 
    0.5175136, 0.5201827, 0.5227067, 0.5221539, 0.5240071, 0.5191005, 
    0.5211585, 0.5203632, 0.5224366, 0.5178925, 0.521763, 0.5169029, 
    0.5173291, 0.5186473, 0.5212982, 0.5218842, 0.5225103, 0.5221239, 
    0.5202504, 0.5199433, 0.5186152, 0.5182486, 0.5172363, 0.5163983, 
    0.5171641, 0.5179682, 0.5202511, 0.5223079, 0.5245497, 0.5250981, 
    0.5277171, 0.5255856, 0.529103, 0.5261132, 0.5312877, 0.5219868, 
    0.5260248, 0.5187072, 0.5194958, 0.5209222, 0.5241923, 0.5224268, 
    0.5244914, 0.5199313, 0.5175645, 0.5169517, 0.5158089, 0.5169779, 
    0.5168828, 0.5180013, 0.5176418, 0.5203269, 0.5188847, 0.5229808, 
    0.524475, 0.528693, 0.5312777, 0.5339073, 0.5350681, 0.5354213, 0.535569,
  0.5311409, 0.5336103, 0.53313, 0.5351228, 0.5340171, 0.5353222, 0.5316414, 
    0.5337085, 0.5323887, 0.531363, 0.5389929, 0.5352116, 0.5429236, 
    0.5405093, 0.5465766, 0.5425479, 0.5473894, 0.54646, 0.5492572, 
    0.5484556, 0.552036, 0.5496271, 0.553893, 0.5514605, 0.551841, 0.5495477, 
    0.5359721, 0.5385221, 0.5358211, 0.5361846, 0.5360214, 0.53404, 
    0.5330421, 0.5309521, 0.5313314, 0.5328664, 0.536348, 0.5351657, 
    0.5381457, 0.5380784, 0.5413988, 0.5399013, 0.5454862, 0.543898, 
    0.548489, 0.547334, 0.5484348, 0.5481009, 0.5484391, 0.5467452, 
    0.5474709, 0.5459806, 0.5401818, 0.5418853, 0.5368071, 0.5337572, 
    0.531732, 0.5302957, 0.5304988, 0.5308859, 0.5328754, 0.5347466, 
    0.5361732, 0.5371279, 0.5380687, 0.5409185, 0.5424271, 0.5458076, 
    0.5451971, 0.5462312, 0.5472191, 0.5488785, 0.5486053, 0.5493366, 
    0.5462037, 0.5482857, 0.5448494, 0.545789, 0.5383254, 0.5354846, 
    0.5342785, 0.5332224, 0.5306549, 0.5324278, 0.5317289, 0.5333918, 
    0.5344489, 0.533926, 0.537154, 0.5358987, 0.5425165, 0.5396647, 
    0.5471038, 0.5453224, 0.5475309, 0.5464038, 0.5483354, 0.5465969, 
    0.5496088, 0.550265, 0.5498165, 0.5515392, 0.5465006, 0.5484349, 
    0.5339114, 0.5339966, 0.5343939, 0.532648, 0.5325412, 0.5309417, 
    0.5323648, 0.5329711, 0.5345101, 0.5354209, 0.5362868, 0.5381913, 
    0.5403196, 0.5432973, 0.5454378, 0.5468734, 0.545993, 0.5467702, 
    0.5459014, 0.5454942, 0.5500191, 0.5474778, 0.5512914, 0.5510802, 
    0.5493541, 0.5511041, 0.5340565, 0.5335658, 0.5318628, 0.5331955, 
    0.5307676, 0.5321265, 0.5329082, 0.5359252, 0.5365881, 0.5372033, 
    0.5384182, 0.539978, 0.5427158, 0.5450994, 0.5472765, 0.5471169, 
    0.5471731, 0.5476598, 0.5464547, 0.5478576, 0.5480932, 0.5474774, 
    0.551052, 0.5500304, 0.5510758, 0.5504105, 0.5337253, 0.534551, 
    0.5341048, 0.534944, 0.5343528, 0.5369823, 0.537771, 0.5414633, 
    0.5399473, 0.5423601, 0.5401922, 0.5405763, 0.5424392, 0.5403093, 
    0.5449681, 0.5418093, 0.5476786, 0.5445224, 0.5478765, 0.5472671, 
    0.5482761, 0.5491801, 0.5503175, 0.5524173, 0.5519309, 0.5536875, 
    0.5357823, 0.536854, 0.5367594, 0.5378811, 0.5387109, 0.5405098, 
    0.5433969, 0.542311, 0.5443047, 0.5447052, 0.5416761, 0.5435358, 
    0.5375712, 0.5385344, 0.5379608, 0.5358669, 0.5425614, 0.5391244, 
    0.5454732, 0.5436096, 0.5490512, 0.5463442, 0.5516632, 0.5539398, 
    0.5560829, 0.5585899, 0.5374388, 0.5367104, 0.5380145, 0.5398196, 
    0.5414948, 0.5437232, 0.5439512, 0.5443689, 0.5454508, 0.5463608, 
    0.5445011, 0.546589, 0.5387582, 0.5428598, 0.5364353, 0.538369, 
    0.5397131, 0.5391232, 0.5421868, 0.5429093, 0.5458465, 0.5443277, 
    0.553378, 0.5493713, 0.5604994, 0.5573863, 0.536456, 0.5374362, 
    0.5408494, 0.539225, 0.5438719, 0.5450167, 0.5459474, 0.5471377, 
    0.5472661, 0.5479715, 0.5468157, 0.5479258, 0.5437279, 0.5456033, 
    0.5404589, 0.5417105, 0.5411347, 0.5405031, 0.5424524, 0.5445305, 
    0.5445746, 0.5452412, 0.5471208, 0.5438908, 0.553896, 0.5477144, 
    0.5385052, 0.5403947, 0.5406643, 0.5399323, 0.5449019, 0.5431005, 
    0.5479543, 0.5466419, 0.5487925, 0.5477237, 0.5475665, 0.5461941, 
    0.5453401, 0.5431831, 0.541429, 0.5400383, 0.5403616, 0.5418894, 
    0.5446575, 0.5472779, 0.5467038, 0.548629, 0.5435348, 0.5456702, 
    0.5448449, 0.5469973, 0.5422822, 0.5462978, 0.5412565, 0.5416982, 
    0.5430648, 0.5458153, 0.5464237, 0.5470738, 0.5466726, 0.5447278, 
    0.5444091, 0.5430315, 0.5426514, 0.541602, 0.5407336, 0.5415271, 
    0.5423606, 0.5447285, 0.5468637, 0.549193, 0.5497631, 0.5524875, 0.55027, 
    0.5539305, 0.5508187, 0.5562066, 0.5465303, 0.5507267, 0.5431269, 
    0.5439448, 0.5454251, 0.5488215, 0.5469872, 0.5491323, 0.5443966, 
    0.5419422, 0.5413071, 0.5401229, 0.5413342, 0.5412356, 0.5423949, 
    0.5420223, 0.5448071, 0.543311, 0.5475626, 0.5491154, 0.5535035, 
    0.5561963, 0.5589389, 0.5601506, 0.5605194, 0.5606736,
  0.5352592, 0.5381025, 0.5375492, 0.5398464, 0.5385715, 0.5400766, 0.535835, 
    0.5382156, 0.5366953, 0.5355148, 0.5443176, 0.539949, 0.5488714, 
    0.5460728, 0.5531155, 0.5484356, 0.5540615, 0.55298, 0.5562374, 
    0.5553033, 0.5594807, 0.5566688, 0.5616519, 0.5588084, 0.5592529, 
    0.5565763, 0.5408266, 0.5437729, 0.5406523, 0.541072, 0.5408835, 
    0.5385979, 0.5374479, 0.535042, 0.5354784, 0.5372455, 0.5412607, 
    0.539896, 0.5433377, 0.5432599, 0.5471033, 0.5453688, 0.5518475, 
    0.5500024, 0.5553422, 0.553997, 0.555279, 0.5548901, 0.5552841, 
    0.5533118, 0.5541564, 0.5524224, 0.5456935, 0.5476671, 0.5417908, 
    0.5382718, 0.5359394, 0.5342872, 0.5345206, 0.5349658, 0.5372558, 
    0.5394126, 0.5410588, 0.5421614, 0.5432487, 0.5465468, 0.5482955, 
    0.5522211, 0.5515115, 0.5527138, 0.5538632, 0.5557961, 0.5554777, 
    0.5563301, 0.5526819, 0.5551053, 0.5511075, 0.5521995, 0.5435455, 
    0.540264, 0.5388727, 0.5376556, 0.5347002, 0.5367404, 0.5359358, 
    0.5378507, 0.5390692, 0.5384664, 0.5421916, 0.540742, 0.5483992, 
    0.5450948, 0.5537291, 0.5516571, 0.5542263, 0.5529145, 0.5551632, 
    0.5531392, 0.5566474, 0.5574129, 0.5568898, 0.5589004, 0.5530271, 
    0.5552791, 0.5384496, 0.5385479, 0.5390058, 0.536994, 0.536871, 
    0.5350301, 0.5366679, 0.537366, 0.5391399, 0.5401905, 0.54119, 0.5433905, 
    0.5458531, 0.5493051, 0.5517913, 0.5534609, 0.5524367, 0.5533409, 
    0.5523303, 0.5518568, 0.5571261, 0.5541644, 0.5586109, 0.5583644, 
    0.5563504, 0.5583922, 0.5386169, 0.5380513, 0.5360899, 0.5376246, 
    0.5348298, 0.5363935, 0.5372936, 0.5407725, 0.5415379, 0.5422484, 
    0.5436527, 0.5454575, 0.5486304, 0.551398, 0.5539301, 0.5537444, 
    0.5538098, 0.5543762, 0.5529737, 0.5546067, 0.554881, 0.5541639, 
    0.5583314, 0.5571392, 0.5583591, 0.5575827, 0.5382351, 0.539187, 
    0.5386726, 0.5396402, 0.5389585, 0.5419931, 0.5429045, 0.547178, 
    0.545422, 0.5482177, 0.5457056, 0.5461504, 0.5483094, 0.5458412, 
    0.5512454, 0.5475792, 0.5543983, 0.5507275, 0.5546287, 0.5539191, 
    0.5550941, 0.5561476, 0.5574741, 0.5599262, 0.5593579, 0.5614115, 
    0.5406075, 0.5418449, 0.5417357, 0.5430318, 0.5439913, 0.5460734, 
    0.5494207, 0.5481608, 0.5504747, 0.5509398, 0.5474247, 0.5495819, 
    0.5426736, 0.5437872, 0.5431239, 0.5407052, 0.5484512, 0.5444697, 
    0.5518324, 0.5496675, 0.5559973, 0.5528452, 0.5590452, 0.5617067, 
    0.5642166, 0.5671582, 0.5425206, 0.5416792, 0.5431859, 0.5452742, 
    0.5472146, 0.5497994, 0.5500641, 0.5505492, 0.5518064, 0.5528646, 
    0.5507028, 0.55313, 0.544046, 0.5487974, 0.5413614, 0.5435959, 0.5451509, 
    0.5444683, 0.5480168, 0.5488548, 0.5522664, 0.5505014, 0.5610494, 
    0.5563705, 0.5694026, 0.5657451, 0.5413854, 0.5425176, 0.5464668, 
    0.5445861, 0.5499721, 0.5513018, 0.5523837, 0.5537686, 0.553918, 
    0.5547394, 0.5533938, 0.5546861, 0.5498049, 0.5519837, 0.5460144, 
    0.5474646, 0.5467972, 0.5460657, 0.5483248, 0.5507368, 0.5507881, 
    0.5515627, 0.5537488, 0.549994, 0.5616553, 0.5544399, 0.5437534, 0.54594, 
    0.5462523, 0.5454046, 0.5511684, 0.5490767, 0.5547193, 0.5531915, 
    0.5556958, 0.5544508, 0.5542676, 0.5526707, 0.5516777, 0.5491726, 
    0.5471383, 0.5455275, 0.5459018, 0.5476719, 0.5508845, 0.5539317, 
    0.5532635, 0.5555053, 0.5495808, 0.5520614, 0.5511021, 0.5536051, 
    0.5481274, 0.5527913, 0.5469384, 0.5474503, 0.5490353, 0.5522301, 
    0.5529377, 0.5536942, 0.5532272, 0.5509661, 0.5505959, 0.5489966, 
    0.5485556, 0.5473388, 0.5463325, 0.5472519, 0.5482184, 0.5509669, 
    0.5534497, 0.5561627, 0.5568274, 0.5600083, 0.5574187, 0.5616957, 
    0.558059, 0.5643616, 0.5530617, 0.5579516, 0.5491073, 0.5500568, 
    0.5517764, 0.5557296, 0.5535934, 0.556092, 0.5505814, 0.5477332, 
    0.546997, 0.5456254, 0.5470284, 0.5469142, 0.5482582, 0.5478261, 
    0.5510583, 0.549321, 0.5542632, 0.5560721, 0.5611962, 0.5643494, 
    0.5675681, 0.5689924, 0.5694262, 0.5696077,
  0.5840976, 0.5875086, 0.5868437, 0.5896073, 0.5880725, 0.5898846, 
    0.5847872, 0.5876446, 0.5858188, 0.5844036, 0.5950114, 0.5897309, 
    0.6005509, 0.5971422, 0.6057471, 0.6000192, 0.6069097, 0.6055806, 
    0.6095905, 0.6084385, 0.613603, 0.610123, 0.6163005, 0.6127695, 
    0.6133204, 0.6100087, 0.5907891, 0.5943512, 0.5905789, 0.5910851, 
    0.5908578, 0.5881042, 0.5867221, 0.5838375, 0.58436, 0.5864791, 
    0.5913129, 0.589667, 0.5938241, 0.5937299, 0.5983957, 0.596287, 
    0.6041912, 0.6019324, 0.6084865, 0.6068304, 0.6084087, 0.6079295, 
    0.6084149, 0.6059882, 0.6070265, 0.6048962, 0.5966813, 0.5990824, 
    0.5919532, 0.5877121, 0.5849124, 0.5829344, 0.5832136, 0.5837463, 
    0.5864915, 0.5890847, 0.5910693, 0.5924011, 0.5937164, 0.5977185, 
    0.5998483, 0.6046493, 0.6037793, 0.6052538, 0.6066659, 0.609046, 
    0.6086535, 0.6097049, 0.6052146, 0.6081945, 0.6032844, 0.6046228, 
    0.5940757, 0.5901105, 0.5884349, 0.5869715, 0.5834284, 0.5858728, 
    0.5849079, 0.587206, 0.5886714, 0.5879461, 0.5924375, 0.590687, 
    0.5999748, 0.5959544, 0.606501, 0.6039577, 0.6071125, 0.6055002, 
    0.6082659, 0.6057761, 0.6100966, 0.6110424, 0.6103959, 0.6128834, 
    0.6056384, 0.6084088, 0.5879259, 0.588044, 0.5885951, 0.5861772, 
    0.5860295, 0.5838232, 0.5857859, 0.5866238, 0.5887564, 0.5900219, 
    0.5912276, 0.593888, 0.5968752, 0.6010804, 0.6041222, 0.6061714, 
    0.6049138, 0.6060239, 0.6047831, 0.6042026, 0.6106879, 0.6070363, 
    0.6125249, 0.6122196, 0.6097299, 0.612254, 0.5881271, 0.587447, 
    0.5850927, 0.5869343, 0.5835835, 0.5854568, 0.5865368, 0.5907238, 
    0.5916477, 0.5925063, 0.5942057, 0.5963947, 0.6002568, 0.6036403, 
    0.6067482, 0.6065198, 0.6066002, 0.6072969, 0.6055729, 0.6075805, 
    0.6079184, 0.6070357, 0.6121787, 0.6107041, 0.6122131, 0.6112524, 
    0.5876679, 0.5888132, 0.5881941, 0.5893589, 0.5885381, 0.5921977, 
    0.5932998, 0.5984868, 0.5963516, 0.5997534, 0.5966961, 0.5972366, 
    0.5998653, 0.5968608, 0.6034534, 0.5989752, 0.6073241, 0.6028193, 
    0.6076077, 0.6067347, 0.6081808, 0.6094796, 0.6111181, 0.6141557, 
    0.6134506, 0.6160014, 0.5905248, 0.5920186, 0.5918867, 0.5934538, 
    0.5946159, 0.5971429, 0.6012216, 0.5996841, 0.60251, 0.6030792, 
    0.5987871, 0.6014184, 0.5930204, 0.5943686, 0.5935653, 0.5906426, 
    0.6000383, 0.5951958, 0.6041727, 0.601523, 0.6092943, 0.6054151, 
    0.613063, 0.6163687, 0.619499, 0.623184, 0.5928354, 0.5918184, 0.5936404, 
    0.5961721, 0.5985312, 0.6016843, 0.6020079, 0.6026012, 0.6041408, 
    0.6054389, 0.6027891, 0.6057648, 0.5946822, 0.6004606, 0.5914346, 
    0.5941368, 0.5960224, 0.5951942, 0.5995085, 0.6005306, 0.6047048, 
    0.6025427, 0.615551, 0.6097547, 0.6260078, 0.6214116, 0.5914636, 
    0.5928317, 0.5976212, 0.595337, 0.6018954, 0.6035225, 0.6048487, 
    0.6065495, 0.6067333, 0.607744, 0.6060889, 0.6076784, 0.6016911, 
    0.6043581, 0.5970713, 0.5988357, 0.5980232, 0.5971336, 0.5998841, 
    0.6028308, 0.6028935, 0.6038421, 0.6065252, 0.6019221, 0.6163048, 
    0.6073753, 0.5943276, 0.5969808, 0.5973604, 0.5963304, 0.6033591, 
    0.6008015, 0.6077192, 0.6058404, 0.6089224, 0.6073886, 0.6071634, 
    0.6052009, 0.603983, 0.6009186, 0.5984383, 0.5964796, 0.5969344, 
    0.5990883, 0.6030115, 0.6067501, 0.6059289, 0.6086875, 0.6014171, 
    0.6044534, 0.6032779, 0.6063486, 0.5996433, 0.6053489, 0.598195, 
    0.5988182, 0.6007509, 0.6046603, 0.6055287, 0.6064581, 0.6058843, 
    0.6031114, 0.6026583, 0.6007037, 0.6001655, 0.5986825, 0.5974579, 
    0.5985767, 0.5997543, 0.6031124, 0.6061576, 0.6094982, 0.6103189, 
    0.6142576, 0.6110495, 0.6163551, 0.6118417, 0.6196803, 0.6056809, 
    0.6117087, 0.6008388, 0.6019989, 0.604104, 0.6089641, 0.6063341, 
    0.609411, 0.6026406, 0.5991629, 0.5982664, 0.5965986, 0.5983046, 
    0.5981656, 0.5998029, 0.5992761, 0.6032243, 0.6010998, 0.6071578, 
    0.6093865, 0.6157336, 0.6196651, 0.623699, 0.6254908, 0.6260375, 0.6262662,
  0.6622251, 0.667787, 0.6666976, 0.6712429, 0.6687129, 0.6717016, 0.6633443, 
    0.6680101, 0.6650231, 0.6627214, 0.6802661, 0.6714472, 0.6897115, 
    0.6838751, 0.6987642, 0.6887959, 0.7008165, 0.6984711, 0.7055877, 
    0.7035307, 0.7128337, 0.7065421, 0.7177787, 0.711318, 0.7123192, 
    0.706337, 0.6732006, 0.679154, 0.6728517, 0.6736924, 0.6733148, 
    0.6687651, 0.6664985, 0.6618038, 0.6626507, 0.6661011, 0.6740712, 
    0.6713416, 0.6782681, 0.6781098, 0.6860123, 0.682423, 0.6960332, 
    0.6920996, 0.7036162, 0.7006762, 0.7034775, 0.7026251, 0.7034886, 
    0.6991889, 0.7010233, 0.6972684, 0.683092, 0.6871875, 0.6751375, 
    0.6681209, 0.6635476, 0.6603438, 0.6607947, 0.6616562, 0.6661214, 
    0.6703799, 0.6736662, 0.6758848, 0.6780871, 0.6848564, 0.688502, 
    0.6968355, 0.6953132, 0.6978964, 0.7003853, 0.7046142, 0.7039137, 
    0.7057924, 0.6978275, 0.7030964, 0.6944497, 0.696789, 0.6786907, 
    0.6720755, 0.669309, 0.6669068, 0.6611419, 0.6651114, 0.6635405, 
    0.6672908, 0.6696985, 0.6685052, 0.6759457, 0.6730312, 0.6887196, 
    0.6818596, 0.7000939, 0.6956249, 0.7011755, 0.6983296, 0.7032234, 
    0.6988153, 0.7064946, 0.7081949, 0.707032, 0.7115249, 0.6985729, 
    0.7034777, 0.6684719, 0.6686662, 0.6695728, 0.665608, 0.665367, 
    0.6617807, 0.6649695, 0.6663378, 0.6698384, 0.6719288, 0.6739292, 
    0.6783753, 0.6834213, 0.6906251, 0.6959125, 0.6995119, 0.6972994, 
    0.6992519, 0.6970701, 0.6960531, 0.7075568, 0.7010406, 0.7108743, 
    0.710321, 0.7058374, 0.7103833, 0.6688027, 0.6676859, 0.6638409, 
    0.6668458, 0.6613927, 0.6644333, 0.6661956, 0.6730922, 0.6746284, 
    0.6760606, 0.6789091, 0.6826057, 0.6892048, 0.6950704, 0.7005307, 
    0.7001271, 0.7002691, 0.7015024, 0.6984575, 0.7020053, 0.7026053, 
    0.7010396, 0.710247, 0.7075859, 0.7103093, 0.7085733, 0.6680484, 
    0.6699321, 0.6689128, 0.6708325, 0.6694789, 0.6755454, 0.6773884, 
    0.6861679, 0.6825325, 0.6883391, 0.683117, 0.6840357, 0.6885313, 
    0.6833967, 0.6947443, 0.6870038, 0.7015504, 0.6936398, 0.7020535, 
    0.7005069, 0.703072, 0.7053893, 0.7083312, 0.713842, 0.7125562, 
    0.7172273, 0.672762, 0.6752465, 0.6750265, 0.6776467, 0.6795995, 
    0.6838763, 0.6908692, 0.6882198, 0.6931019, 0.6940922, 0.6866817, 
    0.6912096, 0.6769205, 0.6791831, 0.6778337, 0.6729575, 0.6888287, 
    0.6805774, 0.6960008, 0.6913906, 0.7050577, 0.69818, 0.711851, 0.7179045, 
    0.7237219, 0.7306815, 0.6766108, 0.6749127, 0.6779597, 0.6822283, 
    0.6862438, 0.6916698, 0.6922304, 0.6932604, 0.6959449, 0.6982217, 
    0.6935872, 0.6987953, 0.6797112, 0.6895558, 0.6742736, 0.6787933, 
    0.6819748, 0.6805746, 0.6879184, 0.6896765, 0.6969327, 0.6931587, 
    0.7163987, 0.7058818, 0.7360995, 0.7273188, 0.6743218, 0.6766047, 
    0.6846905, 0.6808156, 0.6920354, 0.6948648, 0.6971852, 0.7001796, 
    0.7005044, 0.7022954, 0.6993665, 0.702179, 0.6916814, 0.6963252, 
    0.6837546, 0.6867649, 0.685376, 0.6838604, 0.6885635, 0.6936597, 
    0.6937689, 0.6954229, 0.7001367, 0.6920817, 0.7177866, 0.7016412, 
    0.6791143, 0.6836007, 0.6842464, 0.6824967, 0.6945799, 0.6901437, 
    0.7022516, 0.6989285, 0.7043934, 0.7016648, 0.7012656, 0.6978035, 
    0.6956691, 0.6903458, 0.6860851, 0.6827497, 0.6835218, 0.6871974, 
    0.6939742, 0.7005342, 0.6990844, 0.7039744, 0.6912072, 0.6964923, 
    0.6944383, 0.6998248, 0.6881498, 0.6980637, 0.6856694, 0.686735, 
    0.6900563, 0.6968548, 0.6983797, 0.7000182, 0.6990059, 0.6941482, 
    0.6933598, 0.689975, 0.6890477, 0.6865026, 0.6844125, 0.6863217, 
    0.6883404, 0.6941499, 0.6994876, 0.7054225, 0.7068936, 0.7140281, 
    0.7082077, 0.7178792, 0.7096372, 0.7240614, 0.6986477, 0.709397, 
    0.6902081, 0.6922148, 0.6958807, 0.7044679, 0.6997992, 0.7052665, 
    0.6933289, 0.6873254, 0.6857913, 0.6829515, 0.6858565, 0.6856191, 
    0.6884239, 0.6875196, 0.6943448, 0.6906587, 0.7012558, 0.7052227, 
    0.7167343, 0.7240329, 0.731664, 0.7351019, 0.7361569, 0.7365991,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.506774e-11, 3.522342e-11, 3.519307e-11, 3.531871e-11, 3.524898e-11, 
    3.533118e-11, 3.509911e-11, 3.522932e-11, 3.514615e-11, 3.508145e-11, 
    3.556242e-11, 3.532402e-11, 3.581065e-11, 3.565821e-11, 3.604128e-11, 
    3.578679e-11, 3.609261e-11, 3.603389e-11, 3.621064e-11, 3.615992e-11, 
    3.638605e-11, 3.623392e-11, 3.650343e-11, 3.634967e-11, 3.637364e-11, 
    3.622871e-11, 3.537228e-11, 3.553298e-11, 3.536268e-11, 3.53856e-11, 
    3.537528e-11, 3.525023e-11, 3.518724e-11, 3.505553e-11, 3.507938e-11, 
    3.517611e-11, 3.539562e-11, 3.532103e-11, 3.5509e-11, 3.550476e-11, 
    3.571422e-11, 3.561971e-11, 3.597232e-11, 3.587197e-11, 3.616199e-11, 
    3.608893e-11, 3.615848e-11, 3.613733e-11, 3.615864e-11, 3.605161e-11, 
    3.609737e-11, 3.600324e-11, 3.563785e-11, 3.574532e-11, 3.54248e-11, 
    3.523227e-11, 3.510466e-11, 3.501417e-11, 3.502687e-11, 3.505125e-11, 
    3.517659e-11, 3.529457e-11, 3.538455e-11, 3.544472e-11, 3.550403e-11, 
    3.568374e-11, 3.577902e-11, 3.59925e-11, 3.595397e-11, 3.601919e-11, 
    3.608163e-11, 3.618642e-11, 3.616915e-11, 3.621529e-11, 3.60173e-11, 
    3.614882e-11, 3.593168e-11, 3.599102e-11, 3.552038e-11, 3.534131e-11, 
    3.526512e-11, 3.519855e-11, 3.503667e-11, 3.514841e-11, 3.51043e-11, 
    3.520912e-11, 3.527575e-11, 3.524273e-11, 3.544632e-11, 3.536706e-11, 
    3.57846e-11, 3.560461e-11, 3.60744e-11, 3.596179e-11, 3.610128e-11, 
    3.603008e-11, 3.615201e-11, 3.60422e-11, 3.623242e-11, 3.627388e-11, 
    3.624546e-11, 3.635438e-11, 3.603587e-11, 3.615807e-11, 3.524202e-11, 
    3.524741e-11, 3.527242e-11, 3.516222e-11, 3.515548e-11, 3.505463e-11, 
    3.514428e-11, 3.518249e-11, 3.527953e-11, 3.533689e-11, 3.539146e-11, 
    3.551163e-11, 3.564585e-11, 3.583381e-11, 3.596904e-11, 3.605969e-11, 
    3.600405e-11, 3.605309e-11, 3.599818e-11, 3.597241e-11, 3.625822e-11, 
    3.609764e-11, 3.63386e-11, 3.632527e-11, 3.621608e-11, 3.632666e-11, 
    3.52511e-11, 3.522012e-11, 3.511271e-11, 3.519669e-11, 3.504359e-11, 
    3.512922e-11, 3.517842e-11, 3.536862e-11, 3.541045e-11, 3.544925e-11, 
    3.552588e-11, 3.562425e-11, 3.579706e-11, 3.594755e-11, 3.608512e-11, 
    3.607498e-11, 3.60785e-11, 3.610917e-11, 3.603302e-11, 3.61216e-11, 
    3.613642e-11, 3.609754e-11, 3.632336e-11, 3.62588e-11, 3.632483e-11, 
    3.628273e-11, 3.523013e-11, 3.528213e-11, 3.525395e-11, 3.530685e-11, 
    3.526949e-11, 3.54353e-11, 3.5485e-11, 3.571799e-11, 3.56223e-11, 
    3.577461e-11, 3.56377e-11, 3.566194e-11, 3.577937e-11, 3.5645e-11, 
    3.593909e-11, 3.573951e-11, 3.611033e-11, 3.591074e-11, 3.612276e-11, 
    3.608421e-11, 3.614791e-11, 3.620502e-11, 3.627683e-11, 3.640953e-11, 
    3.637872e-11, 3.648978e-11, 3.535975e-11, 3.542725e-11, 3.542132e-11, 
    3.549203e-11, 3.554432e-11, 3.565789e-11, 3.584011e-11, 3.57715e-11, 
    3.589736e-11, 3.592265e-11, 3.57313e-11, 3.584868e-11, 3.547212e-11, 
    3.553279e-11, 3.549664e-11, 3.536446e-11, 3.578692e-11, 3.556988e-11, 
    3.59708e-11, 3.585303e-11, 3.619676e-11, 3.602567e-11, 3.636177e-11, 
    3.65056e-11, 3.664118e-11, 3.679955e-11, 3.546414e-11, 3.541815e-11, 
    3.550037e-11, 3.561423e-11, 3.571994e-11, 3.586067e-11, 3.587504e-11, 
    3.590135e-11, 3.596966e-11, 3.602715e-11, 3.590956e-11, 3.604145e-11, 
    3.554676e-11, 3.580578e-11, 3.540025e-11, 3.55222e-11, 3.560699e-11, 
    3.556979e-11, 3.576317e-11, 3.580872e-11, 3.599414e-11, 3.589827e-11, 
    3.646994e-11, 3.621674e-11, 3.692032e-11, 3.672338e-11, 3.540205e-11, 
    3.546383e-11, 3.567914e-11, 3.557665e-11, 3.586997e-11, 3.594227e-11, 
    3.6001e-11, 3.607617e-11, 3.608423e-11, 3.61288e-11, 3.60557e-11, 
    3.612585e-11, 3.586055e-11, 3.597903e-11, 3.565413e-11, 3.573306e-11, 
    3.569671e-11, 3.565679e-11, 3.57798e-11, 3.591096e-11, 3.591378e-11, 
    3.595578e-11, 3.607427e-11, 3.587045e-11, 3.650239e-11, 3.611167e-11, 
    3.553124e-11, 3.565034e-11, 3.566739e-11, 3.562121e-11, 3.593491e-11, 
    3.582114e-11, 3.612772e-11, 3.604474e-11, 3.618058e-11, 3.611305e-11, 
    3.610302e-11, 3.601634e-11, 3.596229e-11, 3.582604e-11, 3.571519e-11, 
    3.562746e-11, 3.564778e-11, 3.574419e-11, 3.591889e-11, 3.608447e-11, 
    3.604812e-11, 3.616977e-11, 3.584789e-11, 3.598274e-11, 3.59305e-11, 
    3.606653e-11, 3.576951e-11, 3.602293e-11, 3.570473e-11, 3.573255e-11, 
    3.581877e-11, 3.599243e-11, 3.603088e-11, 3.607193e-11, 3.604653e-11, 
    3.592363e-11, 3.590347e-11, 3.581643e-11, 3.579235e-11, 3.572614e-11, 
    3.567123e-11, 3.572131e-11, 3.577382e-11, 3.59234e-11, 3.605822e-11, 
    3.620534e-11, 3.624139e-11, 3.641335e-11, 3.627321e-11, 3.650437e-11, 
    3.630763e-11, 3.664831e-11, 3.60376e-11, 3.630276e-11, 3.582273e-11, 
    3.587432e-11, 3.596772e-11, 3.618223e-11, 3.606637e-11, 3.620185e-11, 
    3.590267e-11, 3.574755e-11, 3.570748e-11, 3.563273e-11, 3.570911e-11, 
    3.57029e-11, 3.577605e-11, 3.575247e-11, 3.592825e-11, 3.583379e-11, 
    3.610224e-11, 3.620034e-11, 3.647767e-11, 3.664783e-11, 3.682134e-11, 
    3.689792e-11, 3.692124e-11, 3.693094e-11,
  1.781549e-11, 1.79512e-11, 1.79248e-11, 1.803447e-11, 1.797361e-11, 
    1.804547e-11, 1.784298e-11, 1.795659e-11, 1.788404e-11, 1.78277e-11, 
    1.824801e-11, 1.803938e-11, 1.846581e-11, 1.833202e-11, 1.866883e-11, 
    1.844495e-11, 1.87141e-11, 1.866239e-11, 1.881827e-11, 1.877357e-11, 
    1.897341e-11, 1.883892e-11, 1.907735e-11, 1.894127e-11, 1.896253e-11, 
    1.883448e-11, 1.808132e-11, 1.822198e-11, 1.807299e-11, 1.809302e-11, 
    1.808404e-11, 1.797486e-11, 1.791992e-11, 1.780515e-11, 1.782597e-11, 
    1.791028e-11, 1.810203e-11, 1.803687e-11, 1.820131e-11, 1.819759e-11, 
    1.83813e-11, 1.829838e-11, 1.860821e-11, 1.851996e-11, 1.877543e-11, 
    1.871106e-11, 1.87724e-11, 1.87538e-11, 1.877264e-11, 1.867827e-11, 
    1.871868e-11, 1.863572e-11, 1.83139e-11, 1.840825e-11, 1.812737e-11, 
    1.795923e-11, 1.784795e-11, 1.776913e-11, 1.778027e-11, 1.780149e-11, 
    1.791078e-11, 1.801378e-11, 1.809242e-11, 1.81451e-11, 1.819706e-11, 
    1.835461e-11, 1.843827e-11, 1.862606e-11, 1.859214e-11, 1.864964e-11, 
    1.870466e-11, 1.879714e-11, 1.878191e-11, 1.882269e-11, 1.864814e-11, 
    1.876407e-11, 1.857283e-11, 1.862506e-11, 1.82111e-11, 1.805445e-11, 
    1.798794e-11, 1.792987e-11, 1.778883e-11, 1.788618e-11, 1.784777e-11, 
    1.793921e-11, 1.799738e-11, 1.796861e-11, 1.814654e-11, 1.807728e-11, 
    1.844323e-11, 1.828526e-11, 1.869824e-11, 1.85991e-11, 1.872203e-11, 
    1.865927e-11, 1.876685e-11, 1.867002e-11, 1.883788e-11, 1.88745e-11, 
    1.884947e-11, 1.89457e-11, 1.866466e-11, 1.877239e-11, 1.79678e-11, 
    1.797249e-11, 1.799436e-11, 1.789828e-11, 1.789241e-11, 1.780457e-11, 
    1.788273e-11, 1.791605e-11, 1.800077e-11, 1.805093e-11, 1.809868e-11, 
    1.820382e-11, 1.83215e-11, 1.848657e-11, 1.860553e-11, 1.868541e-11, 
    1.863642e-11, 1.867967e-11, 1.863132e-11, 1.860868e-11, 1.886077e-11, 
    1.871905e-11, 1.893185e-11, 1.892005e-11, 1.882365e-11, 1.892138e-11, 
    1.797578e-11, 1.794879e-11, 1.785514e-11, 1.792841e-11, 1.779502e-11, 
    1.786963e-11, 1.791257e-11, 1.807871e-11, 1.811531e-11, 1.814924e-11, 
    1.821636e-11, 1.830262e-11, 1.845431e-11, 1.858669e-11, 1.870787e-11, 
    1.869898e-11, 1.870211e-11, 1.87292e-11, 1.86621e-11, 1.874023e-11, 
    1.875334e-11, 1.871905e-11, 1.891847e-11, 1.886142e-11, 1.89198e-11, 
    1.888265e-11, 1.795756e-11, 1.800301e-11, 1.797845e-11, 1.802465e-11, 
    1.799209e-11, 1.813701e-11, 1.818055e-11, 1.838484e-11, 1.830092e-11, 
    1.843457e-11, 1.831449e-11, 1.833574e-11, 1.843889e-11, 1.832097e-11, 
    1.857937e-11, 1.8404e-11, 1.873026e-11, 1.855456e-11, 1.874128e-11, 
    1.870734e-11, 1.876356e-11, 1.881396e-11, 1.887745e-11, 1.899477e-11, 
    1.896758e-11, 1.906587e-11, 1.807086e-11, 1.812995e-11, 1.812476e-11, 
    1.818669e-11, 1.823253e-11, 1.833207e-11, 1.849212e-11, 1.843188e-11, 
    1.854255e-11, 1.85648e-11, 1.839669e-11, 1.849982e-11, 1.816955e-11, 
    1.822274e-11, 1.819108e-11, 1.807551e-11, 1.844573e-11, 1.825536e-11, 
    1.860749e-11, 1.850393e-11, 1.880677e-11, 1.865591e-11, 1.895262e-11, 
    1.907994e-11, 1.920013e-11, 1.934084e-11, 1.816225e-11, 1.812206e-11, 
    1.819406e-11, 1.829382e-11, 1.838662e-11, 1.851024e-11, 1.852291e-11, 
    1.854611e-11, 1.860626e-11, 1.865688e-11, 1.855343e-11, 1.866958e-11, 
    1.823505e-11, 1.84623e-11, 1.810686e-11, 1.821359e-11, 1.828794e-11, 
    1.825533e-11, 1.8425e-11, 1.846507e-11, 1.862823e-11, 1.854383e-11, 
    1.904847e-11, 1.882458e-11, 1.944829e-11, 1.927324e-11, 1.810802e-11, 
    1.816212e-11, 1.835085e-11, 1.826096e-11, 1.851851e-11, 1.858211e-11, 
    1.863388e-11, 1.870011e-11, 1.870728e-11, 1.874657e-11, 1.86822e-11, 
    1.874404e-11, 1.85105e-11, 1.861473e-11, 1.832926e-11, 1.839858e-11, 
    1.836668e-11, 1.833171e-11, 1.843973e-11, 1.855505e-11, 1.855754e-11, 
    1.859458e-11, 1.869902e-11, 1.851956e-11, 1.907738e-11, 1.873211e-11, 
    1.822118e-11, 1.832564e-11, 1.834062e-11, 1.83001e-11, 1.857573e-11, 
    1.847568e-11, 1.874562e-11, 1.867253e-11, 1.879235e-11, 1.873277e-11, 
    1.872401e-11, 1.864761e-11, 1.860009e-11, 1.848025e-11, 1.838297e-11, 
    1.830598e-11, 1.832387e-11, 1.840848e-11, 1.856212e-11, 1.870792e-11, 
    1.867594e-11, 1.878324e-11, 1.849979e-11, 1.861843e-11, 1.857253e-11, 
    1.869231e-11, 1.843027e-11, 1.865323e-11, 1.837344e-11, 1.839791e-11, 
    1.847369e-11, 1.862647e-11, 1.866038e-11, 1.869656e-11, 1.867424e-11, 
    1.856603e-11, 1.854834e-11, 1.847186e-11, 1.845075e-11, 1.839258e-11, 
    1.834447e-11, 1.838842e-11, 1.843461e-11, 1.856609e-11, 1.868485e-11, 
    1.881467e-11, 1.88465e-11, 1.899862e-11, 1.887471e-11, 1.90793e-11, 
    1.890525e-11, 1.920694e-11, 1.866623e-11, 1.89002e-11, 1.847715e-11, 
    1.852256e-11, 1.860478e-11, 1.879391e-11, 1.869174e-11, 1.881126e-11, 
    1.854765e-11, 1.841139e-11, 1.837624e-11, 1.831065e-11, 1.837774e-11, 
    1.837228e-11, 1.843655e-11, 1.841589e-11, 1.857046e-11, 1.848737e-11, 
    1.872378e-11, 1.881032e-11, 1.905555e-11, 1.920644e-11, 1.936053e-11, 
    1.942868e-11, 1.944944e-11, 1.945812e-11,
  1.677788e-11, 1.692675e-11, 1.689777e-11, 1.701816e-11, 1.695133e-11, 
    1.703023e-11, 1.680802e-11, 1.693266e-11, 1.685305e-11, 1.679126e-11, 
    1.725282e-11, 1.702354e-11, 1.749245e-11, 1.734519e-11, 1.771615e-11, 
    1.746949e-11, 1.776607e-11, 1.770903e-11, 1.788097e-11, 1.783165e-11, 
    1.80523e-11, 1.790376e-11, 1.816716e-11, 1.801679e-11, 1.804027e-11, 
    1.789887e-11, 1.706959e-11, 1.72242e-11, 1.706045e-11, 1.708245e-11, 
    1.707258e-11, 1.695271e-11, 1.689243e-11, 1.676653e-11, 1.678936e-11, 
    1.688185e-11, 1.709235e-11, 1.702078e-11, 1.720144e-11, 1.719735e-11, 
    1.739941e-11, 1.730818e-11, 1.764931e-11, 1.755207e-11, 1.78337e-11, 
    1.776269e-11, 1.783036e-11, 1.780984e-11, 1.783063e-11, 1.772654e-11, 
    1.77711e-11, 1.767963e-11, 1.732524e-11, 1.742907e-11, 1.712019e-11, 
    1.693558e-11, 1.681347e-11, 1.672705e-11, 1.673926e-11, 1.676253e-11, 
    1.688239e-11, 1.699543e-11, 1.708179e-11, 1.713966e-11, 1.719676e-11, 
    1.737006e-11, 1.746213e-11, 1.766899e-11, 1.76316e-11, 1.769498e-11, 
    1.775564e-11, 1.785766e-11, 1.784085e-11, 1.788585e-11, 1.769332e-11, 
    1.782117e-11, 1.761031e-11, 1.766787e-11, 1.721224e-11, 1.704008e-11, 
    1.696708e-11, 1.690333e-11, 1.674864e-11, 1.68554e-11, 1.681328e-11, 
    1.691357e-11, 1.697743e-11, 1.694584e-11, 1.714124e-11, 1.706516e-11, 
    1.746759e-11, 1.729376e-11, 1.774856e-11, 1.763927e-11, 1.77748e-11, 
    1.770559e-11, 1.782424e-11, 1.771744e-11, 1.790262e-11, 1.794305e-11, 
    1.791542e-11, 1.802167e-11, 1.771153e-11, 1.783036e-11, 1.694495e-11, 
    1.69501e-11, 1.697411e-11, 1.686868e-11, 1.686224e-11, 1.67659e-11, 
    1.685162e-11, 1.688817e-11, 1.698114e-11, 1.703622e-11, 1.708866e-11, 
    1.72042e-11, 1.733362e-11, 1.751531e-11, 1.764635e-11, 1.773441e-11, 
    1.768039e-11, 1.772808e-11, 1.767477e-11, 1.764981e-11, 1.792789e-11, 
    1.777152e-11, 1.800637e-11, 1.799334e-11, 1.788692e-11, 1.799481e-11, 
    1.695372e-11, 1.692409e-11, 1.682136e-11, 1.690173e-11, 1.675543e-11, 
    1.683724e-11, 1.688436e-11, 1.706673e-11, 1.710693e-11, 1.714422e-11, 
    1.721798e-11, 1.731284e-11, 1.747978e-11, 1.76256e-11, 1.775917e-11, 
    1.774937e-11, 1.775282e-11, 1.778271e-11, 1.770871e-11, 1.779487e-11, 
    1.780934e-11, 1.77715e-11, 1.79916e-11, 1.79286e-11, 1.799307e-11, 
    1.795204e-11, 1.693372e-11, 1.698361e-11, 1.695664e-11, 1.700736e-11, 
    1.697162e-11, 1.713079e-11, 1.717864e-11, 1.740331e-11, 1.731097e-11, 
    1.745805e-11, 1.732589e-11, 1.734927e-11, 1.746283e-11, 1.733302e-11, 
    1.761753e-11, 1.742441e-11, 1.778387e-11, 1.759021e-11, 1.779603e-11, 
    1.775859e-11, 1.782061e-11, 1.787622e-11, 1.79463e-11, 1.807589e-11, 
    1.804585e-11, 1.815446e-11, 1.70581e-11, 1.712302e-11, 1.711731e-11, 
    1.718536e-11, 1.723576e-11, 1.734523e-11, 1.752141e-11, 1.745508e-11, 
    1.757696e-11, 1.760146e-11, 1.741634e-11, 1.752989e-11, 1.716654e-11, 
    1.722501e-11, 1.719019e-11, 1.706321e-11, 1.747034e-11, 1.726088e-11, 
    1.764851e-11, 1.753442e-11, 1.786828e-11, 1.77019e-11, 1.802932e-11, 
    1.817002e-11, 1.830293e-11, 1.845869e-11, 1.715851e-11, 1.711435e-11, 
    1.719347e-11, 1.730317e-11, 1.740526e-11, 1.754136e-11, 1.755532e-11, 
    1.758088e-11, 1.764715e-11, 1.770295e-11, 1.758895e-11, 1.771695e-11, 
    1.723856e-11, 1.748857e-11, 1.709765e-11, 1.721495e-11, 1.72967e-11, 
    1.726083e-11, 1.744751e-11, 1.749162e-11, 1.767138e-11, 1.757837e-11, 
    1.813524e-11, 1.788796e-11, 1.85777e-11, 1.838384e-11, 1.709892e-11, 
    1.715836e-11, 1.73659e-11, 1.726702e-11, 1.755047e-11, 1.762054e-11, 
    1.76776e-11, 1.775063e-11, 1.775853e-11, 1.780187e-11, 1.773087e-11, 
    1.779907e-11, 1.754166e-11, 1.765649e-11, 1.734214e-11, 1.741842e-11, 
    1.738332e-11, 1.734483e-11, 1.746372e-11, 1.759074e-11, 1.759347e-11, 
    1.763428e-11, 1.774947e-11, 1.755163e-11, 1.816723e-11, 1.778596e-11, 
    1.722328e-11, 1.733818e-11, 1.735464e-11, 1.731007e-11, 1.761351e-11, 
    1.75033e-11, 1.780082e-11, 1.77202e-11, 1.785237e-11, 1.778664e-11, 
    1.777698e-11, 1.769273e-11, 1.764036e-11, 1.750834e-11, 1.740125e-11, 
    1.731653e-11, 1.733622e-11, 1.742933e-11, 1.759852e-11, 1.775924e-11, 
    1.772398e-11, 1.784231e-11, 1.752985e-11, 1.766058e-11, 1.761e-11, 
    1.774202e-11, 1.745331e-11, 1.769898e-11, 1.739075e-11, 1.741768e-11, 
    1.750112e-11, 1.766945e-11, 1.770681e-11, 1.774671e-11, 1.772209e-11, 
    1.760283e-11, 1.758333e-11, 1.749909e-11, 1.747585e-11, 1.741182e-11, 
    1.735887e-11, 1.740724e-11, 1.745809e-11, 1.760289e-11, 1.77338e-11, 
    1.787701e-11, 1.791214e-11, 1.808017e-11, 1.794331e-11, 1.816936e-11, 
    1.797706e-11, 1.83105e-11, 1.771329e-11, 1.797145e-11, 1.750492e-11, 
    1.755493e-11, 1.764553e-11, 1.785411e-11, 1.77414e-11, 1.787325e-11, 
    1.758257e-11, 1.743254e-11, 1.739383e-11, 1.732167e-11, 1.739548e-11, 
    1.738947e-11, 1.746021e-11, 1.743747e-11, 1.760771e-11, 1.751617e-11, 
    1.777673e-11, 1.787221e-11, 1.814305e-11, 1.830992e-11, 1.848047e-11, 
    1.855596e-11, 1.857897e-11, 1.858859e-11,
  1.721998e-11, 1.738378e-11, 1.735188e-11, 1.748443e-11, 1.741085e-11, 
    1.749772e-11, 1.725313e-11, 1.73903e-11, 1.730267e-11, 1.72347e-11, 
    1.774304e-11, 1.749035e-11, 1.80074e-11, 1.784488e-11, 1.825451e-11, 
    1.798206e-11, 1.830969e-11, 1.824663e-11, 1.843675e-11, 1.838219e-11, 
    1.862639e-11, 1.846196e-11, 1.87536e-11, 1.858707e-11, 1.861307e-11, 
    1.845655e-11, 1.754107e-11, 1.771148e-11, 1.7531e-11, 1.755524e-11, 
    1.754436e-11, 1.741236e-11, 1.734602e-11, 1.72075e-11, 1.723261e-11, 
    1.733437e-11, 1.756615e-11, 1.748731e-11, 1.768635e-11, 1.768185e-11, 
    1.79047e-11, 1.780405e-11, 1.818063e-11, 1.807321e-11, 1.838447e-11, 
    1.830595e-11, 1.838077e-11, 1.835807e-11, 1.838107e-11, 1.826598e-11, 
    1.831525e-11, 1.821413e-11, 1.782288e-11, 1.793743e-11, 1.759681e-11, 
    1.739352e-11, 1.725914e-11, 1.716408e-11, 1.71775e-11, 1.72031e-11, 
    1.733497e-11, 1.745939e-11, 1.75545e-11, 1.761826e-11, 1.76812e-11, 
    1.787234e-11, 1.797393e-11, 1.820239e-11, 1.816106e-11, 1.82311e-11, 
    1.829815e-11, 1.841096e-11, 1.839237e-11, 1.844216e-11, 1.822926e-11, 
    1.837062e-11, 1.813754e-11, 1.820115e-11, 1.76983e-11, 1.750856e-11, 
    1.742819e-11, 1.735801e-11, 1.718783e-11, 1.730526e-11, 1.725892e-11, 
    1.736928e-11, 1.743957e-11, 1.740479e-11, 1.762001e-11, 1.753618e-11, 
    1.797996e-11, 1.778815e-11, 1.829032e-11, 1.816954e-11, 1.831933e-11, 
    1.824282e-11, 1.8374e-11, 1.825592e-11, 1.846071e-11, 1.850544e-11, 
    1.847487e-11, 1.859246e-11, 1.824938e-11, 1.838077e-11, 1.740381e-11, 
    1.740948e-11, 1.743592e-11, 1.731987e-11, 1.731279e-11, 1.720681e-11, 
    1.73011e-11, 1.734132e-11, 1.744365e-11, 1.750432e-11, 1.756208e-11, 
    1.76894e-11, 1.783212e-11, 1.803263e-11, 1.817736e-11, 1.827468e-11, 
    1.821497e-11, 1.826768e-11, 1.820877e-11, 1.818118e-11, 1.848867e-11, 
    1.831571e-11, 1.857553e-11, 1.85611e-11, 1.844334e-11, 1.856273e-11, 
    1.741347e-11, 1.738085e-11, 1.726781e-11, 1.735624e-11, 1.719528e-11, 
    1.728529e-11, 1.733714e-11, 1.753793e-11, 1.75822e-11, 1.762329e-11, 
    1.770459e-11, 1.780919e-11, 1.799341e-11, 1.815444e-11, 1.830205e-11, 
    1.829122e-11, 1.829503e-11, 1.832808e-11, 1.824627e-11, 1.834152e-11, 
    1.835753e-11, 1.831569e-11, 1.855917e-11, 1.848945e-11, 1.85608e-11, 
    1.851539e-11, 1.739145e-11, 1.744637e-11, 1.741668e-11, 1.747253e-11, 
    1.743317e-11, 1.760851e-11, 1.766124e-11, 1.790901e-11, 1.780713e-11, 
    1.796942e-11, 1.782359e-11, 1.784938e-11, 1.797472e-11, 1.783145e-11, 
    1.814554e-11, 1.79323e-11, 1.832936e-11, 1.811537e-11, 1.834281e-11, 
    1.830141e-11, 1.836998e-11, 1.84315e-11, 1.850903e-11, 1.86525e-11, 
    1.861923e-11, 1.873953e-11, 1.752841e-11, 1.759994e-11, 1.759364e-11, 
    1.766864e-11, 1.77242e-11, 1.784492e-11, 1.803937e-11, 1.796613e-11, 
    1.81007e-11, 1.812777e-11, 1.792337e-11, 1.804873e-11, 1.764789e-11, 
    1.771236e-11, 1.767396e-11, 1.753405e-11, 1.798299e-11, 1.77519e-11, 
    1.817975e-11, 1.805373e-11, 1.842272e-11, 1.823876e-11, 1.860093e-11, 
    1.875679e-11, 1.890408e-11, 1.907688e-11, 1.763904e-11, 1.759037e-11, 
    1.767757e-11, 1.779854e-11, 1.791116e-11, 1.80614e-11, 1.807681e-11, 
    1.810503e-11, 1.817824e-11, 1.823991e-11, 1.811396e-11, 1.825538e-11, 
    1.772731e-11, 1.800312e-11, 1.757199e-11, 1.770127e-11, 1.77914e-11, 
    1.775184e-11, 1.795777e-11, 1.800647e-11, 1.820503e-11, 1.810226e-11, 
    1.871826e-11, 1.84445e-11, 1.920897e-11, 1.899382e-11, 1.757338e-11, 
    1.763888e-11, 1.786773e-11, 1.775867e-11, 1.807145e-11, 1.814885e-11, 
    1.821189e-11, 1.829261e-11, 1.830134e-11, 1.834927e-11, 1.827077e-11, 
    1.834616e-11, 1.806172e-11, 1.818857e-11, 1.784151e-11, 1.792568e-11, 
    1.788693e-11, 1.784448e-11, 1.797567e-11, 1.811593e-11, 1.811894e-11, 
    1.816404e-11, 1.829138e-11, 1.807273e-11, 1.875373e-11, 1.833171e-11, 
    1.771043e-11, 1.783715e-11, 1.78553e-11, 1.780613e-11, 1.814108e-11, 
    1.801937e-11, 1.83481e-11, 1.825897e-11, 1.840512e-11, 1.833242e-11, 
    1.832174e-11, 1.822861e-11, 1.817074e-11, 1.802494e-11, 1.790673e-11, 
    1.781326e-11, 1.783497e-11, 1.793772e-11, 1.812453e-11, 1.830213e-11, 
    1.826315e-11, 1.839399e-11, 1.804868e-11, 1.819309e-11, 1.813721e-11, 
    1.828309e-11, 1.796419e-11, 1.823556e-11, 1.789513e-11, 1.792486e-11, 
    1.801695e-11, 1.82029e-11, 1.824417e-11, 1.828828e-11, 1.826106e-11, 
    1.812929e-11, 1.810775e-11, 1.801471e-11, 1.798907e-11, 1.791838e-11, 
    1.785997e-11, 1.791333e-11, 1.796946e-11, 1.812935e-11, 1.827401e-11, 
    1.843237e-11, 1.847123e-11, 1.865726e-11, 1.850575e-11, 1.875609e-11, 
    1.854314e-11, 1.891252e-11, 1.825136e-11, 1.85369e-11, 1.802115e-11, 
    1.807638e-11, 1.817647e-11, 1.840706e-11, 1.82824e-11, 1.842823e-11, 
    1.81069e-11, 1.794126e-11, 1.789854e-11, 1.781893e-11, 1.790036e-11, 
    1.789373e-11, 1.79718e-11, 1.794669e-11, 1.813467e-11, 1.803358e-11, 
    1.832147e-11, 1.842708e-11, 1.87269e-11, 1.891185e-11, 1.910102e-11, 
    1.918483e-11, 1.921037e-11, 1.922105e-11,
  1.87948e-11, 1.897033e-11, 1.893613e-11, 1.907825e-11, 1.899934e-11, 
    1.90925e-11, 1.883031e-11, 1.897732e-11, 1.888339e-11, 1.881056e-11, 
    1.93558e-11, 1.90846e-11, 1.963983e-11, 1.946515e-11, 1.990568e-11, 
    1.961259e-11, 1.996508e-11, 1.989718e-11, 2.010193e-11, 2.004315e-11, 
    2.030639e-11, 2.01291e-11, 2.044363e-11, 2.026396e-11, 2.029201e-11, 
    2.012327e-11, 1.9139e-11, 1.932192e-11, 1.912819e-11, 1.91542e-11, 
    1.914253e-11, 1.900096e-11, 1.892986e-11, 1.878142e-11, 1.880832e-11, 
    1.891736e-11, 1.916591e-11, 1.908133e-11, 1.92949e-11, 1.929006e-11, 
    1.952942e-11, 1.942129e-11, 1.982615e-11, 1.971059e-11, 2.00456e-11, 
    1.996104e-11, 2.004163e-11, 2.001717e-11, 2.004195e-11, 1.991801e-11, 
    1.997106e-11, 1.98622e-11, 1.944151e-11, 1.956461e-11, 1.919881e-11, 
    1.898078e-11, 1.883674e-11, 1.873492e-11, 1.87493e-11, 1.877672e-11, 
    1.8918e-11, 1.905139e-11, 1.91534e-11, 1.922182e-11, 1.928937e-11, 
    1.949468e-11, 1.960384e-11, 1.984957e-11, 1.980509e-11, 1.988047e-11, 
    1.995264e-11, 2.007415e-11, 2.005412e-11, 2.010776e-11, 1.987848e-11, 
    2.003069e-11, 1.977978e-11, 1.984822e-11, 1.930777e-11, 1.910412e-11, 
    1.901796e-11, 1.89427e-11, 1.876035e-11, 1.888617e-11, 1.883652e-11, 
    1.895477e-11, 1.903014e-11, 1.899284e-11, 1.922369e-11, 1.913375e-11, 
    1.961033e-11, 1.940422e-11, 1.994421e-11, 1.981421e-11, 1.997545e-11, 
    1.989308e-11, 2.003434e-11, 1.990718e-11, 2.012775e-11, 2.017597e-11, 
    2.014301e-11, 2.026978e-11, 1.990014e-11, 2.004163e-11, 1.89918e-11, 
    1.899787e-11, 1.902621e-11, 1.890183e-11, 1.889424e-11, 1.878068e-11, 
    1.88817e-11, 1.892481e-11, 1.903451e-11, 1.909957e-11, 1.916153e-11, 
    1.929817e-11, 1.945145e-11, 1.966695e-11, 1.982262e-11, 1.992737e-11, 
    1.98631e-11, 1.991984e-11, 1.985642e-11, 1.982674e-11, 2.015789e-11, 
    1.997155e-11, 2.025151e-11, 2.023596e-11, 2.010904e-11, 2.023771e-11, 
    1.900215e-11, 1.896717e-11, 1.884603e-11, 1.894079e-11, 1.876834e-11, 
    1.886476e-11, 1.892034e-11, 1.913563e-11, 1.918312e-11, 1.922722e-11, 
    1.931448e-11, 1.942681e-11, 1.962478e-11, 1.979797e-11, 1.995684e-11, 
    1.994518e-11, 1.994928e-11, 1.998487e-11, 1.989679e-11, 1.999935e-11, 
    2.00166e-11, 1.997153e-11, 2.023388e-11, 2.015873e-11, 2.023563e-11, 
    2.018668e-11, 1.897853e-11, 1.903743e-11, 1.900559e-11, 1.906548e-11, 
    1.902328e-11, 1.921136e-11, 1.926796e-11, 1.953407e-11, 1.94246e-11, 
    1.959899e-11, 1.944227e-11, 1.946999e-11, 1.96047e-11, 1.945072e-11, 
    1.97884e-11, 1.95591e-11, 1.998625e-11, 1.975595e-11, 2.000074e-11, 
    1.995615e-11, 2.003e-11, 2.009628e-11, 2.017983e-11, 2.033454e-11, 
    2.029865e-11, 2.042843e-11, 1.912541e-11, 1.920216e-11, 1.91954e-11, 
    1.927588e-11, 1.933554e-11, 1.946519e-11, 1.967419e-11, 1.959545e-11, 
    1.974015e-11, 1.976927e-11, 1.954949e-11, 1.968427e-11, 1.925362e-11, 
    1.932283e-11, 1.928161e-11, 1.913147e-11, 1.961358e-11, 1.936529e-11, 
    1.98252e-11, 1.968963e-11, 2.008682e-11, 1.988872e-11, 2.027891e-11, 
    2.044708e-11, 2.060608e-11, 2.079283e-11, 1.924412e-11, 1.919189e-11, 
    1.928547e-11, 1.941538e-11, 1.953636e-11, 1.969788e-11, 1.971445e-11, 
    1.974481e-11, 1.982358e-11, 1.988994e-11, 1.975442e-11, 1.99066e-11, 
    1.933891e-11, 1.963522e-11, 1.917217e-11, 1.931093e-11, 1.940771e-11, 
    1.936522e-11, 1.958646e-11, 1.963881e-11, 1.985241e-11, 1.974182e-11, 
    2.04055e-11, 2.01103e-11, 2.093567e-11, 2.070306e-11, 1.917366e-11, 
    1.924394e-11, 1.948971e-11, 1.937255e-11, 1.970869e-11, 1.979195e-11, 
    1.985978e-11, 1.994669e-11, 1.995608e-11, 2.000769e-11, 1.992316e-11, 
    2.000435e-11, 1.969823e-11, 1.983469e-11, 1.946152e-11, 1.955197e-11, 
    1.951033e-11, 1.946471e-11, 1.96057e-11, 1.975655e-11, 1.975978e-11, 
    1.980829e-11, 1.99454e-11, 1.971006e-11, 2.04438e-11, 1.998883e-11, 
    1.932075e-11, 1.945686e-11, 1.947634e-11, 1.942352e-11, 1.978359e-11, 
    1.965268e-11, 2.000643e-11, 1.991046e-11, 2.006785e-11, 1.998955e-11, 
    1.997805e-11, 1.987778e-11, 1.981551e-11, 1.965868e-11, 1.95316e-11, 
    1.943117e-11, 1.94545e-11, 1.956491e-11, 1.97658e-11, 1.995694e-11, 
    1.991498e-11, 2.005586e-11, 1.968421e-11, 1.983956e-11, 1.977943e-11, 
    1.993643e-11, 1.959336e-11, 1.98853e-11, 1.951914e-11, 1.955108e-11, 
    1.965009e-11, 1.985013e-11, 1.989453e-11, 1.994202e-11, 1.991271e-11, 
    1.977091e-11, 1.974773e-11, 1.964768e-11, 1.962011e-11, 1.954412e-11, 
    1.948135e-11, 1.95387e-11, 1.959904e-11, 1.977097e-11, 1.992666e-11, 
    2.009722e-11, 2.013909e-11, 2.03397e-11, 2.017631e-11, 2.044635e-11, 
    2.021665e-11, 2.061524e-11, 1.990229e-11, 2.02099e-11, 1.96546e-11, 
    1.971399e-11, 1.982168e-11, 2.006995e-11, 1.993569e-11, 2.009276e-11, 
    1.974683e-11, 1.956873e-11, 1.952279e-11, 1.943727e-11, 1.952475e-11, 
    1.951763e-11, 1.960153e-11, 1.957455e-11, 1.977669e-11, 1.966796e-11, 
    1.997776e-11, 2.009152e-11, 2.041481e-11, 2.061449e-11, 2.081892e-11, 
    2.090955e-11, 2.093718e-11, 2.094874e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
