netcdf ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-12-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-12-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to patch-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to patch-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "timestep fractional area burned" ;
		FAREA_BURNED:units = "proportion" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "patch-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total patch-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float RSCANOPY(time, lndgrid) ;
		RSCANOPY:long_name = "canopy resistance" ;
		RSCANOPY:units = " s m-1" ;
		RSCANOPY:cell_methods = "time: mean" ;
		RSCANOPY:_FillValue = 1.e+36f ;
		RSCANOPY:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new Patches" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total patch-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C eallocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 10/28/14 13:17:34" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-12-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 11202 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "10/28/14" ;

 time_written =
  "13:17:34" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  5.065059e-14, 5.07875e-14, 5.076091e-14, 5.087123e-14, 5.081006e-14, 
    5.088227e-14, 5.067837e-14, 5.079292e-14, 5.071982e-14, 5.066294e-14, 
    5.1085e-14, 5.087615e-14, 5.130174e-14, 5.116879e-14, 5.150255e-14, 
    5.128103e-14, 5.154717e-14, 5.149621e-14, 5.164964e-14, 5.160571e-14, 
    5.180164e-14, 5.166991e-14, 5.190315e-14, 5.177022e-14, 5.179101e-14, 
    5.166555e-14, 5.091825e-14, 5.1059e-14, 5.09099e-14, 5.092998e-14, 
    5.092098e-14, 5.081131e-14, 5.075598e-14, 5.064015e-14, 5.066119e-14, 
    5.074628e-14, 5.093901e-14, 5.087365e-14, 5.10384e-14, 5.103468e-14, 
    5.121782e-14, 5.113528e-14, 5.144272e-14, 5.135543e-14, 5.160754e-14, 
    5.154418e-14, 5.160456e-14, 5.158626e-14, 5.16048e-14, 5.151186e-14, 
    5.155169e-14, 5.146989e-14, 5.115073e-14, 5.124461e-14, 5.096441e-14, 
    5.079556e-14, 5.06834e-14, 5.060371e-14, 5.061498e-14, 5.063645e-14, 
    5.074677e-14, 5.085045e-14, 5.092939e-14, 5.098216e-14, 5.103415e-14, 
    5.119125e-14, 5.127441e-14, 5.146034e-14, 5.142685e-14, 5.148361e-14, 
    5.153788e-14, 5.162887e-14, 5.161391e-14, 5.165397e-14, 5.148214e-14, 
    5.159635e-14, 5.140775e-14, 5.145936e-14, 5.104813e-14, 5.089129e-14, 
    5.082445e-14, 5.076601e-14, 5.062364e-14, 5.072197e-14, 5.068321e-14, 
    5.077543e-14, 5.083397e-14, 5.080502e-14, 5.098361e-14, 5.091421e-14, 
    5.127934e-14, 5.11222e-14, 5.153155e-14, 5.143372e-14, 5.155499e-14, 
    5.149313e-14, 5.159909e-14, 5.150374e-14, 5.166889e-14, 5.170481e-14, 
    5.168026e-14, 5.177457e-14, 5.149844e-14, 5.160454e-14, 5.080421e-14, 
    5.080893e-14, 5.083093e-14, 5.073417e-14, 5.072826e-14, 5.063956e-14, 
    5.07185e-14, 5.075209e-14, 5.083737e-14, 5.088776e-14, 5.093566e-14, 
    5.10409e-14, 5.115831e-14, 5.132234e-14, 5.144007e-14, 5.151892e-14, 
    5.147058e-14, 5.151325e-14, 5.146554e-14, 5.144318e-14, 5.169134e-14, 
    5.155205e-14, 5.176101e-14, 5.174946e-14, 5.165492e-14, 5.175076e-14, 
    5.081224e-14, 5.078507e-14, 5.069065e-14, 5.076455e-14, 5.06299e-14, 
    5.070527e-14, 5.074858e-14, 5.091562e-14, 5.095233e-14, 5.098631e-14, 
    5.105343e-14, 5.113951e-14, 5.129034e-14, 5.142145e-14, 5.154104e-14, 
    5.153229e-14, 5.153537e-14, 5.156205e-14, 5.149592e-14, 5.157291e-14, 
    5.158581e-14, 5.155205e-14, 5.174791e-14, 5.169199e-14, 5.174921e-14, 
    5.171281e-14, 5.079391e-14, 5.083963e-14, 5.081492e-14, 5.086136e-14, 
    5.082864e-14, 5.097406e-14, 5.101763e-14, 5.122133e-14, 5.11378e-14, 
    5.127075e-14, 5.115133e-14, 5.117249e-14, 5.127502e-14, 5.115779e-14, 
    5.14142e-14, 5.124037e-14, 5.156309e-14, 5.138965e-14, 5.157395e-14, 
    5.154053e-14, 5.159587e-14, 5.16454e-14, 5.170771e-14, 5.182254e-14, 
    5.179597e-14, 5.189196e-14, 5.090776e-14, 5.096699e-14, 5.09618e-14, 
    5.102377e-14, 5.106958e-14, 5.116884e-14, 5.132784e-14, 5.126809e-14, 
    5.13778e-14, 5.13998e-14, 5.123313e-14, 5.133547e-14, 5.100663e-14, 
    5.105979e-14, 5.102816e-14, 5.091242e-14, 5.128182e-14, 5.109236e-14, 
    5.1442e-14, 5.133955e-14, 5.163833e-14, 5.14898e-14, 5.178133e-14, 
    5.190566e-14, 5.202267e-14, 5.215911e-14, 5.099933e-14, 5.09591e-14, 
    5.103115e-14, 5.113072e-14, 5.122311e-14, 5.13458e-14, 5.135836e-14, 
    5.138131e-14, 5.14408e-14, 5.149077e-14, 5.138855e-14, 5.15033e-14, 
    5.107206e-14, 5.129826e-14, 5.094386e-14, 5.105065e-14, 5.112487e-14, 
    5.109234e-14, 5.126126e-14, 5.130103e-14, 5.146249e-14, 5.137907e-14, 
    5.187496e-14, 5.165582e-14, 5.226298e-14, 5.209362e-14, 5.094503e-14, 
    5.09992e-14, 5.118753e-14, 5.109796e-14, 5.135399e-14, 5.141692e-14, 
    5.146808e-14, 5.15334e-14, 5.154046e-14, 5.157915e-14, 5.151575e-14, 
    5.157666e-14, 5.134606e-14, 5.144916e-14, 5.116605e-14, 5.1235e-14, 
    5.120329e-14, 5.116848e-14, 5.127588e-14, 5.139015e-14, 5.139263e-14, 
    5.142924e-14, 5.153227e-14, 5.135503e-14, 5.190313e-14, 5.156487e-14, 
    5.105825e-14, 5.116242e-14, 5.117735e-14, 5.1137e-14, 5.141061e-14, 
    5.131154e-14, 5.157821e-14, 5.150621e-14, 5.162417e-14, 5.156557e-14, 
    5.155694e-14, 5.148162e-14, 5.14347e-14, 5.131607e-14, 5.121948e-14, 
    5.114286e-14, 5.116068e-14, 5.124484e-14, 5.139715e-14, 5.154109e-14, 
    5.150956e-14, 5.161521e-14, 5.133544e-14, 5.145281e-14, 5.140745e-14, 
    5.152571e-14, 5.126649e-14, 5.148713e-14, 5.121001e-14, 5.123434e-14, 
    5.130957e-14, 5.146074e-14, 5.149423e-14, 5.152989e-14, 5.150789e-14, 
    5.140102e-14, 5.138352e-14, 5.130775e-14, 5.12868e-14, 5.122905e-14, 
    5.118119e-14, 5.12249e-14, 5.127079e-14, 5.140108e-14, 5.151836e-14, 
    5.16461e-14, 5.167735e-14, 5.182628e-14, 5.170501e-14, 5.1905e-14, 
    5.17349e-14, 5.202925e-14, 5.149997e-14, 5.172998e-14, 5.131301e-14, 
    5.135801e-14, 5.143931e-14, 5.162568e-14, 5.152515e-14, 5.164273e-14, 
    5.138283e-14, 5.124772e-14, 5.121279e-14, 5.114751e-14, 5.121429e-14, 
    5.120886e-14, 5.127272e-14, 5.125221e-14, 5.14054e-14, 5.132314e-14, 
    5.155671e-14, 5.164182e-14, 5.188189e-14, 5.202878e-14, 5.217819e-14, 
    5.224405e-14, 5.22641e-14, 5.227248e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -7.470118e-15, -7.463324e-15, -7.464646e-15, -7.459169e-15, -7.462208e-15, 
    -7.458621e-15, -7.468743e-15, -7.463052e-15, -7.466686e-15, -7.46951e-15, 
    -7.448549e-15, -7.458925e-15, -7.437819e-15, -7.444415e-15, 
    -7.427872e-15, -7.438842e-15, -7.425665e-15, -7.428194e-15, 
    -7.420599e-15, -7.422774e-15, -7.39021e-15, -7.419595e-15, -7.385129e-15, 
    -7.391795e-15, -7.390747e-15, -7.41981e-15, -7.45684e-15, -7.449839e-15, 
    -7.457254e-15, -7.456255e-15, -7.456705e-15, -7.462143e-15, 
    -7.464883e-15, -7.470642e-15, -7.469596e-15, -7.465369e-15, 
    -7.455806e-15, -7.459054e-15, -7.450884e-15, -7.451068e-15, 
    -7.441986e-15, -7.446079e-15, -7.430842e-15, -7.435169e-15, 
    -7.422684e-15, -7.425819e-15, -7.422829e-15, -7.423736e-15, 
    -7.422817e-15, -7.427418e-15, -7.425447e-15, -7.429498e-15, -7.44531e-15, 
    -7.440656e-15, -7.454549e-15, -7.462914e-15, -7.468492e-15, -7.47245e-15, 
    -7.47189e-15, -7.470822e-15, -7.465344e-15, -7.460205e-15, -7.45629e-15, 
    -7.453672e-15, -7.451095e-15, -7.443288e-15, -7.439174e-15, 
    -7.429965e-15, -7.43163e-15, -7.428814e-15, -7.426132e-15, -7.421625e-15, 
    -7.422367e-15, -7.420381e-15, -7.428891e-15, -7.423232e-15, 
    -7.432578e-15, -7.430019e-15, -7.450376e-15, -7.458178e-15, 
    -7.461483e-15, -7.464391e-15, -7.471459e-15, -7.466576e-15, -7.4685e-15, 
    -7.463928e-15, -7.461022e-15, -7.462459e-15, -7.4536e-15, -7.457042e-15, 
    -7.43893e-15, -7.446723e-15, -7.426444e-15, -7.431289e-15, -7.425285e-15, 
    -7.428348e-15, -7.423099e-15, -7.427823e-15, -7.419644e-15, 
    -7.395107e-15, -7.419079e-15, -7.391579e-15, -7.428085e-15, 
    -7.422828e-15, -7.462499e-15, -7.462265e-15, -7.461174e-15, 
    -7.465969e-15, -7.466264e-15, -7.47067e-15, -7.466751e-15, -7.465083e-15, 
    -7.460855e-15, -7.458353e-15, -7.455977e-15, -7.450758e-15, 
    -7.444932e-15, -7.436803e-15, -7.430974e-15, -7.427072e-15, 
    -7.429466e-15, -7.427352e-15, -7.429714e-15, -7.430823e-15, 
    -7.395799e-15, -7.425427e-15, -7.392262e-15, -7.392844e-15, 
    -7.420333e-15, -7.392779e-15, -7.4621e-15, -7.46345e-15, -7.468133e-15, 
    -7.464468e-15, -7.47115e-15, -7.467406e-15, -7.465253e-15, -7.456966e-15, 
    -7.455152e-15, -7.453464e-15, -7.450138e-15, -7.445869e-15, 
    -7.438389e-15, -7.431894e-15, -7.425977e-15, -7.42641e-15, -7.426257e-15, 
    -7.424934e-15, -7.42821e-15, -7.424397e-15, -7.423756e-15, -7.42543e-15, 
    -7.392923e-15, -7.395766e-15, -7.392857e-15, -7.394701e-15, 
    -7.463012e-15, -7.460742e-15, -7.461968e-15, -7.459662e-15, 
    -7.461285e-15, -7.454066e-15, -7.451904e-15, -7.441805e-15, 
    -7.445952e-15, -7.439359e-15, -7.445283e-15, -7.444232e-15, 
    -7.439136e-15, -7.444964e-15, -7.432248e-15, -7.440858e-15, 
    -7.424883e-15, -7.433459e-15, -7.424345e-15, -7.426002e-15, 
    -7.423261e-15, -7.420807e-15, -7.39496e-15, -7.389166e-15, -7.390501e-15, 
    -7.385691e-15, -7.457362e-15, -7.45442e-15, -7.454683e-15, -7.451608e-15, 
    -7.449335e-15, -7.444416e-15, -7.436533e-15, -7.439497e-15, 
    -7.434061e-15, -7.432969e-15, -7.44123e-15, -7.436153e-15, -7.452455e-15, 
    -7.449813e-15, -7.451389e-15, -7.457127e-15, -7.438809e-15, 
    -7.448199e-15, -7.430878e-15, -7.435954e-15, -7.421156e-15, 
    -7.428505e-15, -7.391237e-15, -7.384998e-15, -7.379166e-15, 
    -7.372362e-15, -7.452819e-15, -7.454817e-15, -7.451244e-15, 
    -7.446298e-15, -7.441723e-15, -7.435644e-15, -7.435024e-15, 
    -7.433885e-15, -7.43094e-15, -7.428465e-15, -7.433521e-15, -7.427845e-15, 
    -7.449194e-15, -7.437996e-15, -7.455569e-15, -7.450265e-15, -7.44659e-15, 
    -7.448206e-15, -7.439837e-15, -7.437865e-15, -7.42986e-15, -7.433998e-15, 
    -7.386532e-15, -7.420283e-15, -7.367204e-15, -7.375624e-15, 
    -7.455514e-15, -7.452828e-15, -7.443484e-15, -7.447928e-15, -7.43524e-15, 
    -7.43212e-15, -7.429589e-15, -7.426351e-15, -7.426004e-15, -7.424086e-15, 
    -7.427229e-15, -7.424212e-15, -7.43563e-15, -7.430525e-15, -7.444556e-15, 
    -7.441134e-15, -7.442709e-15, -7.444435e-15, -7.439111e-15, 
    -7.433441e-15, -7.433326e-15, -7.431508e-15, -7.426381e-15, 
    -7.435189e-15, -7.385112e-15, -7.424771e-15, -7.4499e-15, -7.444724e-15, 
    -7.443992e-15, -7.445995e-15, -7.432433e-15, -7.437341e-15, 
    -7.424135e-15, -7.427701e-15, -7.421859e-15, -7.424761e-15, 
    -7.425187e-15, -7.428918e-15, -7.43124e-15, -7.437115e-15, -7.441903e-15, 
    -7.445705e-15, -7.444822e-15, -7.440646e-15, -7.433095e-15, -7.42597e-15, 
    -7.427529e-15, -7.422303e-15, -7.436159e-15, -7.43034e-15, -7.432586e-15, 
    -7.426734e-15, -7.439574e-15, -7.42862e-15, -7.442376e-15, -7.44117e-15, 
    -7.43744e-15, -7.429942e-15, -7.428294e-15, -7.426525e-15, -7.427618e-15, 
    -7.432906e-15, -7.433775e-15, -7.437531e-15, -7.438566e-15, 
    -7.441433e-15, -7.443805e-15, -7.441636e-15, -7.439358e-15, 
    -7.432906e-15, -7.427096e-15, -7.420771e-15, -7.419226e-15, 
    -7.388969e-15, -7.395092e-15, -7.385018e-15, -7.393563e-15, 
    -7.378822e-15, -7.427995e-15, -7.39382e-15, -7.437271e-15, -7.435042e-15, 
    -7.431005e-15, -7.421774e-15, -7.426762e-15, -7.420932e-15, 
    -7.433809e-15, -7.440498e-15, -7.442238e-15, -7.445473e-15, 
    -7.442164e-15, -7.442433e-15, -7.439268e-15, -7.440286e-15, 
    -7.432691e-15, -7.436769e-15, -7.425197e-15, -7.420979e-15, 
    -7.386193e-15, -7.378855e-15, -7.371422e-15, -7.368146e-15, 
    -7.367151e-15, -7.366734e-15 ;

 CH4_SURF_DIFF_UNSAT =
  4.838033e-14, 4.786322e-14, 4.796389e-14, 4.754587e-14, 4.777791e-14, 
    4.750399e-14, 4.827565e-14, 4.784262e-14, 4.811921e-14, 4.833389e-14, 
    4.673166e-14, 4.752721e-14, 4.590192e-14, 4.641199e-14, 4.512808e-14, 
    4.598133e-14, 4.495558e-14, 4.515284e-14, 4.455873e-14, 4.472913e-14, 
    4.383215e-14, 4.448003e-14, 4.343679e-14, 4.395464e-14, 4.387367e-14, 
    4.449692e-14, 4.736749e-14, 4.683087e-14, 4.73992e-14, 4.73228e-14, 
    4.735711e-14, 4.777309e-14, 4.798228e-14, 4.841985e-14, 4.834051e-14, 
    4.801912e-14, 4.728844e-14, 4.753688e-14, 4.691026e-14, 4.692444e-14, 
    4.622421e-14, 4.654027e-14, 4.535936e-14, 4.569579e-14, 4.472202e-14, 
    4.496737e-14, 4.473353e-14, 4.480448e-14, 4.473261e-14, 4.509232e-14, 
    4.493828e-14, 4.525454e-14, 4.64811e-14, 4.612145e-14, 4.719193e-14, 
    4.783236e-14, 4.825667e-14, 4.855705e-14, 4.851462e-14, 4.843368e-14, 
    4.801724e-14, 4.762486e-14, 4.732521e-14, 4.712448e-14, 4.692648e-14, 
    4.632555e-14, 4.600689e-14, 4.529121e-14, 4.542065e-14, 4.520138e-14, 
    4.499176e-14, 4.463922e-14, 4.469731e-14, 4.454181e-14, 4.520723e-14, 
    4.476521e-14, 4.549433e-14, 4.529518e-14, 4.687229e-14, 4.74699e-14, 
    4.772303e-14, 4.794453e-14, 4.848198e-14, 4.811099e-14, 4.825732e-14, 
    4.790905e-14, 4.768733e-14, 4.779704e-14, 4.711899e-14, 4.738289e-14, 
    4.598799e-14, 4.659016e-14, 4.501622e-14, 4.53941e-14, 4.492555e-14, 
    4.516481e-14, 4.475465e-14, 4.512382e-14, 4.448393e-14, 4.420894e-14, 
    4.443971e-14, 4.39379e-14, 4.514426e-14, 4.47335e-14, 4.78001e-14, 
    4.778221e-14, 4.769888e-14, 4.806486e-14, 4.808724e-14, 4.842201e-14, 
    4.81242e-14, 4.799719e-14, 4.76745e-14, 4.748328e-14, 4.730134e-14, 
    4.690064e-14, 4.645201e-14, 4.582289e-14, 4.536963e-14, 4.506515e-14, 
    4.525194e-14, 4.508704e-14, 4.527135e-14, 4.535769e-14, 4.426127e-14, 
    4.493683e-14, 4.399062e-14, 4.403554e-14, 4.453809e-14, 4.403048e-14, 
    4.776965e-14, 4.787256e-14, 4.82293e-14, 4.795019e-14, 4.845843e-14, 
    4.817408e-14, 4.801035e-14, 4.737731e-14, 4.7238e-14, 4.710861e-14, 
    4.685288e-14, 4.65241e-14, 4.594588e-14, 4.544133e-14, 4.497958e-14, 
    4.501345e-14, 4.500153e-14, 4.48982e-14, 4.515399e-14, 4.485617e-14, 
    4.480611e-14, 4.493693e-14, 4.404155e-14, 4.425888e-14, 4.403649e-14, 
    4.417799e-14, 4.783913e-14, 4.76659e-14, 4.775952e-14, 4.758342e-14, 
    4.770748e-14, 4.715506e-14, 4.69891e-14, 4.621055e-14, 4.653056e-14, 
    4.602109e-14, 4.64789e-14, 4.639785e-14, 4.600431e-14, 4.645421e-14, 
    4.546912e-14, 4.613744e-14, 4.489418e-14, 4.556351e-14, 4.485215e-14, 
    4.498158e-14, 4.476727e-14, 4.45751e-14, 4.419779e-14, 4.375104e-14, 
    4.385455e-14, 4.348058e-14, 4.740737e-14, 4.718208e-14, 4.720198e-14, 
    4.696597e-14, 4.67912e-14, 4.641191e-14, 4.580182e-14, 4.60315e-14, 
    4.560969e-14, 4.552488e-14, 4.616565e-14, 4.577243e-14, 4.703118e-14, 
    4.682834e-14, 4.694918e-14, 4.738958e-14, 4.597851e-14, 4.670403e-14, 
    4.536211e-14, 4.575684e-14, 4.460251e-14, 4.517741e-14, 4.391151e-14, 
    4.342679e-14, 4.29699e-14, 4.243443e-14, 4.705906e-14, 4.721228e-14, 
    4.69379e-14, 4.655747e-14, 4.620394e-14, 4.573278e-14, 4.568454e-14, 
    4.55961e-14, 4.536688e-14, 4.517391e-14, 4.556806e-14, 4.512551e-14, 
    4.678115e-14, 4.591543e-14, 4.727011e-14, 4.686318e-14, 4.657994e-14, 
    4.670431e-14, 4.605775e-14, 4.5905e-14, 4.528297e-14, 4.560482e-14, 
    4.354647e-14, 4.45344e-14, 4.202601e-14, 4.269163e-14, 4.726576e-14, 
    4.705962e-14, 4.63402e-14, 4.668287e-14, 4.570132e-14, 4.545887e-14, 
    4.52616e-14, 4.500902e-14, 4.498178e-14, 4.483196e-14, 4.50774e-14, 
    4.484168e-14, 4.573177e-14, 4.533455e-14, 4.642265e-14, 4.615837e-14, 
    4.628002e-14, 4.641331e-14, 4.60016e-14, 4.556185e-14, 4.555254e-14, 
    4.541129e-14, 4.501248e-14, 4.569733e-14, 4.343609e-14, 4.488646e-14, 
    4.683455e-14, 4.643616e-14, 4.63793e-14, 4.653376e-14, 4.548319e-14, 
    4.586453e-14, 4.483562e-14, 4.511428e-14, 4.465752e-14, 4.488462e-14, 
    4.4918e-14, 4.520926e-14, 4.539034e-14, 4.584705e-14, 4.621784e-14, 
    4.651138e-14, 4.644317e-14, 4.612058e-14, 4.553494e-14, 4.497927e-14, 
    4.510111e-14, 4.469227e-14, 4.577266e-14, 4.532034e-14, 4.549526e-14, 
    4.503883e-14, 4.603758e-14, 4.518713e-14, 4.625429e-14, 4.616099e-14, 
    4.58721e-14, 4.528956e-14, 4.516057e-14, 4.502258e-14, 4.510776e-14, 
    4.552006e-14, 4.558757e-14, 4.587915e-14, 4.595952e-14, 4.618132e-14, 
    4.636469e-14, 4.619713e-14, 4.602098e-14, 4.551993e-14, 4.506717e-14, 
    4.457235e-14, 4.44511e-14, 4.373605e-14, 4.420788e-14, 4.342873e-14, 
    4.409109e-14, 4.294341e-14, 4.513787e-14, 4.411071e-14, 4.585897e-14, 
    4.568589e-14, 4.53723e-14, 4.465129e-14, 4.504098e-14, 4.458522e-14, 
    4.559022e-14, 4.610939e-14, 4.62436e-14, 4.649353e-14, 4.623788e-14, 
    4.625869e-14, 4.601375e-14, 4.60925e-14, 4.550327e-14, 4.582002e-14, 
    4.491881e-14, 4.458884e-14, 4.351977e-14, 4.294568e-14, 4.235986e-14, 
    4.210068e-14, 4.202173e-14, 4.198872e-14 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931953e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 1.931952e-23, 
    1.931951e-23, 1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 
    1.93195e-23, 1.931951e-23, 1.931948e-23, 1.931949e-23, 1.931947e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931945e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931945e-23, 
    1.931946e-23, 1.931951e-23, 1.93195e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 
    1.931952e-23, 1.931951e-23, 1.931951e-23, 1.93195e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.931947e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931949e-23, 1.931949e-23, 1.931951e-23, 
    1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931952e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 1.93195e-23, 
    1.931949e-23, 1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 1.931947e-23, 
    1.931946e-23, 1.931948e-23, 1.931947e-23, 1.93195e-23, 1.931951e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 
    1.931949e-23, 1.93195e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 1.931945e-23, 
    1.931946e-23, 1.931945e-23, 1.931947e-23, 1.931946e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 
    1.931947e-23, 1.931945e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931953e-23, 
    1.931953e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 
    1.931946e-23, 1.931947e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931945e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931951e-23, 1.93195e-23, 1.931949e-23, 1.93195e-23, 
    1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931949e-23, 
    1.931947e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931945e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931948e-23, 1.93195e-23, 
    1.93195e-23, 1.93195e-23, 1.931951e-23, 1.931948e-23, 1.93195e-23, 
    1.931947e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 
    1.931944e-23, 1.931943e-23, 1.931942e-23, 1.93195e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.93195e-23, 1.931948e-23, 1.931951e-23, 1.93195e-23, 1.93195e-23, 
    1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931944e-23, 1.931946e-23, 1.931941e-23, 1.931943e-23, 1.931951e-23, 
    1.93195e-23, 1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931946e-23, 1.931948e-23, 1.931947e-23, 1.931949e-23, 1.931949e-23, 
    1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931944e-23, 1.931947e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.93195e-23, 1.931948e-23, 
    1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931949e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931947e-23, 1.931949e-23, 1.931947e-23, 1.931949e-23, 1.931949e-23, 
    1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931948e-23, 1.931948e-23, 1.931948e-23, 1.931948e-23, 1.931949e-23, 
    1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931946e-23, 1.931946e-23, 1.931945e-23, 1.931945e-23, 1.931944e-23, 
    1.931945e-23, 1.931943e-23, 1.931947e-23, 1.931945e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 
    1.931948e-23, 1.931949e-23, 1.931949e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931946e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931941e-23, 1.931941e-23, 1.931941e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975388e-24, 1.975386e-24, 1.975387e-24, 1.975385e-24, 1.975386e-24, 
    1.975385e-24, 1.975387e-24, 1.975386e-24, 1.975387e-24, 1.975388e-24, 
    1.975383e-24, 1.975385e-24, 1.975381e-24, 1.975382e-24, 1.975379e-24, 
    1.975381e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 
    1.975376e-24, 1.975377e-24, 1.975375e-24, 1.975376e-24, 1.975376e-24, 
    1.975378e-24, 1.975385e-24, 1.975384e-24, 1.975385e-24, 1.975385e-24, 
    1.975385e-24, 1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975385e-24, 1.975385e-24, 1.975384e-24, 1.975384e-24, 
    1.975382e-24, 1.975383e-24, 1.97538e-24, 1.97538e-24, 1.975378e-24, 
    1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975383e-24, 1.975382e-24, 1.975384e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975385e-24, 1.975384e-24, 1.975384e-24, 
    1.975382e-24, 1.975381e-24, 1.975379e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 1.975379e-24, 
    1.975378e-24, 1.97538e-24, 1.975379e-24, 1.975384e-24, 1.975385e-24, 
    1.975386e-24, 1.975386e-24, 1.975388e-24, 1.975387e-24, 1.975387e-24, 
    1.975386e-24, 1.975386e-24, 1.975386e-24, 1.975384e-24, 1.975385e-24, 
    1.975381e-24, 1.975383e-24, 1.975379e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975379e-24, 1.975377e-24, 1.975377e-24, 
    1.975377e-24, 1.975376e-24, 1.975379e-24, 1.975378e-24, 1.975386e-24, 
    1.975386e-24, 1.975386e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.97538e-24, 1.975377e-24, 
    1.975379e-24, 1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975386e-24, 1.975386e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975385e-24, 1.975385e-24, 1.975384e-24, 
    1.975384e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 
    1.975378e-24, 1.975379e-24, 1.975377e-24, 1.975377e-24, 1.975377e-24, 
    1.975377e-24, 1.975386e-24, 1.975386e-24, 1.975386e-24, 1.975386e-24, 
    1.975386e-24, 1.975384e-24, 1.975384e-24, 1.975382e-24, 1.975383e-24, 
    1.975381e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.975383e-24, 
    1.97538e-24, 1.975382e-24, 1.975379e-24, 1.97538e-24, 1.975378e-24, 
    1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975377e-24, 1.975376e-24, 
    1.975376e-24, 1.975375e-24, 1.975385e-24, 1.975384e-24, 1.975384e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975382e-24, 1.975381e-24, 1.975384e-24, 
    1.975384e-24, 1.975384e-24, 1.975385e-24, 1.975381e-24, 1.975383e-24, 
    1.97538e-24, 1.975381e-24, 1.975378e-24, 1.975379e-24, 1.975376e-24, 
    1.975375e-24, 1.975374e-24, 1.975372e-24, 1.975384e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.97538e-24, 1.975379e-24, 1.97538e-24, 1.975379e-24, 
    1.975383e-24, 1.975381e-24, 1.975385e-24, 1.975384e-24, 1.975383e-24, 
    1.975383e-24, 1.975381e-24, 1.975381e-24, 1.975379e-24, 1.97538e-24, 
    1.975375e-24, 1.975378e-24, 1.975371e-24, 1.975373e-24, 1.975385e-24, 
    1.975384e-24, 1.975382e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975378e-24, 1.975381e-24, 1.97538e-24, 1.975382e-24, 1.975382e-24, 
    1.975382e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.97538e-24, 1.975375e-24, 1.975379e-24, 
    1.975384e-24, 1.975382e-24, 1.975382e-24, 1.975383e-24, 1.97538e-24, 
    1.975381e-24, 1.975378e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.97538e-24, 1.975381e-24, 1.975382e-24, 
    1.975383e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975381e-24, 1.975379e-24, 1.97538e-24, 
    1.975379e-24, 1.975381e-24, 1.975379e-24, 1.975382e-24, 1.975382e-24, 
    1.975381e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.97538e-24, 1.97538e-24, 1.975381e-24, 1.975381e-24, 1.975382e-24, 
    1.975382e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 1.975379e-24, 
    1.975378e-24, 1.975377e-24, 1.975376e-24, 1.975377e-24, 1.975375e-24, 
    1.975377e-24, 1.975374e-24, 1.975379e-24, 1.975377e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975378e-24, 
    1.97538e-24, 1.975382e-24, 1.975382e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.975381e-24, 1.975382e-24, 1.97538e-24, 1.975381e-24, 
    1.975379e-24, 1.975378e-24, 1.975375e-24, 1.975374e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24 ;

 CONC_CH4_SAT =
  3.522518e-08, 3.522421e-08, 3.522441e-08, 3.522359e-08, 3.522406e-08, 
    3.52235e-08, 3.522501e-08, 3.522415e-08, 3.522472e-08, 3.522512e-08, 
    3.522185e-08, 3.522355e-08, 3.522016e-08, 3.522129e-08, 3.521843e-08, 
    3.522031e-08, 3.521805e-08, 3.521853e-08, 3.521717e-08, 3.521757e-08, 
    3.511421e-08, 3.521699e-08, 3.511297e-08, 3.511466e-08, 3.511437e-08, 
    3.521702e-08, 3.522326e-08, 3.522205e-08, 3.522332e-08, 3.522315e-08, 
    3.522323e-08, 3.522404e-08, 3.522441e-08, 3.522529e-08, 3.522514e-08, 
    3.522451e-08, 3.522308e-08, 3.52236e-08, 3.522235e-08, 3.522238e-08, 
    3.522089e-08, 3.522157e-08, 3.5219e-08, 3.521976e-08, 3.521755e-08, 
    3.521811e-08, 3.521757e-08, 3.521774e-08, 3.521757e-08, 3.521839e-08, 
    3.521804e-08, 3.521877e-08, 3.522144e-08, 3.522066e-08, 3.52229e-08, 
    3.522409e-08, 3.522496e-08, 3.522554e-08, 3.522546e-08, 3.522529e-08, 
    3.52245e-08, 3.522377e-08, 3.522318e-08, 3.522278e-08, 3.522239e-08, 
    3.522103e-08, 3.522038e-08, 3.521882e-08, 3.521914e-08, 3.521862e-08, 
    3.521817e-08, 3.521735e-08, 3.521749e-08, 3.521712e-08, 3.521866e-08, 
    3.521763e-08, 3.521932e-08, 3.521886e-08, 3.522213e-08, 3.522347e-08, 
    3.522389e-08, 3.522437e-08, 3.522539e-08, 3.522468e-08, 3.522496e-08, 
    3.522432e-08, 3.522389e-08, 3.522411e-08, 3.522277e-08, 3.522329e-08, 
    3.522035e-08, 3.522166e-08, 3.521822e-08, 3.521908e-08, 3.521802e-08, 
    3.521857e-08, 3.521761e-08, 3.521848e-08, 3.521699e-08, 3.511561e-08, 
    3.521687e-08, 3.511462e-08, 3.521852e-08, 3.521756e-08, 3.522411e-08, 
    3.522407e-08, 3.522392e-08, 3.522459e-08, 3.522464e-08, 3.522528e-08, 
    3.522473e-08, 3.522447e-08, 3.522388e-08, 3.522349e-08, 3.522313e-08, 
    3.522232e-08, 3.522136e-08, 3.522e-08, 3.521902e-08, 3.521835e-08, 
    3.521877e-08, 3.52184e-08, 3.521881e-08, 3.521901e-08, 3.511585e-08, 
    3.521803e-08, 3.51148e-08, 3.511496e-08, 3.52171e-08, 3.511494e-08, 
    3.522405e-08, 3.522426e-08, 3.522492e-08, 3.52244e-08, 3.522536e-08, 
    3.522481e-08, 3.522448e-08, 3.522325e-08, 3.522301e-08, 3.522274e-08, 
    3.522223e-08, 3.522154e-08, 3.522028e-08, 3.521917e-08, 3.521815e-08, 
    3.521823e-08, 3.52182e-08, 3.521795e-08, 3.521854e-08, 3.521786e-08, 
    3.521773e-08, 3.521804e-08, 3.511498e-08, 3.511585e-08, 3.511496e-08, 
    3.511549e-08, 3.522419e-08, 3.522385e-08, 3.522403e-08, 3.522368e-08, 
    3.522392e-08, 3.52228e-08, 3.522245e-08, 3.522083e-08, 3.522155e-08, 
    3.522044e-08, 3.522145e-08, 3.522126e-08, 3.522034e-08, 3.52214e-08, 
    3.521921e-08, 3.522065e-08, 3.521794e-08, 3.521938e-08, 3.521785e-08, 
    3.521815e-08, 3.521766e-08, 3.52172e-08, 3.511557e-08, 3.511398e-08, 
    3.511433e-08, 3.511312e-08, 3.522334e-08, 3.522287e-08, 3.522294e-08, 
    3.522246e-08, 3.522209e-08, 3.522131e-08, 3.521998e-08, 3.522049e-08, 
    3.521957e-08, 3.521937e-08, 3.522079e-08, 3.52199e-08, 3.522257e-08, 
    3.522213e-08, 3.522241e-08, 3.522329e-08, 3.522034e-08, 3.522187e-08, 
    3.5219e-08, 3.521988e-08, 3.521726e-08, 3.521856e-08, 3.511452e-08, 
    3.511291e-08, 3.511157e-08, 3.510991e-08, 3.522264e-08, 3.522296e-08, 
    3.522241e-08, 3.522157e-08, 3.522085e-08, 3.521983e-08, 3.521973e-08, 
    3.521953e-08, 3.521903e-08, 3.521859e-08, 3.521944e-08, 3.521848e-08, 
    3.522197e-08, 3.522021e-08, 3.522306e-08, 3.522219e-08, 3.522164e-08, 
    3.522191e-08, 3.522056e-08, 3.522022e-08, 3.521881e-08, 3.521956e-08, 
    3.511328e-08, 3.521706e-08, 3.510873e-08, 3.511069e-08, 3.522307e-08, 
    3.522266e-08, 3.522113e-08, 3.522187e-08, 3.521977e-08, 3.521922e-08, 
    3.521879e-08, 3.52182e-08, 3.521815e-08, 3.521779e-08, 3.521837e-08, 
    3.521783e-08, 3.521982e-08, 3.521895e-08, 3.522134e-08, 3.522076e-08, 
    3.522103e-08, 3.522132e-08, 3.522043e-08, 3.521942e-08, 3.521944e-08, 
    3.52191e-08, 3.521806e-08, 3.521976e-08, 3.511287e-08, 3.521779e-08, 
    3.522219e-08, 3.522131e-08, 3.522123e-08, 3.522157e-08, 3.521928e-08, 
    3.522012e-08, 3.521781e-08, 3.521846e-08, 3.52174e-08, 3.521793e-08, 
    3.5218e-08, 3.521867e-08, 3.521907e-08, 3.522007e-08, 3.522088e-08, 
    3.522153e-08, 3.522138e-08, 3.522067e-08, 3.521937e-08, 3.521813e-08, 
    3.52184e-08, 3.521749e-08, 3.521993e-08, 3.52189e-08, 3.521928e-08, 
    3.521828e-08, 3.522049e-08, 3.521848e-08, 3.522098e-08, 3.522078e-08, 
    3.522014e-08, 3.52188e-08, 3.521856e-08, 3.521822e-08, 3.521844e-08, 
    3.521934e-08, 3.521951e-08, 3.522016e-08, 3.522032e-08, 3.522083e-08, 
    3.522122e-08, 3.522085e-08, 3.522045e-08, 3.521936e-08, 3.521832e-08, 
    3.521718e-08, 3.521692e-08, 3.511387e-08, 3.511558e-08, 3.511284e-08, 
    3.511504e-08, 3.511139e-08, 3.521843e-08, 3.511517e-08, 3.522012e-08, 
    3.521974e-08, 3.521899e-08, 3.521733e-08, 3.521828e-08, 3.521718e-08, 
    3.521951e-08, 3.522062e-08, 3.522095e-08, 3.522148e-08, 3.522094e-08, 
    3.522099e-08, 3.522046e-08, 3.522063e-08, 3.521932e-08, 3.522004e-08, 
    3.521799e-08, 3.521721e-08, 3.511323e-08, 3.511146e-08, 3.510974e-08, 
    3.510896e-08, 3.510873e-08, 3.510863e-08,
  6.096772e-11, 6.10464e-11, 6.103116e-11, 6.109448e-11, 6.105943e-11, 
    6.110083e-11, 6.098376e-11, 6.104946e-11, 6.100757e-11, 6.097492e-11, 
    6.121701e-11, 6.109733e-11, 6.135022e-11, 6.126701e-11, 6.147609e-11, 
    6.133717e-11, 6.150409e-11, 6.147226e-11, 6.156847e-11, 6.154093e-11, 
    6.14207e-11, 6.158117e-11, 6.148339e-11, 6.140151e-11, 6.141423e-11, 
    6.157842e-11, 6.112159e-11, 6.120206e-11, 6.111679e-11, 6.112828e-11, 
    6.112316e-11, 6.106009e-11, 6.102818e-11, 6.096183e-11, 6.097391e-11, 
    6.10227e-11, 6.113345e-11, 6.109598e-11, 6.11907e-11, 6.118857e-11, 
    6.129776e-11, 6.124635e-11, 6.143874e-11, 6.138407e-11, 6.154208e-11, 
    6.150235e-11, 6.154019e-11, 6.152874e-11, 6.154034e-11, 6.148206e-11, 
    6.150703e-11, 6.145578e-11, 6.12557e-11, 6.131451e-11, 6.114809e-11, 
    6.105083e-11, 6.098661e-11, 6.094088e-11, 6.094734e-11, 6.095963e-11, 
    6.102299e-11, 6.108265e-11, 6.112805e-11, 6.115837e-11, 6.118826e-11, 
    6.128082e-11, 6.133309e-11, 6.14497e-11, 6.142882e-11, 6.146431e-11, 
    6.14984e-11, 6.155541e-11, 6.154605e-11, 6.157112e-11, 6.146348e-11, 
    6.153498e-11, 6.141689e-11, 6.144919e-11, 6.119578e-11, 6.110612e-11, 
    6.106746e-11, 6.103407e-11, 6.095231e-11, 6.100875e-11, 6.098649e-11, 
    6.103956e-11, 6.107317e-11, 6.105658e-11, 6.11592e-11, 6.111929e-11, 
    6.133619e-11, 6.123875e-11, 6.149443e-11, 6.143312e-11, 6.150914e-11, 
    6.147039e-11, 6.153672e-11, 6.147702e-11, 6.15805e-11, 6.136153e-11, 
    6.158759e-11, 6.140425e-11, 6.14737e-11, 6.154013e-11, 6.105608e-11, 
    6.105878e-11, 6.107145e-11, 6.101575e-11, 6.101237e-11, 6.096147e-11, 
    6.100682e-11, 6.102607e-11, 6.107517e-11, 6.110409e-11, 6.113161e-11, 
    6.119209e-11, 6.126038e-11, 6.136321e-11, 6.143709e-11, 6.148655e-11, 
    6.145626e-11, 6.148299e-11, 6.145309e-11, 6.14391e-11, 6.13534e-11, 
    6.150722e-11, 6.139592e-11, 6.138885e-11, 6.157169e-11, 6.138965e-11, 
    6.106069e-11, 6.104511e-11, 6.09908e-11, 6.103331e-11, 6.095593e-11, 
    6.099918e-11, 6.102399e-11, 6.112e-11, 6.114122e-11, 6.116071e-11, 
    6.119932e-11, 6.124878e-11, 6.134317e-11, 6.142537e-11, 6.150042e-11, 
    6.149493e-11, 6.149686e-11, 6.151354e-11, 6.147211e-11, 6.152035e-11, 
    6.152839e-11, 6.150729e-11, 6.13879e-11, 6.135385e-11, 6.13887e-11, 
    6.136647e-11, 6.105019e-11, 6.107644e-11, 6.106225e-11, 6.108889e-11, 
    6.107007e-11, 6.115355e-11, 6.117856e-11, 6.129983e-11, 6.124777e-11, 
    6.133086e-11, 6.125611e-11, 6.126933e-11, 6.133332e-11, 6.126019e-11, 
    6.142072e-11, 6.13117e-11, 6.15142e-11, 6.140522e-11, 6.1521e-11, 
    6.150009e-11, 6.153478e-11, 6.156576e-11, 6.136334e-11, 6.143369e-11, 
    6.141736e-11, 6.147655e-11, 6.11156e-11, 6.114955e-11, 6.114667e-11, 
    6.118227e-11, 6.120857e-11, 6.126711e-11, 6.136672e-11, 6.132932e-11, 
    6.13981e-11, 6.141186e-11, 6.130742e-11, 6.137146e-11, 6.117235e-11, 
    6.120281e-11, 6.118476e-11, 6.111821e-11, 6.133778e-11, 6.122154e-11, 
    6.143829e-11, 6.137409e-11, 6.156133e-11, 6.146815e-11, 6.140836e-11, 
    6.148482e-11, 6.155738e-11, 6.164167e-11, 6.11682e-11, 6.114512e-11, 
    6.118654e-11, 6.12436e-11, 6.130109e-11, 6.137798e-11, 6.13859e-11, 
    6.140027e-11, 6.143759e-11, 6.14689e-11, 6.140469e-11, 6.147676e-11, 
    6.120964e-11, 6.134813e-11, 6.113629e-11, 6.119753e-11, 6.124028e-11, 
    6.122165e-11, 6.132507e-11, 6.134998e-11, 6.145107e-11, 6.13989e-11, 
    6.146584e-11, 6.157214e-11, 6.17062e-11, 6.160115e-11, 6.113703e-11, 
    6.116817e-11, 6.127872e-11, 6.122489e-11, 6.138317e-11, 6.142258e-11, 
    6.14547e-11, 6.149554e-11, 6.150003e-11, 6.152424e-11, 6.148456e-11, 
    6.152272e-11, 6.137815e-11, 6.14428e-11, 6.126538e-11, 6.130854e-11, 
    6.128873e-11, 6.126691e-11, 6.133422e-11, 6.140568e-11, 6.140739e-11, 
    6.143025e-11, 6.149431e-11, 6.138382e-11, 6.148297e-11, 6.151481e-11, 
    6.120211e-11, 6.12629e-11, 6.127241e-11, 6.124738e-11, 6.141862e-11, 
    6.135652e-11, 6.152368e-11, 6.147858e-11, 6.15525e-11, 6.151576e-11, 
    6.151035e-11, 6.146317e-11, 6.143373e-11, 6.135933e-11, 6.12988e-11, 
    6.125085e-11, 6.126202e-11, 6.131468e-11, 6.141009e-11, 6.150036e-11, 
    6.148057e-11, 6.154689e-11, 6.137154e-11, 6.144502e-11, 6.141657e-11, 
    6.149077e-11, 6.132828e-11, 6.146612e-11, 6.129294e-11, 6.130818e-11, 
    6.135529e-11, 6.144988e-11, 6.147106e-11, 6.149335e-11, 6.147964e-11, 
    6.141254e-11, 6.140163e-11, 6.135419e-11, 6.134099e-11, 6.130488e-11, 
    6.127487e-11, 6.130224e-11, 6.133093e-11, 6.141265e-11, 6.148611e-11, 
    6.156618e-11, 6.158583e-11, 6.143577e-11, 6.136152e-11, 6.14841e-11, 
    6.137943e-11, 6.156106e-11, 6.147437e-11, 6.137667e-11, 6.13575e-11, 
    6.13857e-11, 6.143649e-11, 6.155323e-11, 6.149042e-11, 6.156396e-11, 
    6.140122e-11, 6.13164e-11, 6.129467e-11, 6.125373e-11, 6.129561e-11, 
    6.129221e-11, 6.133225e-11, 6.13194e-11, 6.141537e-11, 6.136384e-11, 
    6.151016e-11, 6.156343e-11, 6.147028e-11, 6.156101e-11, 6.165369e-11, 
    6.169452e-11, 6.170696e-11, 6.171214e-11,
  2.833864e-14, 2.840811e-14, 2.839463e-14, 2.845063e-14, 2.841961e-14, 
    2.845624e-14, 2.835277e-14, 2.841081e-14, 2.837379e-14, 2.834497e-14, 
    2.855925e-14, 2.845314e-14, 2.867521e-14, 2.860317e-14, 2.87844e-14, 
    2.866391e-14, 2.880873e-14, 2.878105e-14, 2.88647e-14, 2.884074e-14, 
    2.882827e-14, 2.887576e-14, 2.888325e-14, 2.881141e-14, 2.882259e-14, 
    2.887338e-14, 2.847461e-14, 2.854599e-14, 2.847035e-14, 2.848053e-14, 
    2.847599e-14, 2.84202e-14, 2.839202e-14, 2.833342e-14, 2.834408e-14, 
    2.838717e-14, 2.848511e-14, 2.845193e-14, 2.853583e-14, 2.853394e-14, 
    2.862976e-14, 2.858522e-14, 2.875194e-14, 2.870451e-14, 2.884174e-14, 
    2.880719e-14, 2.88401e-14, 2.883014e-14, 2.884023e-14, 2.878957e-14, 
    2.881126e-14, 2.876674e-14, 2.859339e-14, 2.864427e-14, 2.849807e-14, 
    2.841205e-14, 2.83553e-14, 2.831495e-14, 2.832065e-14, 2.83315e-14, 
    2.838742e-14, 2.844014e-14, 2.848031e-14, 2.850717e-14, 2.853367e-14, 
    2.861515e-14, 2.866037e-14, 2.876147e-14, 2.874333e-14, 2.877415e-14, 
    2.880376e-14, 2.885334e-14, 2.88452e-14, 2.886702e-14, 2.877342e-14, 
    2.883558e-14, 2.873297e-14, 2.876101e-14, 2.854043e-14, 2.846091e-14, 
    2.842675e-14, 2.83972e-14, 2.832503e-14, 2.837484e-14, 2.835519e-14, 
    2.840204e-14, 2.843176e-14, 2.841708e-14, 2.850791e-14, 2.847257e-14, 
    2.866305e-14, 2.857849e-14, 2.880031e-14, 2.874706e-14, 2.881309e-14, 
    2.877941e-14, 2.883709e-14, 2.878518e-14, 2.887518e-14, 2.877627e-14, 
    2.888136e-14, 2.881381e-14, 2.878229e-14, 2.884005e-14, 2.841664e-14, 
    2.841904e-14, 2.843023e-14, 2.838102e-14, 2.837804e-14, 2.83331e-14, 
    2.837313e-14, 2.839014e-14, 2.843352e-14, 2.845911e-14, 2.848347e-14, 
    2.853707e-14, 2.859744e-14, 2.868645e-14, 2.875051e-14, 2.879345e-14, 
    2.876715e-14, 2.879037e-14, 2.876439e-14, 2.875224e-14, 2.876908e-14, 
    2.881144e-14, 2.88065e-14, 2.880029e-14, 2.886752e-14, 2.880099e-14, 
    2.842072e-14, 2.840695e-14, 2.835899e-14, 2.839652e-14, 2.832822e-14, 
    2.836639e-14, 2.838831e-14, 2.847321e-14, 2.849198e-14, 2.850925e-14, 
    2.854348e-14, 2.858738e-14, 2.866909e-14, 2.874035e-14, 2.880551e-14, 
    2.880074e-14, 2.880241e-14, 2.881693e-14, 2.878092e-14, 2.882284e-14, 
    2.882984e-14, 2.881148e-14, 2.879946e-14, 2.876948e-14, 2.880016e-14, 
    2.878061e-14, 2.841143e-14, 2.843464e-14, 2.842209e-14, 2.844567e-14, 
    2.842902e-14, 2.850293e-14, 2.85251e-14, 2.863157e-14, 2.858649e-14, 
    2.865843e-14, 2.859374e-14, 2.860517e-14, 2.866059e-14, 2.859726e-14, 
    2.873633e-14, 2.864186e-14, 2.881749e-14, 2.87229e-14, 2.882341e-14, 
    2.880522e-14, 2.883538e-14, 2.886235e-14, 2.877786e-14, 2.883965e-14, 
    2.882533e-14, 2.887724e-14, 2.846929e-14, 2.849938e-14, 2.849681e-14, 
    2.852836e-14, 2.855169e-14, 2.860324e-14, 2.868948e-14, 2.865707e-14, 
    2.871668e-14, 2.872861e-14, 2.863812e-14, 2.869359e-14, 2.851958e-14, 
    2.85466e-14, 2.853057e-14, 2.847162e-14, 2.866443e-14, 2.856322e-14, 
    2.875155e-14, 2.869586e-14, 2.88585e-14, 2.87775e-14, 2.881743e-14, 
    2.888451e-14, 2.894815e-14, 2.902222e-14, 2.851589e-14, 2.849543e-14, 
    2.853214e-14, 2.85828e-14, 2.863264e-14, 2.869924e-14, 2.87061e-14, 
    2.871856e-14, 2.875094e-14, 2.877813e-14, 2.872242e-14, 2.878495e-14, 
    2.85527e-14, 2.867338e-14, 2.848763e-14, 2.854192e-14, 2.857985e-14, 
    2.85633e-14, 2.865339e-14, 2.867497e-14, 2.876266e-14, 2.871737e-14, 
    2.886787e-14, 2.886793e-14, 2.907893e-14, 2.898661e-14, 2.848827e-14, 
    2.851586e-14, 2.86133e-14, 2.856617e-14, 2.870373e-14, 2.873791e-14, 
    2.876578e-14, 2.880128e-14, 2.880518e-14, 2.882623e-14, 2.879173e-14, 
    2.88249e-14, 2.869938e-14, 2.875547e-14, 2.860175e-14, 2.863909e-14, 
    2.862194e-14, 2.860307e-14, 2.866131e-14, 2.872327e-14, 2.872473e-14, 
    2.874458e-14, 2.88003e-14, 2.87043e-14, 2.888293e-14, 2.881811e-14, 
    2.854595e-14, 2.859963e-14, 2.860783e-14, 2.858613e-14, 2.873448e-14, 
    2.868064e-14, 2.882573e-14, 2.878653e-14, 2.885081e-14, 2.881885e-14, 
    2.881414e-14, 2.877315e-14, 2.874759e-14, 2.868308e-14, 2.863066e-14, 
    2.858918e-14, 2.859884e-14, 2.864441e-14, 2.87271e-14, 2.880547e-14, 
    2.878828e-14, 2.884592e-14, 2.869365e-14, 2.87574e-14, 2.873271e-14, 
    2.879713e-14, 2.865618e-14, 2.877578e-14, 2.862558e-14, 2.863877e-14, 
    2.867957e-14, 2.876164e-14, 2.878e-14, 2.879937e-14, 2.878745e-14, 
    2.872922e-14, 2.871974e-14, 2.867861e-14, 2.866719e-14, 2.863591e-14, 
    2.860995e-14, 2.863364e-14, 2.865848e-14, 2.87293e-14, 2.879309e-14, 
    2.886272e-14, 2.887982e-14, 2.88415e-14, 2.877626e-14, 2.888392e-14, 
    2.879206e-14, 2.895144e-14, 2.878292e-14, 2.878961e-14, 2.868147e-14, 
    2.870592e-14, 2.875001e-14, 2.885148e-14, 2.879683e-14, 2.886081e-14, 
    2.871938e-14, 2.864592e-14, 2.862708e-14, 2.859168e-14, 2.862789e-14, 
    2.862495e-14, 2.865961e-14, 2.864848e-14, 2.873166e-14, 2.868697e-14, 
    2.881399e-14, 2.886034e-14, 2.887174e-14, 2.895136e-14, 2.903275e-14, 
    2.906865e-14, 2.907959e-14, 2.908416e-14,
  3.913097e-18, 3.92695e-18, 3.92426e-18, 3.93544e-18, 3.929244e-18, 
    3.936562e-18, 3.915913e-18, 3.927492e-18, 3.920103e-18, 3.914356e-18, 
    3.957168e-18, 3.935942e-18, 3.979898e-18, 3.965868e-18, 4.001198e-18, 
    3.977699e-18, 4.00595e-18, 4.000542e-18, 4.016889e-18, 4.012203e-18, 
    4.016815e-18, 4.019053e-18, 4.027611e-18, 4.013502e-18, 4.015697e-18, 
    4.018586e-18, 3.940229e-18, 3.954514e-18, 3.939379e-18, 3.941415e-18, 
    3.940506e-18, 3.929364e-18, 3.923742e-18, 3.912055e-18, 3.914179e-18, 
    3.922773e-18, 3.942331e-18, 3.935699e-18, 3.952471e-18, 3.952092e-18, 
    3.971045e-18, 3.962359e-18, 3.994859e-18, 3.985606e-18, 4.012399e-18, 
    4.005648e-18, 4.012078e-18, 4.01013e-18, 4.012103e-18, 4.002205e-18, 
    4.006443e-18, 3.997747e-18, 3.963966e-18, 3.973869e-18, 3.944921e-18, 
    3.927742e-18, 3.916416e-18, 3.908375e-18, 3.909511e-18, 3.911673e-18, 
    3.922822e-18, 3.933344e-18, 3.941368e-18, 3.946738e-18, 3.952038e-18, 
    3.968205e-18, 3.977007e-18, 3.996721e-18, 3.993178e-18, 3.999196e-18, 
    4.004977e-18, 4.014668e-18, 4.013075e-18, 4.017343e-18, 3.999051e-18, 
    4.011196e-18, 3.991157e-18, 3.996629e-18, 3.953402e-18, 3.937491e-18, 
    3.930675e-18, 3.924774e-18, 3.910383e-18, 3.920313e-18, 3.916395e-18, 
    3.925737e-18, 3.931671e-18, 3.928739e-18, 3.946885e-18, 3.939821e-18, 
    3.977529e-18, 3.961012e-18, 4.004303e-18, 3.993907e-18, 4.0068e-18, 
    4.000222e-18, 4.01149e-18, 4.001348e-18, 4.018939e-18, 4.006597e-18, 
    4.020149e-18, 4.013972e-18, 4.000784e-18, 4.01207e-18, 3.928653e-18, 
    3.92913e-18, 3.931365e-18, 3.921547e-18, 3.920951e-18, 3.911993e-18, 
    3.91997e-18, 3.923365e-18, 3.932021e-18, 3.937132e-18, 3.942001e-18, 
    3.95272e-18, 3.964755e-18, 3.982088e-18, 3.99458e-18, 4.002963e-18, 
    3.997826e-18, 4.00236e-18, 3.997289e-18, 3.994917e-18, 4.005182e-18, 
    4.006478e-18, 4.012536e-18, 4.011316e-18, 4.017442e-18, 4.011454e-18, 
    3.929467e-18, 3.926717e-18, 3.917152e-18, 3.924636e-18, 3.911019e-18, 
    3.918628e-18, 3.923001e-18, 3.939951e-18, 3.943701e-18, 3.947155e-18, 
    3.954002e-18, 3.962791e-18, 3.978704e-18, 3.992597e-18, 4.005317e-18, 
    4.004386e-18, 4.004713e-18, 4.007549e-18, 4.000515e-18, 4.008705e-18, 
    4.010074e-18, 4.006485e-18, 4.011153e-18, 4.00526e-18, 4.01129e-18, 
    4.007449e-18, 3.927612e-18, 3.932245e-18, 3.92974e-18, 3.934448e-18, 
    3.931125e-18, 3.945893e-18, 3.950328e-18, 3.971399e-18, 3.962613e-18, 
    3.976629e-18, 3.964033e-18, 3.966258e-18, 3.977053e-18, 3.964718e-18, 
    3.991816e-18, 3.973403e-18, 4.00766e-18, 3.989197e-18, 4.008816e-18, 
    4.005262e-18, 4.011156e-18, 4.01643e-18, 4.00691e-18, 4.019047e-18, 
    4.016234e-18, 4.026429e-18, 3.939166e-18, 3.945182e-18, 3.944666e-18, 
    3.950977e-18, 3.955646e-18, 3.965882e-18, 3.982678e-18, 3.976362e-18, 
    3.987978e-18, 3.990308e-18, 3.97267e-18, 3.98348e-18, 3.949222e-18, 
    3.95463e-18, 3.95142e-18, 3.939633e-18, 3.977796e-18, 3.957957e-18, 
    3.994783e-18, 3.983921e-18, 4.015676e-18, 3.99985e-18, 4.014683e-18, 
    4.027862e-18, 4.040367e-18, 4.054943e-18, 3.948483e-18, 3.944391e-18, 
    3.951732e-18, 3.961877e-18, 3.971605e-18, 3.98458e-18, 3.985917e-18, 
    3.988346e-18, 3.994662e-18, 3.99997e-18, 3.9891e-18, 4.001303e-18, 
    3.955856e-18, 3.979542e-18, 3.942832e-18, 3.953694e-18, 3.961285e-18, 
    3.957969e-18, 3.975644e-18, 3.979848e-18, 3.996952e-18, 3.988113e-18, 
    4.024592e-18, 4.017524e-18, 4.066113e-18, 4.047934e-18, 3.942959e-18, 
    3.948476e-18, 3.967841e-18, 3.958545e-18, 3.985455e-18, 3.992122e-18, 
    3.99756e-18, 4.004494e-18, 4.005254e-18, 4.009368e-18, 4.002626e-18, 
    4.009107e-18, 3.984607e-18, 3.995547e-18, 3.965591e-18, 3.97286e-18, 
    3.96952e-18, 3.965847e-18, 3.977188e-18, 3.989268e-18, 3.98955e-18, 
    3.993424e-18, 4.00431e-18, 3.985565e-18, 4.027555e-18, 4.007789e-18, 
    3.954496e-18, 3.965182e-18, 3.966776e-18, 3.96254e-18, 3.991453e-18, 
    3.980954e-18, 4.00927e-18, 4.001611e-18, 4.014172e-18, 4.007925e-18, 
    4.007006e-18, 3.998998e-18, 3.99401e-18, 3.981431e-18, 3.97122e-18, 
    3.963146e-18, 3.965024e-18, 3.973897e-18, 3.990013e-18, 4.005312e-18, 
    4.001954e-18, 4.013217e-18, 3.983489e-18, 3.995926e-18, 3.991108e-18, 
    4.003682e-18, 3.976189e-18, 3.999521e-18, 3.97023e-18, 3.972798e-18, 
    3.980746e-18, 3.996754e-18, 4.000337e-18, 4.004121e-18, 4.001791e-18, 
    3.990427e-18, 3.988578e-18, 3.980559e-18, 3.978335e-18, 3.97224e-18, 
    3.967188e-18, 3.971798e-18, 3.976638e-18, 3.990442e-18, 4.002892e-18, 
    4.016502e-18, 4.019846e-18, 4.019415e-18, 4.006598e-18, 4.027751e-18, 
    4.009708e-18, 4.04102e-18, 4.000911e-18, 4.009222e-18, 3.981116e-18, 
    3.985881e-18, 3.994484e-18, 4.014306e-18, 4.003623e-18, 4.016131e-18, 
    3.988507e-18, 3.974191e-18, 3.970522e-18, 3.963632e-18, 3.97068e-18, 
    3.970107e-18, 3.976855e-18, 3.974687e-18, 3.990901e-18, 3.982188e-18, 
    4.006976e-18, 4.016038e-18, 4.025351e-18, 4.041e-18, 4.057014e-18, 
    4.064086e-18, 4.066242e-18, 4.067142e-18,
  1.685924e-22, 1.693935e-22, 1.692378e-22, 1.69885e-22, 1.695261e-22, 
    1.699499e-22, 1.68755e-22, 1.694249e-22, 1.689973e-22, 1.686651e-22, 
    1.71145e-22, 1.69914e-22, 1.724785e-22, 1.716502e-22, 1.73738e-22, 
    1.723488e-22, 1.740193e-22, 1.736989e-22, 1.746671e-22, 1.743894e-22, 
    1.749556e-22, 1.747954e-22, 1.755979e-22, 1.747583e-22, 1.748889e-22, 
    1.747678e-22, 1.701622e-22, 1.70991e-22, 1.70113e-22, 1.70231e-22, 
    1.701783e-22, 1.695331e-22, 1.692081e-22, 1.68532e-22, 1.686548e-22, 
    1.691518e-22, 1.702841e-22, 1.698998e-22, 1.708717e-22, 1.708498e-22, 
    1.719555e-22, 1.714456e-22, 1.733627e-22, 1.728155e-22, 1.74401e-22, 
    1.740011e-22, 1.74382e-22, 1.742666e-22, 1.743835e-22, 1.737974e-22, 
    1.740483e-22, 1.735335e-22, 1.71538e-22, 1.721223e-22, 1.704341e-22, 
    1.694396e-22, 1.687842e-22, 1.683195e-22, 1.683851e-22, 1.685101e-22, 
    1.691547e-22, 1.697634e-22, 1.702281e-22, 1.705394e-22, 1.708466e-22, 
    1.717885e-22, 1.723078e-22, 1.734729e-22, 1.732632e-22, 1.736193e-22, 
    1.739614e-22, 1.745356e-22, 1.744411e-22, 1.746942e-22, 1.736106e-22, 
    1.743299e-22, 1.731436e-22, 1.734673e-22, 1.709265e-22, 1.700036e-22, 
    1.696093e-22, 1.692675e-22, 1.684355e-22, 1.690096e-22, 1.68783e-22, 
    1.693231e-22, 1.696665e-22, 1.694968e-22, 1.705479e-22, 1.701385e-22, 
    1.723386e-22, 1.713675e-22, 1.739215e-22, 1.733063e-22, 1.740694e-22, 
    1.736799e-22, 1.743473e-22, 1.737465e-22, 1.747888e-22, 1.743474e-22, 
    1.748606e-22, 1.747861e-22, 1.737132e-22, 1.743817e-22, 1.694919e-22, 
    1.695195e-22, 1.696488e-22, 1.690809e-22, 1.690464e-22, 1.685285e-22, 
    1.689896e-22, 1.69186e-22, 1.696867e-22, 1.699828e-22, 1.702648e-22, 
    1.708863e-22, 1.715846e-22, 1.726077e-22, 1.733461e-22, 1.738421e-22, 
    1.735381e-22, 1.738064e-22, 1.735063e-22, 1.733659e-22, 1.742632e-22, 
    1.740504e-22, 1.747007e-22, 1.746281e-22, 1.747001e-22, 1.746363e-22, 
    1.69539e-22, 1.693798e-22, 1.688267e-22, 1.692594e-22, 1.684722e-22, 
    1.68912e-22, 1.691651e-22, 1.701463e-22, 1.703633e-22, 1.705636e-22, 
    1.709606e-22, 1.714706e-22, 1.724078e-22, 1.732289e-22, 1.739815e-22, 
    1.739264e-22, 1.739457e-22, 1.741138e-22, 1.736973e-22, 1.741823e-22, 
    1.742634e-22, 1.740507e-22, 1.746184e-22, 1.742677e-22, 1.746266e-22, 
    1.74398e-22, 1.694316e-22, 1.696998e-22, 1.695548e-22, 1.698274e-22, 
    1.69635e-22, 1.704906e-22, 1.707478e-22, 1.719767e-22, 1.714604e-22, 
    1.722853e-22, 1.715418e-22, 1.716731e-22, 1.723108e-22, 1.715821e-22, 
    1.731829e-22, 1.720951e-22, 1.741203e-22, 1.730283e-22, 1.741888e-22, 
    1.739782e-22, 1.743274e-22, 1.7464e-22, 1.743659e-22, 1.750882e-22, 
    1.749207e-22, 1.755274e-22, 1.701006e-22, 1.704493e-22, 1.704192e-22, 
    1.707851e-22, 1.71056e-22, 1.716508e-22, 1.726425e-22, 1.722693e-22, 
    1.729557e-22, 1.730934e-22, 1.720513e-22, 1.7269e-22, 1.706834e-22, 
    1.709973e-22, 1.708109e-22, 1.701277e-22, 1.723543e-22, 1.711903e-22, 
    1.733582e-22, 1.727159e-22, 1.745953e-22, 1.736581e-22, 1.748285e-22, 
    1.75613e-22, 1.763574e-22, 1.772268e-22, 1.706405e-22, 1.704033e-22, 
    1.708289e-22, 1.714178e-22, 1.719886e-22, 1.727549e-22, 1.728338e-22, 
    1.729775e-22, 1.733509e-22, 1.73665e-22, 1.730223e-22, 1.737438e-22, 
    1.710687e-22, 1.724573e-22, 1.70313e-22, 1.70943e-22, 1.713833e-22, 
    1.711908e-22, 1.722269e-22, 1.724752e-22, 1.734866e-22, 1.729636e-22, 
    1.754185e-22, 1.747051e-22, 1.778933e-22, 1.768087e-22, 1.703203e-22, 
    1.7064e-22, 1.717666e-22, 1.712242e-22, 1.728065e-22, 1.732007e-22, 
    1.735223e-22, 1.739329e-22, 1.739778e-22, 1.742215e-22, 1.738222e-22, 
    1.74206e-22, 1.727565e-22, 1.734033e-22, 1.716336e-22, 1.720627e-22, 
    1.718654e-22, 1.716487e-22, 1.723181e-22, 1.730322e-22, 1.730486e-22, 
    1.732778e-22, 1.73923e-22, 1.72813e-22, 1.755953e-22, 1.741289e-22, 
    1.709892e-22, 1.716099e-22, 1.717036e-22, 1.71456e-22, 1.731612e-22, 
    1.725406e-22, 1.742157e-22, 1.737621e-22, 1.745061e-22, 1.74136e-22, 
    1.740815e-22, 1.736074e-22, 1.733124e-22, 1.725688e-22, 1.719659e-22, 
    1.71491e-22, 1.716002e-22, 1.721239e-22, 1.730762e-22, 1.739813e-22, 
    1.737826e-22, 1.744495e-22, 1.726903e-22, 1.734258e-22, 1.731409e-22, 
    1.738847e-22, 1.722592e-22, 1.736393e-22, 1.719073e-22, 1.720589e-22, 
    1.725283e-22, 1.734751e-22, 1.736867e-22, 1.739108e-22, 1.737727e-22, 
    1.731006e-22, 1.729912e-22, 1.725172e-22, 1.723859e-22, 1.72026e-22, 
    1.717278e-22, 1.719999e-22, 1.722858e-22, 1.731014e-22, 1.738381e-22, 
    1.746443e-22, 1.748425e-22, 1.751105e-22, 1.743478e-22, 1.75607e-22, 
    1.745335e-22, 1.76397e-22, 1.737212e-22, 1.745041e-22, 1.725501e-22, 
    1.728317e-22, 1.733406e-22, 1.745145e-22, 1.738813e-22, 1.746225e-22, 
    1.72987e-22, 1.721415e-22, 1.719246e-22, 1.715188e-22, 1.719339e-22, 
    1.719001e-22, 1.722984e-22, 1.721704e-22, 1.731285e-22, 1.726134e-22, 
    1.740799e-22, 1.746169e-22, 1.754633e-22, 1.763954e-22, 1.7735e-22, 
    1.777721e-22, 1.779009e-22, 1.779546e-22,
  2.342864e-27, 2.35708e-27, 2.354314e-27, 2.365813e-27, 2.359434e-27, 
    2.366968e-27, 2.345747e-27, 2.357639e-27, 2.350046e-27, 2.34415e-27, 
    2.388243e-27, 2.366329e-27, 2.412009e-27, 2.397227e-27, 2.434519e-27, 
    2.409695e-27, 2.439552e-27, 2.433816e-27, 2.451153e-27, 2.446177e-27, 
    2.459573e-27, 2.453452e-27, 2.471121e-27, 2.456023e-27, 2.458373e-27, 
    2.452957e-27, 2.37074e-27, 2.385501e-27, 2.369864e-27, 2.371965e-27, 
    2.371025e-27, 2.35956e-27, 2.35379e-27, 2.341791e-27, 2.343968e-27, 
    2.352789e-27, 2.37291e-27, 2.366074e-27, 2.383364e-27, 2.382973e-27, 
    2.402672e-27, 2.393587e-27, 2.427802e-27, 2.418021e-27, 2.446385e-27, 
    2.439224e-27, 2.446045e-27, 2.443977e-27, 2.446072e-27, 2.435578e-27, 
    2.440069e-27, 2.430856e-27, 2.395228e-27, 2.405649e-27, 2.375577e-27, 
    2.357905e-27, 2.346265e-27, 2.338026e-27, 2.339187e-27, 2.341403e-27, 
    2.352841e-27, 2.36365e-27, 2.371911e-27, 2.377448e-27, 2.382916e-27, 
    2.3997e-27, 2.408961e-27, 2.429776e-27, 2.426022e-27, 2.432394e-27, 
    2.438513e-27, 2.448796e-27, 2.447104e-27, 2.451639e-27, 2.432235e-27, 
    2.445113e-27, 2.423883e-27, 2.429673e-27, 2.384353e-27, 2.367919e-27, 
    2.360918e-27, 2.354843e-27, 2.340081e-27, 2.350265e-27, 2.346244e-27, 
    2.355829e-27, 2.361929e-27, 2.358912e-27, 2.377599e-27, 2.370318e-27, 
    2.409511e-27, 2.392198e-27, 2.437799e-27, 2.426793e-27, 2.440445e-27, 
    2.433474e-27, 2.445424e-27, 2.434667e-27, 2.453334e-27, 2.448638e-27, 
    2.454622e-27, 2.45652e-27, 2.43407e-27, 2.44604e-27, 2.358825e-27, 
    2.359317e-27, 2.361613e-27, 2.351531e-27, 2.350919e-27, 2.341729e-27, 
    2.349909e-27, 2.353396e-27, 2.362287e-27, 2.367549e-27, 2.372565e-27, 
    2.383624e-27, 2.39606e-27, 2.414314e-27, 2.427505e-27, 2.436377e-27, 
    2.430937e-27, 2.435739e-27, 2.430369e-27, 2.427858e-27, 2.447123e-27, 
    2.440108e-27, 2.454985e-27, 2.453681e-27, 2.451745e-27, 2.453828e-27, 
    2.359663e-27, 2.356834e-27, 2.347019e-27, 2.354697e-27, 2.340731e-27, 
    2.348533e-27, 2.353026e-27, 2.370458e-27, 2.374315e-27, 2.37788e-27, 
    2.384946e-27, 2.394034e-27, 2.410744e-27, 2.425412e-27, 2.438872e-27, 
    2.437885e-27, 2.438232e-27, 2.441241e-27, 2.433785e-27, 2.442467e-27, 
    2.443921e-27, 2.440112e-27, 2.453506e-27, 2.447202e-27, 2.453653e-27, 
    2.449545e-27, 2.357754e-27, 2.36252e-27, 2.359943e-27, 2.364788e-27, 
    2.36137e-27, 2.376585e-27, 2.381163e-27, 2.403053e-27, 2.393852e-27, 
    2.408558e-27, 2.395294e-27, 2.397637e-27, 2.409019e-27, 2.396013e-27, 
    2.424591e-27, 2.405166e-27, 2.441358e-27, 2.421831e-27, 2.442584e-27, 
    2.438813e-27, 2.445065e-27, 2.450668e-27, 2.448969e-27, 2.461953e-27, 
    2.458941e-27, 2.469851e-27, 2.369643e-27, 2.375847e-27, 2.37531e-27, 
    2.381823e-27, 2.386646e-27, 2.397238e-27, 2.414933e-27, 2.40827e-27, 
    2.420525e-27, 2.422988e-27, 2.404379e-27, 2.415782e-27, 2.380014e-27, 
    2.385604e-27, 2.382282e-27, 2.370127e-27, 2.40979e-27, 2.389042e-27, 
    2.427721e-27, 2.416243e-27, 2.449867e-27, 2.433088e-27, 2.457283e-27, 
    2.471397e-27, 2.484877e-27, 2.500961e-27, 2.379249e-27, 2.375026e-27, 
    2.382601e-27, 2.393096e-27, 2.403261e-27, 2.41694e-27, 2.418348e-27, 
    2.420916e-27, 2.42759e-27, 2.433207e-27, 2.421719e-27, 2.434618e-27, 
    2.386883e-27, 2.411628e-27, 2.373422e-27, 2.384639e-27, 2.392481e-27, 
    2.389048e-27, 2.407511e-27, 2.411944e-27, 2.430019e-27, 2.420667e-27, 
    2.467899e-27, 2.451839e-27, 2.513298e-27, 2.493224e-27, 2.37355e-27, 
    2.379239e-27, 2.399303e-27, 2.389642e-27, 2.41786e-27, 2.424907e-27, 
    2.430655e-27, 2.438004e-27, 2.438806e-27, 2.44317e-27, 2.43602e-27, 
    2.442892e-27, 2.416969e-27, 2.428527e-27, 2.396929e-27, 2.404584e-27, 
    2.401063e-27, 2.397199e-27, 2.40914e-27, 2.421897e-27, 2.422186e-27, 
    2.426286e-27, 2.437841e-27, 2.417977e-27, 2.471088e-27, 2.441524e-27, 
    2.385455e-27, 2.396512e-27, 2.398179e-27, 2.393772e-27, 2.424199e-27, 
    2.413113e-27, 2.443066e-27, 2.434945e-27, 2.448267e-27, 2.441638e-27, 
    2.440664e-27, 2.432178e-27, 2.426902e-27, 2.413618e-27, 2.402857e-27, 
    2.394394e-27, 2.396334e-27, 2.405677e-27, 2.422683e-27, 2.438871e-27, 
    2.435315e-27, 2.447253e-27, 2.415786e-27, 2.428933e-27, 2.423839e-27, 
    2.437141e-27, 2.408089e-27, 2.432762e-27, 2.40181e-27, 2.404514e-27, 
    2.412894e-27, 2.429816e-27, 2.433596e-27, 2.437609e-27, 2.435135e-27, 
    2.423119e-27, 2.421162e-27, 2.412694e-27, 2.410352e-27, 2.403926e-27, 
    2.398609e-27, 2.403463e-27, 2.408565e-27, 2.42313e-27, 2.436308e-27, 
    2.450746e-27, 2.454296e-27, 2.462361e-27, 2.448649e-27, 2.471299e-27, 
    2.451996e-27, 2.485622e-27, 2.434222e-27, 2.45146e-27, 2.413281e-27, 
    2.41831e-27, 2.427411e-27, 2.448423e-27, 2.437078e-27, 2.450358e-27, 
    2.421086e-27, 2.405991e-27, 2.402118e-27, 2.394888e-27, 2.402284e-27, 
    2.401681e-27, 2.408788e-27, 2.406503e-27, 2.423615e-27, 2.414412e-27, 
    2.440635e-27, 2.450256e-27, 2.4687e-27, 2.485585e-27, 2.503234e-27, 
    2.511051e-27, 2.513435e-27, 2.514432e-27,
  1.04139e-32, 1.049388e-32, 1.04783e-32, 1.05431e-32, 1.050713e-32, 
    1.054961e-32, 1.04301e-32, 1.049704e-32, 1.045428e-32, 1.042112e-32, 
    1.067099e-32, 1.0546e-32, 1.080725e-32, 1.072278e-32, 1.09362e-32, 
    1.079403e-32, 1.096508e-32, 1.093214e-32, 1.103172e-32, 1.100311e-32, 
    1.109436e-32, 1.104494e-32, 1.116104e-32, 1.107386e-32, 1.108743e-32, 
    1.104209e-32, 1.057087e-32, 1.065512e-32, 1.056594e-32, 1.057779e-32, 
    1.057249e-32, 1.050785e-32, 1.047538e-32, 1.040785e-32, 1.042009e-32, 
    1.046973e-32, 1.058313e-32, 1.054455e-32, 1.064269e-32, 1.064042e-32, 
    1.075387e-32, 1.070188e-32, 1.089765e-32, 1.084162e-32, 1.100431e-32, 
    1.096318e-32, 1.100236e-32, 1.099047e-32, 1.100251e-32, 1.094226e-32, 
    1.096803e-32, 1.091516e-32, 1.071136e-32, 1.077088e-32, 1.059818e-32, 
    1.049855e-32, 1.043301e-32, 1.03867e-32, 1.039322e-32, 1.040568e-32, 
    1.047002e-32, 1.053089e-32, 1.057748e-32, 1.060873e-32, 1.06401e-32, 
    1.073693e-32, 1.078982e-32, 1.090898e-32, 1.088745e-32, 1.0924e-32, 
    1.09591e-32, 1.101818e-32, 1.100844e-32, 1.103452e-32, 1.092307e-32, 
    1.099701e-32, 1.087519e-32, 1.090838e-32, 1.064848e-32, 1.055496e-32, 
    1.051553e-32, 1.048129e-32, 1.039825e-32, 1.045552e-32, 1.04329e-32, 
    1.048683e-32, 1.052119e-32, 1.050419e-32, 1.060959e-32, 1.056849e-32, 
    1.079296e-32, 1.069384e-32, 1.0955e-32, 1.089187e-32, 1.097019e-32, 
    1.093017e-32, 1.099879e-32, 1.093702e-32, 1.104427e-32, 1.103126e-32, 
    1.105168e-32, 1.107671e-32, 1.09336e-32, 1.100234e-32, 1.05037e-32, 
    1.050647e-32, 1.051941e-32, 1.046265e-32, 1.04592e-32, 1.040751e-32, 
    1.045351e-32, 1.047314e-32, 1.05232e-32, 1.055288e-32, 1.058117e-32, 
    1.06442e-32, 1.071613e-32, 1.082042e-32, 1.089595e-32, 1.094683e-32, 
    1.091562e-32, 1.094317e-32, 1.091237e-32, 1.089797e-32, 1.102253e-32, 
    1.096826e-32, 1.106786e-32, 1.106033e-32, 1.103514e-32, 1.106118e-32, 
    1.050842e-32, 1.049248e-32, 1.043725e-32, 1.048045e-32, 1.04019e-32, 
    1.044577e-32, 1.047106e-32, 1.05693e-32, 1.059105e-32, 1.061118e-32, 
    1.065184e-32, 1.070446e-32, 1.08e-32, 1.088396e-32, 1.096115e-32, 
    1.095548e-32, 1.095748e-32, 1.097476e-32, 1.093196e-32, 1.09818e-32, 
    1.099016e-32, 1.096828e-32, 1.105932e-32, 1.102297e-32, 1.106017e-32, 
    1.103648e-32, 1.049767e-32, 1.052452e-32, 1.051e-32, 1.053731e-32, 
    1.051804e-32, 1.060388e-32, 1.062998e-32, 1.075606e-32, 1.070341e-32, 
    1.078751e-32, 1.071174e-32, 1.072512e-32, 1.079017e-32, 1.071584e-32, 
    1.087927e-32, 1.076814e-32, 1.097543e-32, 1.086348e-32, 1.098247e-32, 
    1.096082e-32, 1.099672e-32, 1.102894e-32, 1.103316e-32, 1.110808e-32, 
    1.109069e-32, 1.115369e-32, 1.056469e-32, 1.059971e-32, 1.059666e-32, 
    1.063377e-32, 1.066169e-32, 1.072283e-32, 1.082396e-32, 1.078584e-32, 
    1.085596e-32, 1.087007e-32, 1.076361e-32, 1.082882e-32, 1.062333e-32, 
    1.065568e-32, 1.063644e-32, 1.056742e-32, 1.079456e-32, 1.067557e-32, 
    1.089719e-32, 1.083145e-32, 1.102433e-32, 1.092798e-32, 1.108112e-32, 
    1.116266e-32, 1.124072e-32, 1.133456e-32, 1.061891e-32, 1.059506e-32, 
    1.063827e-32, 1.069905e-32, 1.075723e-32, 1.083544e-32, 1.08435e-32, 
    1.08582e-32, 1.089643e-32, 1.092865e-32, 1.086281e-32, 1.093674e-32, 
    1.066311e-32, 1.080506e-32, 1.058602e-32, 1.065009e-32, 1.069547e-32, 
    1.067559e-32, 1.07815e-32, 1.080685e-32, 1.091037e-32, 1.085677e-32, 
    1.114244e-32, 1.103569e-32, 1.140756e-32, 1.12894e-32, 1.058673e-32, 
    1.061885e-32, 1.073463e-32, 1.067903e-32, 1.08407e-32, 1.088106e-32, 
    1.091401e-32, 1.095618e-32, 1.096077e-32, 1.098584e-32, 1.094478e-32, 
    1.098424e-32, 1.083561e-32, 1.090181e-32, 1.072106e-32, 1.076478e-32, 
    1.074467e-32, 1.072261e-32, 1.079081e-32, 1.086384e-32, 1.086547e-32, 
    1.088897e-32, 1.095532e-32, 1.084137e-32, 1.116091e-32, 1.097646e-32, 
    1.065479e-32, 1.071871e-32, 1.072821e-32, 1.070294e-32, 1.087701e-32, 
    1.081355e-32, 1.098524e-32, 1.093861e-32, 1.101513e-32, 1.097704e-32, 
    1.097144e-32, 1.092274e-32, 1.08925e-32, 1.081644e-32, 1.075492e-32, 
    1.070654e-32, 1.071767e-32, 1.077103e-32, 1.086833e-32, 1.096116e-32, 
    1.094075e-32, 1.10093e-32, 1.082883e-32, 1.090414e-32, 1.087496e-32, 
    1.095122e-32, 1.078482e-32, 1.092616e-32, 1.074893e-32, 1.076438e-32, 
    1.081229e-32, 1.090922e-32, 1.093087e-32, 1.095391e-32, 1.093971e-32, 
    1.087083e-32, 1.085961e-32, 1.081114e-32, 1.079776e-32, 1.076102e-32, 
    1.073065e-32, 1.075837e-32, 1.078754e-32, 1.087089e-32, 1.094645e-32, 
    1.102939e-32, 1.10498e-32, 1.111047e-32, 1.103135e-32, 1.116214e-32, 
    1.10507e-32, 1.124513e-32, 1.093451e-32, 1.104757e-32, 1.08145e-32, 
    1.084328e-32, 1.089543e-32, 1.101605e-32, 1.095086e-32, 1.102717e-32, 
    1.085918e-32, 1.077284e-32, 1.075069e-32, 1.070939e-32, 1.075164e-32, 
    1.074819e-32, 1.07888e-32, 1.077574e-32, 1.087366e-32, 1.082097e-32, 
    1.097128e-32, 1.102658e-32, 1.114705e-32, 1.124487e-32, 1.134781e-32, 
    1.139412e-32, 1.140837e-32, 1.141432e-32,
  1.510159e-38, 1.525776e-38, 1.522729e-38, 1.535419e-38, 1.528368e-38, 
    1.536696e-38, 1.513316e-38, 1.526396e-38, 1.518034e-38, 1.511564e-38, 
    1.560644e-38, 1.535988e-38, 1.587507e-38, 1.570888e-38, 1.613511e-38, 
    1.584903e-38, 1.619381e-38, 1.612682e-38, 1.632962e-38, 1.627123e-38, 
    1.648366e-38, 1.635664e-38, 1.662107e-38, 1.644146e-38, 1.646937e-38, 
    1.635083e-38, 1.540869e-38, 1.557497e-38, 1.539899e-38, 1.54223e-38, 
    1.541186e-38, 1.528511e-38, 1.52216e-38, 1.508979e-38, 1.511365e-38, 
    1.521053e-38, 1.543279e-38, 1.535701e-38, 1.555021e-38, 1.554573e-38, 
    1.576994e-38, 1.566764e-38, 1.605686e-38, 1.594347e-38, 1.627367e-38, 
    1.61899e-38, 1.626971e-38, 1.624547e-38, 1.627002e-38, 1.614737e-38, 
    1.619979e-38, 1.609236e-38, 1.568647e-38, 1.580341e-38, 1.546238e-38, 
    1.526695e-38, 1.513885e-38, 1.504861e-38, 1.506131e-38, 1.508558e-38, 
    1.52111e-38, 1.533022e-38, 1.542165e-38, 1.548312e-38, 1.554508e-38, 
    1.573674e-38, 1.584073e-38, 1.607985e-38, 1.603617e-38, 1.611031e-38, 
    1.61816e-38, 1.630198e-38, 1.628211e-38, 1.633537e-38, 1.61084e-38, 
    1.625882e-38, 1.601133e-38, 1.607859e-38, 1.556183e-38, 1.537743e-38, 
    1.530018e-38, 1.523313e-38, 1.50711e-38, 1.518277e-38, 1.513864e-38, 
    1.524394e-38, 1.531121e-38, 1.527791e-38, 1.54848e-38, 1.5404e-38, 
    1.584692e-38, 1.565169e-38, 1.617327e-38, 1.604513e-38, 1.620416e-38, 
    1.612281e-38, 1.626245e-38, 1.613671e-38, 1.635527e-38, 1.635402e-38, 
    1.637044e-38, 1.644731e-38, 1.612977e-38, 1.626968e-38, 1.527696e-38, 
    1.528239e-38, 1.530772e-38, 1.51967e-38, 1.518996e-38, 1.508912e-38, 
    1.517884e-38, 1.521719e-38, 1.531514e-38, 1.537335e-38, 1.542892e-38, 
    1.555322e-38, 1.569584e-38, 1.590103e-38, 1.60534e-38, 1.615665e-38, 
    1.609327e-38, 1.614921e-38, 1.608668e-38, 1.605748e-38, 1.633611e-38, 
    1.620026e-38, 1.642912e-38, 1.641365e-38, 1.633663e-38, 1.64154e-38, 
    1.52862e-38, 1.5255e-38, 1.514711e-38, 1.523148e-38, 1.507819e-38, 
    1.516375e-38, 1.521316e-38, 1.540562e-38, 1.544833e-38, 1.548795e-38, 
    1.556836e-38, 1.567278e-38, 1.586076e-38, 1.602913e-38, 1.618577e-38, 
    1.617424e-38, 1.61783e-38, 1.621347e-38, 1.612645e-38, 1.622781e-38, 
    1.624486e-38, 1.620027e-38, 1.641158e-38, 1.633699e-38, 1.641332e-38, 
    1.63647e-38, 1.526514e-38, 1.531773e-38, 1.528929e-38, 1.534281e-38, 
    1.530506e-38, 1.547361e-38, 1.552511e-38, 1.577429e-38, 1.56707e-38, 
    1.583615e-38, 1.568721e-38, 1.571347e-38, 1.584146e-38, 1.569524e-38, 
    1.601967e-38, 1.579807e-38, 1.621484e-38, 1.598774e-38, 1.622918e-38, 
    1.618509e-38, 1.62582e-38, 1.632396e-38, 1.63579e-38, 1.651186e-38, 
    1.647606e-38, 1.660587e-38, 1.539653e-38, 1.546538e-38, 1.545937e-38, 
    1.553257e-38, 1.558788e-38, 1.570896e-38, 1.590799e-38, 1.583285e-38, 
    1.597244e-38, 1.600099e-38, 1.578908e-38, 1.591765e-38, 1.551191e-38, 
    1.5576e-38, 1.553785e-38, 1.540191e-38, 1.585005e-38, 1.561545e-38, 
    1.605593e-38, 1.592294e-38, 1.631455e-38, 1.611841e-38, 1.645638e-38, 
    1.662445e-38, 1.678557e-38, 1.698062e-38, 1.550317e-38, 1.545621e-38, 
    1.554147e-38, 1.566205e-38, 1.577656e-38, 1.5931e-38, 1.594726e-38, 
    1.597699e-38, 1.605436e-38, 1.611971e-38, 1.598635e-38, 1.613615e-38, 
    1.559079e-38, 1.587073e-38, 1.543845e-38, 1.556494e-38, 1.565494e-38, 
    1.561545e-38, 1.58243e-38, 1.587423e-38, 1.608266e-38, 1.597409e-38, 
    1.658273e-38, 1.63378e-38, 1.713529e-38, 1.68857e-38, 1.543983e-38, 
    1.550304e-38, 1.573217e-38, 1.562227e-38, 1.594162e-38, 1.602325e-38, 
    1.609e-38, 1.617568e-38, 1.618501e-38, 1.623605e-38, 1.615249e-38, 
    1.623277e-38, 1.593134e-38, 1.606527e-38, 1.57055e-38, 1.579141e-38, 
    1.575184e-38, 1.570852e-38, 1.584263e-38, 1.598842e-38, 1.599168e-38, 
    1.603928e-38, 1.617407e-38, 1.594296e-38, 1.662095e-38, 1.621706e-38, 
    1.557419e-38, 1.570094e-38, 1.571953e-38, 1.566974e-38, 1.601504e-38, 
    1.588745e-38, 1.623482e-38, 1.613996e-38, 1.629574e-38, 1.621811e-38, 
    1.620672e-38, 1.610772e-38, 1.60464e-38, 1.589315e-38, 1.577202e-38, 
    1.567688e-38, 1.569883e-38, 1.580371e-38, 1.599751e-38, 1.618581e-38, 
    1.614434e-38, 1.628385e-38, 1.591765e-38, 1.607002e-38, 1.601091e-38, 
    1.616558e-38, 1.583083e-38, 1.611481e-38, 1.576022e-38, 1.57906e-38, 
    1.588497e-38, 1.608035e-38, 1.612424e-38, 1.617107e-38, 1.614217e-38, 
    1.600255e-38, 1.597984e-38, 1.588269e-38, 1.585633e-38, 1.578398e-38, 
    1.572431e-38, 1.57788e-38, 1.583622e-38, 1.600265e-38, 1.615589e-38, 
    1.632488e-38, 1.636657e-38, 1.651685e-38, 1.635425e-38, 1.662349e-38, 
    1.639405e-38, 1.679474e-38, 1.61317e-38, 1.638754e-38, 1.588931e-38, 
    1.594681e-38, 1.605239e-38, 1.62977e-38, 1.616485e-38, 1.632038e-38, 
    1.597896e-38, 1.580729e-38, 1.576369e-38, 1.568255e-38, 1.576555e-38, 
    1.575878e-38, 1.583867e-38, 1.581295e-38, 1.600827e-38, 1.590208e-38, 
    1.620641e-38, 1.631917e-38, 1.659218e-38, 1.679413e-38, 1.700853e-38, 
    1.710672e-38, 1.713699e-38, 1.714966e-38,
  8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 9.809089e-45, 9.809089e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 9.809089e-45, 9.809089e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 9.809089e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 9.809089e-45, 9.809089e-45, 
    9.809089e-45, 9.809089e-45, 9.809089e-45,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  2.055945e-05, 2.036958e-05, 2.040654e-05, 2.025308e-05, 2.033826e-05, 
    2.02377e-05, 2.052101e-05, 2.036203e-05, 2.046357e-05, 2.054239e-05, 
    1.995421e-05, 2.024622e-05, 1.964962e-05, 1.983683e-05, 1.936562e-05, 
    1.967878e-05, 1.930231e-05, 1.937469e-05, 1.915667e-05, 1.92192e-05, 
    1.894019e-05, 1.912779e-05, 1.879484e-05, 1.898519e-05, 1.895544e-05, 
    1.913399e-05, 2.018758e-05, 1.999063e-05, 2.019922e-05, 2.017118e-05, 
    2.018377e-05, 2.033649e-05, 2.041331e-05, 2.057395e-05, 2.054482e-05, 
    2.042682e-05, 2.015857e-05, 2.024976e-05, 2.001972e-05, 2.002493e-05, 
    1.97679e-05, 1.988391e-05, 1.945048e-05, 1.957395e-05, 1.921659e-05, 
    1.930663e-05, 1.922082e-05, 1.924685e-05, 1.922048e-05, 1.935248e-05, 
    1.929595e-05, 1.941201e-05, 1.98622e-05, 1.973019e-05, 2.012313e-05, 
    2.035827e-05, 2.051404e-05, 2.062433e-05, 2.060875e-05, 2.057903e-05, 
    2.042613e-05, 2.028206e-05, 2.017205e-05, 2.009836e-05, 2.002568e-05, 
    1.980513e-05, 1.968815e-05, 1.942548e-05, 1.947297e-05, 1.939251e-05, 
    1.931558e-05, 1.918621e-05, 1.920752e-05, 1.915046e-05, 1.939465e-05, 
    1.923245e-05, 1.950001e-05, 1.942693e-05, 2.000584e-05, 2.022518e-05, 
    2.031813e-05, 2.039944e-05, 2.059676e-05, 2.046055e-05, 2.051428e-05, 
    2.03864e-05, 2.0305e-05, 2.034527e-05, 2.009635e-05, 2.019323e-05, 
    1.968121e-05, 1.990223e-05, 1.932456e-05, 1.946323e-05, 1.929128e-05, 
    1.937908e-05, 1.922857e-05, 1.936404e-05, 1.912922e-05, 1.90786e-05, 
    1.9113e-05, 1.897904e-05, 1.937154e-05, 1.922081e-05, 2.03464e-05, 
    2.033983e-05, 2.030924e-05, 2.044362e-05, 2.045183e-05, 2.057474e-05, 
    2.04654e-05, 2.041877e-05, 2.030028e-05, 2.023009e-05, 2.016329e-05, 
    2.00162e-05, 1.985153e-05, 1.962061e-05, 1.945425e-05, 1.934251e-05, 
    1.941105e-05, 1.935054e-05, 1.941818e-05, 1.944986e-05, 1.90978e-05, 
    1.929542e-05, 1.899841e-05, 1.901491e-05, 1.91491e-05, 1.901305e-05, 
    2.033522e-05, 2.0373e-05, 2.050399e-05, 2.04015e-05, 2.058812e-05, 
    2.048372e-05, 2.042361e-05, 2.019119e-05, 2.014004e-05, 2.009254e-05, 
    1.999866e-05, 1.987798e-05, 1.966575e-05, 1.948057e-05, 1.93111e-05, 
    1.932353e-05, 1.931916e-05, 1.928124e-05, 1.937511e-05, 1.926582e-05, 
    1.924745e-05, 1.929545e-05, 1.901712e-05, 1.909693e-05, 1.901526e-05, 
    1.906724e-05, 2.036073e-05, 2.029713e-05, 2.03315e-05, 2.026685e-05, 
    2.03124e-05, 2.010961e-05, 2.004869e-05, 1.97629e-05, 1.988035e-05, 
    1.969336e-05, 1.986139e-05, 1.983164e-05, 1.968722e-05, 1.985232e-05, 
    1.949078e-05, 1.973607e-05, 1.927977e-05, 1.952543e-05, 1.926434e-05, 
    1.931184e-05, 1.92332e-05, 1.916268e-05, 1.907451e-05, 1.891036e-05, 
    1.894841e-05, 1.881094e-05, 2.020222e-05, 2.011952e-05, 2.012681e-05, 
    2.004018e-05, 1.997603e-05, 1.983679e-05, 1.961287e-05, 1.969716e-05, 
    1.954235e-05, 1.951122e-05, 1.97464e-05, 1.960209e-05, 2.006412e-05, 
    1.998967e-05, 2.003402e-05, 2.019569e-05, 1.967773e-05, 1.994404e-05, 
    1.945149e-05, 1.959636e-05, 1.917274e-05, 1.938371e-05, 1.896934e-05, 
    1.879118e-05, 1.862317e-05, 1.842629e-05, 2.007435e-05, 2.013059e-05, 
    2.002987e-05, 1.989024e-05, 1.976046e-05, 1.958753e-05, 1.956982e-05, 
    1.953736e-05, 1.945323e-05, 1.938242e-05, 1.952708e-05, 1.936466e-05, 
    1.997237e-05, 1.965457e-05, 2.015183e-05, 2.000246e-05, 1.989848e-05, 
    1.994413e-05, 1.970679e-05, 1.965073e-05, 1.942245e-05, 1.954056e-05, 
    1.883518e-05, 1.914776e-05, 1.827609e-05, 1.852086e-05, 2.015023e-05, 
    2.007455e-05, 1.981048e-05, 1.993626e-05, 1.957598e-05, 1.9487e-05, 
    1.94146e-05, 1.932192e-05, 1.931191e-05, 1.925694e-05, 1.9347e-05, 
    1.92605e-05, 1.958716e-05, 1.944137e-05, 1.984073e-05, 1.974373e-05, 
    1.978838e-05, 1.983731e-05, 1.968619e-05, 1.95248e-05, 1.952137e-05, 
    1.946954e-05, 1.932324e-05, 1.957451e-05, 1.879462e-05, 1.927699e-05, 
    1.999193e-05, 1.984571e-05, 1.982483e-05, 1.988152e-05, 1.949592e-05, 
    1.963589e-05, 1.925828e-05, 1.936054e-05, 1.919292e-05, 1.927626e-05, 
    1.928851e-05, 1.939539e-05, 1.946185e-05, 1.962947e-05, 1.976556e-05, 
    1.98733e-05, 1.984827e-05, 1.972987e-05, 1.951493e-05, 1.9311e-05, 
    1.935572e-05, 1.920567e-05, 1.960216e-05, 1.943617e-05, 1.950036e-05, 
    1.933285e-05, 1.96994e-05, 1.938732e-05, 1.977893e-05, 1.974469e-05, 
    1.963866e-05, 1.942488e-05, 1.937752e-05, 1.932689e-05, 1.935814e-05, 
    1.950947e-05, 1.953423e-05, 1.964125e-05, 1.967075e-05, 1.975215e-05, 
    1.981946e-05, 1.975796e-05, 1.969331e-05, 1.950941e-05, 1.934326e-05, 
    1.916167e-05, 1.911717e-05, 1.890487e-05, 1.907822e-05, 1.879191e-05, 
    1.903535e-05, 1.861346e-05, 1.936922e-05, 1.904254e-05, 1.963384e-05, 
    1.957031e-05, 1.945524e-05, 1.919066e-05, 1.933364e-05, 1.91664e-05, 
    1.953521e-05, 1.972577e-05, 1.977501e-05, 1.986675e-05, 1.977291e-05, 
    1.978055e-05, 1.969065e-05, 1.971955e-05, 1.95033e-05, 1.961954e-05, 
    1.928881e-05, 1.916773e-05, 1.882535e-05, 1.861428e-05, 1.839885e-05, 
    1.830354e-05, 1.827451e-05, 1.826237e-05,
  1.427401e-05, 1.408346e-05, 1.412053e-05, 1.396666e-05, 1.405205e-05, 
    1.395125e-05, 1.423542e-05, 1.407588e-05, 1.417776e-05, 1.425689e-05, 
    1.366751e-05, 1.39598e-05, 1.336343e-05, 1.355026e-05, 1.308059e-05, 
    1.33925e-05, 1.301764e-05, 1.308963e-05, 1.287298e-05, 1.293507e-05, 
    1.265765e-05, 1.284431e-05, 1.251379e-05, 1.270226e-05, 1.267277e-05, 
    1.285046e-05, 1.390105e-05, 1.370392e-05, 1.391272e-05, 1.388463e-05, 
    1.389724e-05, 1.405028e-05, 1.412731e-05, 1.428859e-05, 1.425933e-05, 
    1.414088e-05, 1.3872e-05, 1.396335e-05, 1.373306e-05, 1.373826e-05, 
    1.348144e-05, 1.359729e-05, 1.316504e-05, 1.328801e-05, 1.293248e-05, 
    1.302194e-05, 1.293667e-05, 1.296254e-05, 1.293634e-05, 1.306754e-05, 
    1.301133e-05, 1.312676e-05, 1.357559e-05, 1.34438e-05, 1.383652e-05, 
    1.40721e-05, 1.422842e-05, 1.43392e-05, 1.432354e-05, 1.429369e-05, 
    1.414019e-05, 1.399572e-05, 1.388551e-05, 1.381174e-05, 1.373901e-05, 
    1.351858e-05, 1.340185e-05, 1.314015e-05, 1.318743e-05, 1.310735e-05, 
    1.303084e-05, 1.29023e-05, 1.292347e-05, 1.286681e-05, 1.310948e-05, 
    1.294822e-05, 1.321436e-05, 1.31416e-05, 1.371913e-05, 1.393872e-05, 
    1.403186e-05, 1.411341e-05, 1.43115e-05, 1.417473e-05, 1.422866e-05, 
    1.410034e-05, 1.401871e-05, 1.405909e-05, 1.380972e-05, 1.390672e-05, 
    1.339493e-05, 1.361559e-05, 1.303977e-05, 1.317773e-05, 1.300669e-05, 
    1.309399e-05, 1.294437e-05, 1.307903e-05, 1.284573e-05, 1.279488e-05, 
    1.282963e-05, 1.269616e-05, 1.308649e-05, 1.293667e-05, 1.406022e-05, 
    1.405363e-05, 1.402296e-05, 1.415773e-05, 1.416598e-05, 1.428938e-05, 
    1.417959e-05, 1.41328e-05, 1.401399e-05, 1.394364e-05, 1.387673e-05, 
    1.372953e-05, 1.356493e-05, 1.333451e-05, 1.316879e-05, 1.305762e-05, 
    1.31258e-05, 1.306561e-05, 1.313289e-05, 1.316443e-05, 1.281393e-05, 
    1.30108e-05, 1.271537e-05, 1.273173e-05, 1.286546e-05, 1.272988e-05, 
    1.404901e-05, 1.40869e-05, 1.421833e-05, 1.411549e-05, 1.430282e-05, 
    1.419798e-05, 1.413765e-05, 1.390467e-05, 1.385345e-05, 1.380591e-05, 
    1.371199e-05, 1.359136e-05, 1.337951e-05, 1.319499e-05, 1.30264e-05, 
    1.303876e-05, 1.30344e-05, 1.299671e-05, 1.309005e-05, 1.298139e-05, 
    1.296313e-05, 1.301084e-05, 1.273392e-05, 1.281306e-05, 1.273207e-05, 
    1.278361e-05, 1.407459e-05, 1.401082e-05, 1.404528e-05, 1.398047e-05, 
    1.402613e-05, 1.382298e-05, 1.376201e-05, 1.347644e-05, 1.359373e-05, 
    1.340705e-05, 1.357479e-05, 1.354507e-05, 1.340091e-05, 1.356573e-05, 
    1.320515e-05, 1.344966e-05, 1.299525e-05, 1.323965e-05, 1.297992e-05, 
    1.302713e-05, 1.294897e-05, 1.287894e-05, 1.279082e-05, 1.262813e-05, 
    1.266581e-05, 1.252971e-05, 1.391572e-05, 1.38329e-05, 1.384022e-05, 
    1.375351e-05, 1.368935e-05, 1.355022e-05, 1.33268e-05, 1.341086e-05, 
    1.325653e-05, 1.322552e-05, 1.345998e-05, 1.331605e-05, 1.377747e-05, 
    1.370299e-05, 1.374735e-05, 1.390918e-05, 1.339146e-05, 1.365737e-05, 
    1.316605e-05, 1.331034e-05, 1.288893e-05, 1.30986e-05, 1.268655e-05, 
    1.251015e-05, 1.234413e-05, 1.21499e-05, 1.378771e-05, 1.3844e-05, 
    1.374321e-05, 1.36036e-05, 1.347401e-05, 1.330154e-05, 1.328389e-05, 
    1.325156e-05, 1.316779e-05, 1.309732e-05, 1.324131e-05, 1.307965e-05, 
    1.368567e-05, 1.336837e-05, 1.386526e-05, 1.371578e-05, 1.361184e-05, 
    1.365747e-05, 1.342047e-05, 1.336455e-05, 1.313714e-05, 1.325474e-05, 
    1.255368e-05, 1.286412e-05, 1.200203e-05, 1.224314e-05, 1.386366e-05, 
    1.378791e-05, 1.352394e-05, 1.36496e-05, 1.329003e-05, 1.32014e-05, 
    1.312933e-05, 1.303714e-05, 1.30272e-05, 1.297256e-05, 1.306209e-05, 
    1.29761e-05, 1.330117e-05, 1.315598e-05, 1.355416e-05, 1.345732e-05, 
    1.350188e-05, 1.355074e-05, 1.339991e-05, 1.323904e-05, 1.323563e-05, 
    1.318401e-05, 1.303842e-05, 1.328857e-05, 1.251353e-05, 1.299245e-05, 
    1.370526e-05, 1.355912e-05, 1.353827e-05, 1.35949e-05, 1.321029e-05, 
    1.334974e-05, 1.297389e-05, 1.307555e-05, 1.290897e-05, 1.299176e-05, 
    1.300394e-05, 1.311022e-05, 1.317636e-05, 1.334334e-05, 1.34791e-05, 
    1.358669e-05, 1.356168e-05, 1.344348e-05, 1.32292e-05, 1.302629e-05, 
    1.307075e-05, 1.292164e-05, 1.331613e-05, 1.315079e-05, 1.32147e-05, 
    1.304802e-05, 1.341308e-05, 1.310216e-05, 1.349246e-05, 1.345828e-05, 
    1.335251e-05, 1.313955e-05, 1.309245e-05, 1.304209e-05, 1.307317e-05, 
    1.322376e-05, 1.324844e-05, 1.335509e-05, 1.338451e-05, 1.346572e-05, 
    1.353291e-05, 1.347152e-05, 1.340701e-05, 1.322371e-05, 1.305836e-05, 
    1.287794e-05, 1.283378e-05, 1.262267e-05, 1.279448e-05, 1.251085e-05, 
    1.275194e-05, 1.233451e-05, 1.308417e-05, 1.27591e-05, 1.334771e-05, 
    1.328439e-05, 1.316977e-05, 1.290671e-05, 1.30488e-05, 1.288263e-05, 
    1.324941e-05, 1.343938e-05, 1.348854e-05, 1.358015e-05, 1.348644e-05, 
    1.349407e-05, 1.340436e-05, 1.343319e-05, 1.321763e-05, 1.333345e-05, 
    1.300423e-05, 1.288395e-05, 1.254397e-05, 1.233533e-05, 1.212289e-05, 
    1.202905e-05, 1.200049e-05, 1.198855e-05,
  6.636314e-06, 6.51931e-06, 6.542035e-06, 6.44784e-06, 6.500072e-06, 
    6.438428e-06, 6.612575e-06, 6.514665e-06, 6.577147e-06, 6.625778e-06, 
    6.26566e-06, 6.443645e-06, 6.081769e-06, 6.194593e-06, 5.911926e-06, 
    6.099291e-06, 5.874284e-06, 5.917334e-06, 5.787996e-06, 5.824993e-06, 
    5.660149e-06, 5.770937e-06, 5.575113e-06, 5.686577e-06, 5.669103e-06, 
    5.774596e-06, 6.407778e-06, 6.287767e-06, 6.414896e-06, 6.397758e-06, 
    6.405451e-06, 6.498986e-06, 6.546192e-06, 6.645282e-06, 6.627279e-06, 
    6.554515e-06, 6.390054e-06, 6.445818e-06, 6.305468e-06, 6.308632e-06, 
    6.152977e-06, 6.223075e-06, 5.962515e-06, 6.036367e-06, 5.823448e-06, 
    5.876853e-06, 5.825951e-06, 5.841379e-06, 5.82575e-06, 5.904114e-06, 
    5.870513e-06, 5.939567e-06, 6.209933e-06, 6.130241e-06, 6.368433e-06, 
    6.512354e-06, 6.608273e-06, 6.676453e-06, 6.666808e-06, 6.648423e-06, 
    6.554089e-06, 6.465604e-06, 6.398296e-06, 6.353334e-06, 6.309087e-06, 
    6.17543e-06, 6.104933e-06, 5.947593e-06, 5.975946e-06, 5.927941e-06, 
    5.882172e-06, 5.805464e-06, 5.818078e-06, 5.784328e-06, 5.929218e-06, 
    5.83284e-06, 5.992105e-06, 5.948461e-06, 6.297005e-06, 6.430769e-06, 
    6.48771e-06, 6.537663e-06, 6.659392e-06, 6.575289e-06, 6.608422e-06, 
    6.529651e-06, 6.479666e-06, 6.504383e-06, 6.352105e-06, 6.411235e-06, 
    6.100759e-06, 6.234165e-06, 5.887507e-06, 5.970126e-06, 5.867739e-06, 
    5.919946e-06, 5.830543e-06, 5.910993e-06, 5.771782e-06, 5.741549e-06, 
    5.762205e-06, 5.682964e-06, 5.915457e-06, 5.825945e-06, 6.505073e-06, 
    6.50104e-06, 6.482266e-06, 6.564856e-06, 6.569917e-06, 6.645773e-06, 
    6.578276e-06, 6.54956e-06, 6.476776e-06, 6.433774e-06, 6.392943e-06, 
    6.303322e-06, 6.203475e-06, 6.064348e-06, 5.964763e-06, 5.898182e-06, 
    5.938996e-06, 5.902959e-06, 5.943245e-06, 5.962147e-06, 5.75287e-06, 
    5.870197e-06, 5.694347e-06, 5.704052e-06, 5.783523e-06, 5.702958e-06, 
    6.49821e-06, 6.521418e-06, 6.602073e-06, 6.53894e-06, 6.654042e-06, 
    6.589567e-06, 6.552534e-06, 6.409985e-06, 6.378748e-06, 6.349786e-06, 
    6.292667e-06, 6.219483e-06, 6.091463e-06, 5.980481e-06, 5.879514e-06, 
    5.886901e-06, 5.8843e-06, 5.86178e-06, 5.917585e-06, 5.852629e-06, 
    5.841735e-06, 5.870218e-06, 5.705351e-06, 5.752357e-06, 5.704258e-06, 
    5.734855e-06, 6.513874e-06, 6.474841e-06, 6.495928e-06, 6.456282e-06, 
    6.484204e-06, 6.360181e-06, 6.323075e-06, 6.149956e-06, 6.220919e-06, 
    6.108066e-06, 6.209443e-06, 6.191455e-06, 6.104365e-06, 6.203962e-06, 
    5.986578e-06, 6.133781e-06, 5.860905e-06, 6.007299e-06, 5.851753e-06, 
    5.87995e-06, 5.833286e-06, 5.791549e-06, 5.739138e-06, 5.64267e-06, 
    5.664981e-06, 5.584511e-06, 6.416728e-06, 6.366226e-06, 6.370682e-06, 
    6.317905e-06, 6.278917e-06, 6.194573e-06, 6.059706e-06, 6.110363e-06, 
    6.017437e-06, 5.99881e-06, 6.140016e-06, 6.053235e-06, 6.332474e-06, 
    6.287198e-06, 6.314157e-06, 6.412735e-06, 6.098667e-06, 6.259501e-06, 
    5.963118e-06, 6.049802e-06, 5.797495e-06, 5.922702e-06, 5.677268e-06, 
    5.572967e-06, 5.475235e-06, 5.36144e-06, 6.338705e-06, 6.372987e-06, 
    6.311636e-06, 6.2269e-06, 6.14849e-06, 6.044506e-06, 6.033892e-06, 
    6.01445e-06, 5.964162e-06, 5.921936e-06, 6.008294e-06, 5.91136e-06, 
    6.276683e-06, 6.084747e-06, 6.385945e-06, 6.294968e-06, 6.231895e-06, 
    6.259561e-06, 6.11616e-06, 6.082445e-06, 5.945789e-06, 6.016367e-06, 
    5.598662e-06, 5.782725e-06, 5.275196e-06, 5.415997e-06, 6.384969e-06, 
    6.338828e-06, 6.178671e-06, 6.254788e-06, 6.037582e-06, 5.984328e-06, 
    5.941111e-06, 5.885936e-06, 5.879994e-06, 5.847358e-06, 5.900855e-06, 
    5.849474e-06, 6.044285e-06, 5.957079e-06, 6.196956e-06, 6.138407e-06, 
    6.165333e-06, 6.194884e-06, 6.10376e-06, 6.00693e-06, 6.004883e-06, 
    5.973894e-06, 5.886701e-06, 6.036705e-06, 5.574961e-06, 5.859234e-06, 
    6.288577e-06, 6.199958e-06, 6.187341e-06, 6.221628e-06, 5.989662e-06, 
    6.073524e-06, 5.848156e-06, 5.908908e-06, 5.809436e-06, 5.858823e-06, 
    5.866094e-06, 5.929664e-06, 5.969302e-06, 6.06967e-06, 6.151566e-06, 
    6.216655e-06, 6.201511e-06, 6.13005e-06, 6.001021e-06, 5.879447e-06, 
    5.906035e-06, 5.816984e-06, 6.053284e-06, 5.95397e-06, 5.992313e-06, 
    5.892439e-06, 6.111706e-06, 5.924835e-06, 6.159635e-06, 6.138986e-06, 
    6.075191e-06, 5.947233e-06, 5.919021e-06, 5.888893e-06, 5.907484e-06, 
    5.997756e-06, 6.012578e-06, 6.076744e-06, 6.094474e-06, 6.143482e-06, 
    6.1841e-06, 6.146982e-06, 6.108041e-06, 5.997725e-06, 5.898625e-06, 
    5.790952e-06, 5.76467e-06, 5.639441e-06, 5.741314e-06, 5.573383e-06, 
    5.716052e-06, 5.469588e-06, 5.914068e-06, 5.720296e-06, 6.072297e-06, 
    6.034188e-06, 5.965353e-06, 5.808088e-06, 5.892908e-06, 5.793745e-06, 
    6.01316e-06, 6.127577e-06, 6.157268e-06, 6.212691e-06, 6.156002e-06, 
    6.16061e-06, 6.106442e-06, 6.123841e-06, 5.994069e-06, 6.063714e-06, 
    5.866272e-06, 5.794531e-06, 5.592926e-06, 5.470071e-06, 5.345657e-06, 
    5.290927e-06, 5.274296e-06, 5.267346e-06,
  1.674986e-06, 1.63156e-06, 1.639965e-06, 1.605217e-06, 1.624455e-06, 
    1.601758e-06, 1.666145e-06, 1.629844e-06, 1.65298e-06, 1.67106e-06, 
    1.538702e-06, 1.603675e-06, 1.472494e-06, 1.513002e-06, 1.412193e-06, 
    1.478762e-06, 1.39894e-06, 1.414099e-06, 1.368713e-06, 1.381646e-06, 
    1.324328e-06, 1.362763e-06, 1.295069e-06, 1.333463e-06, 1.32742e-06, 
    1.364038e-06, 1.590511e-06, 1.546725e-06, 1.593121e-06, 1.58684e-06, 
    1.589658e-06, 1.624055e-06, 1.641505e-06, 1.678329e-06, 1.671619e-06, 
    1.644587e-06, 1.584019e-06, 1.604473e-06, 1.553156e-06, 1.554307e-06, 
    1.498018e-06, 1.523284e-06, 1.430067e-06, 1.456293e-06, 1.381105e-06, 
    1.399842e-06, 1.381982e-06, 1.387387e-06, 1.381912e-06, 1.409439e-06, 
    1.397614e-06, 1.42195e-06, 1.518536e-06, 1.489853e-06, 1.576112e-06, 
    1.628991e-06, 1.664545e-06, 1.689968e-06, 1.686364e-06, 1.679501e-06, 
    1.64443e-06, 1.611751e-06, 1.587037e-06, 1.570597e-06, 1.554472e-06, 
    1.506097e-06, 1.480782e-06, 1.424788e-06, 1.434826e-06, 1.417843e-06, 
    1.401713e-06, 1.374815e-06, 1.379226e-06, 1.367433e-06, 1.418294e-06, 
    1.384395e-06, 1.440556e-06, 1.425094e-06, 1.550081e-06, 1.598945e-06, 
    1.619896e-06, 1.638347e-06, 1.683595e-06, 1.65229e-06, 1.6646e-06, 
    1.635383e-06, 1.61693e-06, 1.626046e-06, 1.570148e-06, 1.591778e-06, 
    1.479287e-06, 1.527294e-06, 1.40359e-06, 1.432763e-06, 1.396639e-06, 
    1.415021e-06, 1.38359e-06, 1.411863e-06, 1.363057e-06, 1.352533e-06, 
    1.35972e-06, 1.332213e-06, 1.413437e-06, 1.38198e-06, 1.626301e-06, 
    1.624812e-06, 1.617888e-06, 1.64842e-06, 1.650297e-06, 1.678512e-06, 
    1.653398e-06, 1.642751e-06, 1.615865e-06, 1.600048e-06, 1.585077e-06, 
    1.552376e-06, 1.516206e-06, 1.466271e-06, 1.430864e-06, 1.407348e-06, 
    1.421748e-06, 1.409031e-06, 1.42325e-06, 1.429937e-06, 1.356471e-06, 
    1.397503e-06, 1.336153e-06, 1.339515e-06, 1.367152e-06, 1.339136e-06, 
    1.623768e-06, 1.632338e-06, 1.662239e-06, 1.638819e-06, 1.681597e-06, 
    1.657591e-06, 1.643854e-06, 1.59132e-06, 1.579882e-06, 1.569302e-06, 
    1.548502e-06, 1.521986e-06, 1.47596e-06, 1.436433e-06, 1.400778e-06, 
    1.403377e-06, 1.402462e-06, 1.394546e-06, 1.414188e-06, 1.391333e-06, 
    1.387512e-06, 1.39751e-06, 1.339966e-06, 1.356292e-06, 1.339587e-06, 
    1.350205e-06, 1.629551e-06, 1.615153e-06, 1.622926e-06, 1.608321e-06, 
    1.618602e-06, 1.573098e-06, 1.559565e-06, 1.496933e-06, 1.522505e-06, 
    1.481903e-06, 1.51836e-06, 1.51187e-06, 1.480579e-06, 1.516381e-06, 
    1.438596e-06, 1.491124e-06, 1.394239e-06, 1.445954e-06, 1.391026e-06, 
    1.400931e-06, 1.384551e-06, 1.369954e-06, 1.351694e-06, 1.318296e-06, 
    1.325996e-06, 1.298292e-06, 1.593792e-06, 1.575305e-06, 1.576933e-06, 
    1.557681e-06, 1.543509e-06, 1.512994e-06, 1.464614e-06, 1.482726e-06, 
    1.449556e-06, 1.442937e-06, 1.493361e-06, 1.462306e-06, 1.562988e-06, 
    1.546517e-06, 1.556318e-06, 1.592328e-06, 1.478538e-06, 1.536468e-06, 
    1.430281e-06, 1.461081e-06, 1.37203e-06, 1.415994e-06, 1.330243e-06, 
    1.294334e-06, 1.260978e-06, 1.222501e-06, 1.56526e-06, 1.577776e-06, 
    1.5554e-06, 1.524667e-06, 1.496406e-06, 1.459193e-06, 1.455412e-06, 
    1.448494e-06, 1.43065e-06, 1.415723e-06, 1.446307e-06, 1.411993e-06, 
    1.5427e-06, 1.473558e-06, 1.582515e-06, 1.54934e-06, 1.526473e-06, 
    1.536489e-06, 1.484803e-06, 1.472735e-06, 1.42415e-06, 1.449176e-06, 
    1.303151e-06, 1.366874e-06, 1.193599e-06, 1.2409e-06, 1.582158e-06, 
    1.565305e-06, 1.507264e-06, 1.534759e-06, 1.456726e-06, 1.437797e-06, 
    1.422496e-06, 1.403038e-06, 1.400947e-06, 1.389484e-06, 1.40829e-06, 
    1.390226e-06, 1.459115e-06, 1.428143e-06, 1.513853e-06, 1.492784e-06, 
    1.502461e-06, 1.513106e-06, 1.480361e-06, 1.445822e-06, 1.445094e-06, 
    1.434099e-06, 1.403309e-06, 1.456414e-06, 1.295019e-06, 1.393654e-06, 
    1.547017e-06, 1.514937e-06, 1.510387e-06, 1.522761e-06, 1.43969e-06, 
    1.469547e-06, 1.389764e-06, 1.411128e-06, 1.376203e-06, 1.393507e-06, 
    1.396061e-06, 1.418451e-06, 1.432471e-06, 1.468171e-06, 1.497511e-06, 
    1.520964e-06, 1.515497e-06, 1.489784e-06, 1.443723e-06, 1.400755e-06, 
    1.410116e-06, 1.378843e-06, 1.462323e-06, 1.427043e-06, 1.440631e-06, 
    1.405326e-06, 1.483207e-06, 1.416748e-06, 1.500412e-06, 1.492991e-06, 
    1.470143e-06, 1.424661e-06, 1.414695e-06, 1.404078e-06, 1.410626e-06, 
    1.442563e-06, 1.447829e-06, 1.470698e-06, 1.477037e-06, 1.494606e-06, 
    1.509219e-06, 1.495864e-06, 1.481894e-06, 1.442552e-06, 1.407505e-06, 
    1.369745e-06, 1.360579e-06, 1.317184e-06, 1.352452e-06, 1.294478e-06, 
    1.343679e-06, 1.259061e-06, 1.412948e-06, 1.345151e-06, 1.469109e-06, 
    1.455517e-06, 1.431073e-06, 1.375733e-06, 1.405491e-06, 1.370721e-06, 
    1.448036e-06, 1.488898e-06, 1.499561e-06, 1.519532e-06, 1.499105e-06, 
    1.500762e-06, 1.481321e-06, 1.487557e-06, 1.441254e-06, 1.466044e-06, 
    1.396124e-06, 1.370995e-06, 1.301181e-06, 1.259224e-06, 1.217194e-06, 
    1.198854e-06, 1.193298e-06, 1.190979e-06,
  1.526628e-07, 1.468535e-07, 1.479721e-07, 1.433652e-07, 1.4591e-07, 
    1.429092e-07, 1.514741e-07, 1.466254e-07, 1.497097e-07, 1.521346e-07, 
    1.346795e-07, 1.431619e-07, 1.262101e-07, 1.313707e-07, 1.186529e-07, 
    1.270043e-07, 1.170122e-07, 1.188894e-07, 1.132981e-07, 1.148825e-07, 
    1.079149e-07, 1.125715e-07, 1.044129e-07, 1.09016e-07, 1.082873e-07, 
    1.127272e-07, 1.414297e-07, 1.357178e-07, 1.417725e-07, 1.409479e-07, 
    1.413177e-07, 1.458569e-07, 1.481775e-07, 1.53113e-07, 1.522097e-07, 
    1.485886e-07, 1.405781e-07, 1.43267e-07, 1.365518e-07, 1.367013e-07, 
    1.29454e-07, 1.326912e-07, 1.208772e-07, 1.241649e-07, 1.148161e-07, 
    1.171237e-07, 1.149237e-07, 1.155881e-07, 1.149151e-07, 1.183113e-07, 
    1.168485e-07, 1.198653e-07, 1.32081e-07, 1.284134e-07, 1.395429e-07, 
    1.465122e-07, 1.512593e-07, 1.546839e-07, 1.541969e-07, 1.53271e-07, 
    1.485675e-07, 1.442279e-07, 1.409737e-07, 1.388223e-07, 1.367228e-07, 
    1.304865e-07, 1.272605e-07, 1.202188e-07, 1.214716e-07, 1.193546e-07, 
    1.173549e-07, 1.140447e-07, 1.145855e-07, 1.131417e-07, 1.194106e-07, 
    1.152202e-07, 1.221887e-07, 1.202569e-07, 1.36153e-07, 1.425386e-07, 
    1.453057e-07, 1.477566e-07, 1.538231e-07, 1.496175e-07, 1.512668e-07, 
    1.473619e-07, 1.449128e-07, 1.46121e-07, 1.387638e-07, 1.415961e-07, 
    1.270709e-07, 1.332074e-07, 1.17587e-07, 1.212138e-07, 1.167281e-07, 
    1.190038e-07, 1.151213e-07, 1.186119e-07, 1.126075e-07, 1.113259e-07, 
    1.122006e-07, 1.08865e-07, 1.188073e-07, 1.149235e-07, 1.461549e-07, 
    1.459573e-07, 1.450396e-07, 1.491003e-07, 1.493511e-07, 1.531377e-07, 
    1.497658e-07, 1.483436e-07, 1.447719e-07, 1.426839e-07, 1.407166e-07, 
    1.364505e-07, 1.317818e-07, 1.254232e-07, 1.209766e-07, 1.180522e-07, 
    1.198402e-07, 1.182608e-07, 1.200272e-07, 1.208609e-07, 1.118049e-07, 
    1.168348e-07, 1.093408e-07, 1.097473e-07, 1.131074e-07, 1.097015e-07, 
    1.458188e-07, 1.469569e-07, 1.509499e-07, 1.478194e-07, 1.535536e-07, 
    1.503271e-07, 1.484907e-07, 1.41536e-07, 1.400361e-07, 1.386534e-07, 
    1.359481e-07, 1.325243e-07, 1.26649e-07, 1.216726e-07, 1.172393e-07, 
    1.175606e-07, 1.174474e-07, 1.164699e-07, 1.189004e-07, 1.160739e-07, 
    1.156035e-07, 1.168356e-07, 1.098018e-07, 1.117831e-07, 1.09756e-07, 
    1.110431e-07, 1.465864e-07, 1.446776e-07, 1.457071e-07, 1.437748e-07, 
    1.451343e-07, 1.39149e-07, 1.373848e-07, 1.293156e-07, 1.32591e-07, 
    1.274029e-07, 1.320583e-07, 1.312256e-07, 1.272348e-07, 1.318042e-07, 
    1.219433e-07, 1.285753e-07, 1.16432e-07, 1.228654e-07, 1.160361e-07, 
    1.172582e-07, 1.152393e-07, 1.134498e-07, 1.11224e-07, 1.071899e-07, 
    1.081156e-07, 1.047968e-07, 1.418608e-07, 1.394375e-07, 1.396503e-07, 
    1.371398e-07, 1.353012e-07, 1.313697e-07, 1.25214e-07, 1.275072e-07, 
    1.233176e-07, 1.22487e-07, 1.288602e-07, 1.249227e-07, 1.378304e-07, 
    1.356908e-07, 1.369625e-07, 1.416684e-07, 1.269758e-07, 1.343907e-07, 
    1.209039e-07, 1.247682e-07, 1.137038e-07, 1.191248e-07, 1.086274e-07, 
    1.043254e-07, 1.003796e-07, 9.58897e-08, 1.381263e-07, 1.397605e-07, 
    1.368433e-07, 1.328692e-07, 1.292482e-07, 1.245302e-07, 1.240539e-07, 
    1.231843e-07, 1.209499e-07, 1.190911e-07, 1.229097e-07, 1.18628e-07, 
    1.351966e-07, 1.263448e-07, 1.40381e-07, 1.360567e-07, 1.331017e-07, 
    1.343934e-07, 1.277711e-07, 1.262405e-07, 1.201393e-07, 1.232698e-07, 
    1.053765e-07, 1.130734e-07, 9.256075e-08, 9.802844e-08, 1.403341e-07, 
    1.381321e-07, 1.306356e-07, 1.341701e-07, 1.242194e-07, 1.218433e-07, 
    1.199333e-07, 1.175187e-07, 1.172602e-07, 1.158462e-07, 1.181689e-07, 
    1.159375e-07, 1.245203e-07, 1.206371e-07, 1.314799e-07, 1.287866e-07, 
    1.300214e-07, 1.313841e-07, 1.27207e-07, 1.228488e-07, 1.227575e-07, 
    1.213807e-07, 1.175524e-07, 1.241801e-07, 1.044071e-07, 1.1636e-07, 
    1.357555e-07, 1.31619e-07, 1.310355e-07, 1.326239e-07, 1.220802e-07, 
    1.258372e-07, 1.158806e-07, 1.185207e-07, 1.142148e-07, 1.163418e-07, 
    1.166568e-07, 1.194301e-07, 1.211773e-07, 1.256633e-07, 1.293893e-07, 
    1.323929e-07, 1.316907e-07, 1.284047e-07, 1.225855e-07, 1.172365e-07, 
    1.183952e-07, 1.145385e-07, 1.249248e-07, 1.204999e-07, 1.22198e-07, 
    1.178019e-07, 1.275684e-07, 1.192186e-07, 1.297595e-07, 1.28813e-07, 
    1.259126e-07, 1.20203e-07, 1.189633e-07, 1.176474e-07, 1.184585e-07, 
    1.224401e-07, 1.231007e-07, 1.259827e-07, 1.267855e-07, 1.290188e-07, 
    1.308859e-07, 1.291791e-07, 1.274017e-07, 1.224387e-07, 1.180716e-07, 
    1.134243e-07, 1.123052e-07, 1.070565e-07, 1.113162e-07, 1.043427e-07, 
    1.102517e-07, 1.001545e-07, 1.187467e-07, 1.1043e-07, 1.257818e-07, 
    1.240672e-07, 1.210027e-07, 1.141573e-07, 1.178223e-07, 1.135436e-07, 
    1.231267e-07, 1.282918e-07, 1.296509e-07, 1.322089e-07, 1.295927e-07, 
    1.298043e-07, 1.273289e-07, 1.281212e-07, 1.222761e-07, 1.253945e-07, 
    1.166646e-07, 1.135772e-07, 1.051413e-07, 1.001736e-07, 9.527559e-08, 
    9.316314e-08, 9.252631e-08, 9.226089e-08,
  4.407835e-09, 4.171025e-09, 4.21634e-09, 4.030609e-09, 4.132911e-09, 
    4.012351e-09, 4.359083e-09, 4.161804e-09, 4.286998e-09, 4.386151e-09, 
    3.686933e-09, 4.022465e-09, 3.360266e-09, 3.558295e-09, 3.076124e-09, 
    3.390533e-09, 3.015382e-09, 3.08491e-09, 2.879142e-09, 2.937043e-09, 
    2.684889e-09, 2.8527e-09, 2.560597e-09, 2.724306e-09, 2.698199e-09, 
    2.858359e-09, 3.95328e-09, 3.727563e-09, 3.966947e-09, 3.934098e-09, 
    3.948819e-09, 4.13077e-09, 4.224673e-09, 4.426338e-09, 4.389234e-09, 
    4.241369e-09, 3.919391e-09, 4.026675e-09, 3.760283e-09, 3.766156e-09, 
    3.484374e-09, 3.609476e-09, 3.159018e-09, 3.282671e-09, 2.93461e-09, 
    3.019496e-09, 2.938555e-09, 2.962933e-09, 2.938238e-09, 3.063447e-09, 
    3.009337e-09, 3.121231e-09, 3.5858e-09, 3.444423e-09, 3.878305e-09, 
    4.157229e-09, 4.350288e-09, 4.491076e-09, 4.470978e-09, 4.432838e-09, 
    4.240514e-09, 4.065206e-09, 3.935122e-09, 3.84978e-09, 3.767e-09, 
    3.524141e-09, 3.400313e-09, 3.134418e-09, 3.181273e-09, 3.102207e-09, 
    3.028038e-09, 2.906387e-09, 2.926165e-09, 2.873446e-09, 3.104289e-09, 
    2.949426e-09, 3.208182e-09, 3.13584e-09, 3.744628e-09, 3.997533e-09, 
    4.108556e-09, 4.207599e-09, 4.455567e-09, 4.283242e-09, 4.350595e-09, 
    4.191601e-09, 4.092739e-09, 4.141429e-09, 3.847466e-09, 3.959912e-09, 
    3.393073e-09, 3.629542e-09, 3.036622e-09, 3.171616e-09, 3.004896e-09, 
    3.08916e-09, 2.945799e-09, 3.0746e-09, 2.854008e-09, 2.807532e-09, 
    2.839231e-09, 2.718891e-09, 3.081856e-09, 2.938547e-09, 4.142794e-09, 
    4.134823e-09, 4.097841e-09, 4.262179e-09, 4.272388e-09, 4.427354e-09, 
    4.289281e-09, 4.231418e-09, 4.087068e-09, 4.003341e-09, 3.924898e-09, 
    3.756305e-09, 3.574208e-09, 3.330351e-09, 3.162736e-09, 3.053845e-09, 
    3.120293e-09, 3.061575e-09, 3.127266e-09, 3.158406e-09, 2.824876e-09, 
    3.008831e-09, 2.735967e-09, 2.750579e-09, 2.872198e-09, 2.74893e-09, 
    4.129233e-09, 4.175208e-09, 4.337631e-09, 4.210146e-09, 4.444469e-09, 
    4.312181e-09, 4.237392e-09, 3.957518e-09, 3.897866e-09, 3.843102e-09, 
    3.736585e-09, 3.602996e-09, 3.376983e-09, 3.188812e-09, 3.023766e-09, 
    3.035646e-09, 3.031459e-09, 2.995376e-09, 3.085318e-09, 2.980795e-09, 
    2.9635e-09, 3.008862e-09, 2.75254e-09, 2.824086e-09, 2.75089e-09, 
    2.797304e-09, 4.160226e-09, 4.083279e-09, 4.124729e-09, 4.047025e-09, 
    4.101651e-09, 3.862706e-09, 3.793051e-09, 3.479053e-09, 3.605587e-09, 
    3.405751e-09, 3.584919e-09, 3.552684e-09, 3.399335e-09, 3.575074e-09, 
    3.19897e-09, 3.45063e-09, 2.99398e-09, 3.233639e-09, 2.979402e-09, 
    3.024466e-09, 2.950127e-09, 2.884672e-09, 2.803843e-09, 2.659017e-09, 
    2.692061e-09, 2.574139e-09, 3.970468e-09, 3.874129e-09, 3.882561e-09, 
    3.783403e-09, 3.711242e-09, 3.558255e-09, 3.322407e-09, 3.409737e-09, 
    3.250676e-09, 3.219396e-09, 3.461557e-09, 3.311361e-09, 3.81061e-09, 
    3.7265e-09, 3.776429e-09, 3.962797e-09, 3.389446e-09, 3.675653e-09, 
    3.160015e-09, 3.305506e-09, 2.893938e-09, 3.093658e-09, 2.710375e-09, 
    2.557516e-09, 2.419544e-09, 2.265224e-09, 3.822282e-09, 3.88693e-09, 
    3.771738e-09, 3.616394e-09, 3.476463e-09, 3.296494e-09, 3.278475e-09, 
    3.245648e-09, 3.161738e-09, 3.092403e-09, 3.235303e-09, 3.075197e-09, 
    3.707151e-09, 3.365392e-09, 3.911559e-09, 3.740848e-09, 3.625428e-09, 
    3.675757e-09, 3.419827e-09, 3.36142e-09, 3.13145e-09, 3.248872e-09, 
    2.594632e-09, 2.870962e-09, 2.152691e-09, 2.338373e-09, 3.909697e-09, 
    3.822511e-09, 3.529894e-09, 3.66704e-09, 3.284732e-09, 3.195213e-09, 
    3.123763e-09, 3.034095e-09, 3.024538e-09, 2.972418e-09, 3.058168e-09, 
    2.975778e-09, 3.296118e-09, 3.15004e-09, 3.562518e-09, 3.458734e-09, 
    3.50621e-09, 3.558811e-09, 3.398269e-09, 3.233013e-09, 3.229572e-09, 
    3.177868e-09, 3.035348e-09, 3.283245e-09, 2.560396e-09, 2.991334e-09, 
    3.729034e-09, 3.567905e-09, 3.545338e-09, 3.606863e-09, 3.204107e-09, 
    3.34608e-09, 2.973684e-09, 3.071216e-09, 2.912604e-09, 2.990658e-09, 
    3.002267e-09, 3.105016e-09, 3.17025e-09, 3.339468e-09, 3.481884e-09, 
    3.597896e-09, 3.570678e-09, 3.444086e-09, 3.223102e-09, 3.023662e-09, 
    3.066562e-09, 2.924445e-09, 3.31144e-09, 3.144915e-09, 3.208535e-09, 
    3.044572e-09, 3.412074e-09, 3.097153e-09, 3.496126e-09, 3.459748e-09, 
    3.348943e-09, 3.133828e-09, 3.087655e-09, 3.038856e-09, 3.068906e-09, 
    3.217634e-09, 3.242498e-09, 3.351612e-09, 3.382185e-09, 3.467647e-09, 
    3.539554e-09, 3.473807e-09, 3.405705e-09, 3.21758e-09, 3.054565e-09, 
    2.883744e-09, 2.843028e-09, 2.654268e-09, 2.80718e-09, 2.558126e-09, 
    2.768745e-09, 2.411743e-09, 3.079608e-09, 2.775169e-09, 3.343971e-09, 
    3.278977e-09, 3.163716e-09, 2.910502e-09, 3.045329e-09, 2.888097e-09, 
    3.243477e-09, 3.439764e-09, 3.491944e-09, 3.590759e-09, 3.489708e-09, 
    3.49785e-09, 3.402923e-09, 3.433225e-09, 3.211466e-09, 3.329259e-09, 
    3.002553e-09, 2.889321e-09, 2.58631e-09, 2.412401e-09, 2.24434e-09, 
    2.172933e-09, 2.151535e-09, 2.142635e-09,
  3.551892e-11, 3.275957e-11, 3.328299e-11, 3.115183e-11, 3.232105e-11, 
    3.094438e-11, 3.494603e-11, 3.265334e-11, 3.410351e-11, 3.52638e-11, 
    2.73103e-11, 3.105925e-11, 2.378899e-11, 2.590797e-11, 2.083682e-11, 
    2.410967e-11, 2.021983e-11, 2.092647e-11, 1.885477e-11, 1.943169e-11, 
    1.695514e-11, 1.859292e-11, 1.576969e-11, 1.733604e-11, 1.708349e-11, 
    1.864887e-11, 3.027572e-11, 2.775733e-11, 3.043007e-11, 3.005943e-11, 
    3.022538e-11, 3.229646e-11, 3.33795e-11, 3.5737e-11, 3.530005e-11, 
    3.357304e-11, 2.989389e-11, 3.11071e-11, 2.811871e-11, 2.818371e-11, 
    2.511126e-11, 2.646351e-11, 2.168696e-11, 2.297223e-11, 1.940735e-11, 
    2.026145e-11, 1.944681e-11, 1.969119e-11, 1.944364e-11, 2.070763e-11, 
    2.015869e-11, 2.129827e-11, 2.620612e-11, 2.46835e-11, 2.94327e-11, 
    3.260068e-11, 3.484295e-11, 3.650274e-11, 3.626456e-11, 3.581368e-11, 
    3.356312e-11, 3.154596e-11, 3.007096e-11, 2.911365e-11, 2.819306e-11, 
    2.553905e-11, 2.421353e-11, 2.14337e-11, 2.191678e-11, 2.110332e-11, 
    2.034795e-11, 1.912564e-11, 1.932293e-11, 1.879828e-11, 2.112462e-11, 
    1.955569e-11, 2.219555e-11, 2.144831e-11, 2.794568e-11, 3.077626e-11, 
    3.204167e-11, 3.318186e-11, 3.608221e-11, 3.405976e-11, 3.484655e-11, 
    3.299696e-11, 3.186055e-11, 3.24189e-11, 2.90878e-11, 3.035059e-11, 
    2.413663e-11, 2.668219e-11, 2.043498e-11, 2.181698e-11, 2.011382e-11, 
    2.096988e-11, 1.951934e-11, 2.082127e-11, 1.860584e-11, 1.814797e-11, 
    1.845992e-11, 1.728357e-11, 2.089529e-11, 1.944674e-11, 3.24346e-11, 
    3.2343e-11, 3.191893e-11, 3.38147e-11, 3.393342e-11, 3.574898e-11, 
    3.413012e-11, 3.345765e-11, 3.179567e-11, 3.084212e-11, 2.995584e-11, 
    2.80747e-11, 2.608035e-11, 2.347318e-11, 2.172531e-11, 2.060992e-11, 
    2.128864e-11, 2.068856e-11, 2.136021e-11, 2.168065e-11, 1.831848e-11, 
    2.015358e-11, 1.744917e-11, 1.759123e-11, 1.878591e-11, 1.757518e-11, 
    3.227881e-11, 3.280779e-11, 3.469474e-11, 3.321131e-11, 3.595102e-11, 
    3.439723e-11, 3.352691e-11, 3.032356e-11, 2.965202e-11, 2.903909e-11, 
    2.785682e-11, 2.639299e-11, 2.396595e-11, 2.19948e-11, 2.030467e-11, 
    2.042508e-11, 2.038262e-11, 2.001773e-11, 2.093064e-11, 1.987079e-11, 
    1.969689e-11, 2.01539e-11, 1.761032e-11, 1.831069e-11, 1.759426e-11, 
    1.804764e-11, 3.263516e-11, 3.175235e-11, 3.222711e-11, 3.133867e-11, 
    3.196255e-11, 2.925812e-11, 2.848192e-11, 2.505418e-11, 2.642118e-11, 
    2.427134e-11, 2.619656e-11, 2.584726e-11, 2.420315e-11, 2.608973e-11, 
    2.210002e-11, 2.474984e-11, 2.000365e-11, 2.246018e-11, 1.985677e-11, 
    2.031176e-11, 1.956271e-11, 1.890966e-11, 1.811177e-11, 1.67064e-11, 
    1.702426e-11, 1.589767e-11, 3.046987e-11, 2.938594e-11, 2.948037e-11, 
    2.837484e-11, 2.75775e-11, 2.590753e-11, 2.338951e-11, 2.431372e-11, 
    2.263773e-11, 2.231201e-11, 2.48667e-11, 2.327331e-11, 2.867705e-11, 
    2.774559e-11, 2.829752e-11, 3.038318e-11, 2.409813e-11, 2.718652e-11, 
    2.169724e-11, 2.321178e-11, 1.900173e-11, 2.101587e-11, 1.720114e-11, 
    1.574062e-11, 1.445412e-11, 1.30527e-11, 2.880696e-11, 2.952935e-11, 
    2.824553e-11, 2.653885e-11, 2.502639e-11, 2.311715e-11, 2.292829e-11, 
    2.258529e-11, 2.171502e-11, 2.100303e-11, 2.24775e-11, 2.082736e-11, 
    2.753251e-11, 2.384321e-11, 2.980582e-11, 2.79039e-11, 2.663732e-11, 
    2.718765e-11, 2.442112e-11, 2.380118e-11, 2.14032e-11, 2.261891e-11, 
    1.609191e-11, 1.877367e-11, 1.205688e-11, 1.371193e-11, 2.978489e-11, 
    2.880951e-11, 2.560108e-11, 2.709211e-11, 2.299382e-11, 2.206109e-11, 
    2.132425e-11, 2.040936e-11, 2.031249e-11, 1.978651e-11, 2.065388e-11, 
    1.98203e-11, 2.311321e-11, 2.159443e-11, 2.595367e-11, 2.483649e-11, 
    2.534589e-11, 2.591355e-11, 2.419179e-11, 2.245366e-11, 2.241783e-11, 
    2.188159e-11, 2.04221e-11, 2.297824e-11, 1.576782e-11, 1.9977e-11, 
    2.777352e-11, 2.601205e-11, 2.576783e-11, 2.643506e-11, 2.215328e-11, 
    2.363907e-11, 1.979924e-11, 2.078677e-11, 1.918759e-11, 1.997015e-11, 
    2.008727e-11, 2.113207e-11, 2.180287e-11, 2.35693e-11, 2.508454e-11, 
    2.633752e-11, 2.604208e-11, 2.46799e-11, 2.235055e-11, 2.030363e-11, 
    2.073935e-11, 1.930575e-11, 2.327414e-11, 2.154167e-11, 2.219922e-11, 
    2.051568e-11, 2.43386e-11, 2.105163e-11, 2.523746e-11, 2.484734e-11, 
    2.366931e-11, 2.142764e-11, 2.095451e-11, 2.045766e-11, 2.076323e-11, 
    2.229371e-11, 2.255246e-11, 2.369749e-11, 2.40211e-11, 2.493191e-11, 
    2.570534e-11, 2.499792e-11, 2.427084e-11, 2.229315e-11, 2.061724e-11, 
    1.890045e-11, 1.849738e-11, 1.666087e-11, 1.814454e-11, 1.57464e-11, 
    1.776834e-11, 1.438233e-11, 2.087238e-11, 1.783104e-11, 2.361681e-11, 
    2.293354e-11, 2.173543e-11, 1.916665e-11, 2.052337e-11, 1.894369e-11, 
    2.256266e-11, 2.463375e-11, 2.519253e-11, 2.625998e-11, 2.516851e-11, 
    2.5256e-11, 2.424126e-11, 2.456394e-11, 2.222965e-11, 2.346167e-11, 
    2.009016e-11, 1.895585e-11, 1.601295e-11, 1.438837e-11, 1.286619e-11, 
    1.223432e-11, 1.204676e-11, 1.196899e-11,
  4.485717e-14, 3.795889e-14, 3.923833e-14, 3.411792e-14, 3.689776e-14, 
    3.363232e-14, 4.339431e-14, 3.770095e-14, 4.127178e-14, 4.420377e-14, 
    2.552042e-14, 3.390091e-14, 1.843828e-14, 2.260232e-14, 1.317501e-14, 
    1.904871e-14, 1.216106e-14, 1.332491e-14, 1.003205e-14, 1.091217e-14, 
    7.349246e-15, 9.642337e-15, 5.853651e-15, 7.859727e-15, 7.519674e-15, 
    9.7251e-15, 3.208312e-14, 2.647642e-14, 3.243854e-14, 3.158733e-14, 
    3.19675e-14, 3.683858e-14, 3.94758e-14, 4.541807e-14, 4.42964e-14, 
    3.99533e-14, 3.120962e-14, 3.401297e-14, 2.725799e-14, 2.739943e-14, 
    2.100105e-14, 2.374337e-14, 1.46224e-14, 1.691673e-14, 1.087445e-14, 
    1.222845e-14, 1.093564e-14, 1.131753e-14, 1.093072e-14, 1.29601e-14, 
    1.20623e-14, 1.395351e-14, 2.321225e-14, 2.015883e-14, 3.01655e-14, 
    3.757332e-14, 4.313279e-14, 4.740537e-14, 4.678431e-14, 4.561587e-14, 
    3.992878e-14, 3.504682e-14, 3.161365e-14, 2.945025e-14, 2.74198e-14, 
    2.185569e-14, 1.924794e-14, 1.418524e-14, 1.502343e-14, 1.362254e-14, 
    1.236901e-14, 1.044163e-14, 1.074403e-14, 9.947459e-15, 1.365855e-14, 
    1.110517e-14, 1.551532e-14, 1.42103e-14, 2.688286e-14, 3.324048e-14, 
    3.622701e-14, 3.899003e-14, 4.63106e-14, 4.116253e-14, 4.314191e-14, 
    3.85374e-14, 3.579426e-14, 3.713367e-14, 2.939257e-14, 3.225534e-14, 
    1.910034e-14, 2.419796e-14, 1.251107e-14, 1.484878e-14, 1.199001e-14, 
    1.339773e-14, 1.104846e-14, 1.314905e-14, 9.661437e-15, 8.994432e-15, 
    9.44678e-15, 7.788543e-15, 1.327269e-14, 1.093555e-14, 3.717157e-14, 
    3.695064e-14, 3.593353e-14, 4.055222e-14, 4.08475e-14, 4.544896e-14, 
    4.133827e-14, 3.966835e-14, 3.563968e-14, 3.339379e-14, 3.135078e-14, 
    2.71624e-14, 2.295427e-14, 1.784426e-14, 1.468903e-14, 1.279847e-14, 
    1.39371e-14, 1.292849e-14, 1.405931e-14, 1.461144e-14, 9.240576e-15, 
    1.205406e-14, 8.014055e-15, 8.209605e-15, 9.928974e-15, 8.187415e-15, 
    3.679609e-14, 3.807614e-14, 4.275763e-14, 3.906226e-14, 4.597077e-14, 
    4.200782e-14, 3.983932e-14, 3.219317e-14, 3.066051e-14, 2.928397e-14, 
    2.669073e-14, 2.359742e-14, 1.877421e-14, 1.51605e-14, 1.229861e-14, 
    1.249486e-14, 1.242553e-14, 1.183578e-14, 1.333189e-14, 1.160145e-14, 
    1.132651e-14, 1.205456e-14, 8.236028e-15, 9.229264e-15, 8.213795e-15, 
    8.850831e-15, 3.76568e-14, 3.553661e-14, 3.667175e-14, 3.455723e-14, 
    3.603775e-14, 2.977343e-14, 2.805159e-14, 2.088798e-14, 2.365574e-14, 
    1.935914e-14, 2.319259e-14, 2.247884e-14, 1.922801e-14, 2.297345e-14, 
    1.534612e-14, 2.028867e-14, 1.181325e-14, 1.59878e-14, 1.157919e-14, 
    1.231013e-14, 1.111612e-14, 1.011453e-14, 8.9425e-15, 7.02359e-15, 
    7.440802e-15, 6.00813e-15, 3.253039e-14, 3.006031e-14, 3.027284e-14, 
    2.781679e-14, 2.609027e-14, 2.260142e-14, 1.768807e-14, 1.944081e-14, 
    1.630766e-14, 1.572258e-14, 2.0518e-14, 1.747201e-14, 2.848111e-14, 
    2.645108e-14, 2.764769e-14, 3.233043e-14, 1.902659e-14, 2.52578e-14, 
    1.464026e-14, 1.735799e-14, 1.025347e-14, 1.347506e-14, 7.677303e-15, 
    5.818811e-15, 4.368243e-15, 3.003348e-15, 2.876831e-14, 3.038329e-14, 
    2.753418e-14, 2.389966e-14, 2.083297e-14, 1.718319e-14, 1.683625e-14, 
    1.621293e-14, 1.467113e-14, 1.345343e-14, 1.601887e-14, 1.315919e-14, 
    2.599407e-14, 1.854097e-14, 3.100928e-14, 2.679246e-14, 2.410444e-14, 
    2.526018e-14, 1.964837e-14, 1.846131e-14, 1.413293e-14, 1.627363e-14, 
    6.245907e-15, 9.910715e-15, 2.179756e-15, 3.61635e-15, 3.096174e-14, 
    2.877395e-14, 2.198055e-14, 2.505817e-14, 1.695633e-14, 1.527732e-14, 
    1.399785e-14, 1.246918e-14, 1.231132e-14, 1.146789e-14, 1.28711e-14, 
    1.152135e-14, 1.717592e-14, 1.446209e-14, 2.269542e-14, 2.045863e-14, 
    2.146825e-14, 2.261366e-14, 1.920613e-14, 1.597606e-14, 1.591178e-14, 
    1.496176e-14, 1.249008e-14, 1.692775e-14, 5.851449e-15, 1.177072e-14, 
    2.651115e-14, 2.28146e-14, 2.231761e-14, 2.368445e-14, 1.544036e-14, 
    1.815539e-14, 1.148802e-14, 1.309157e-14, 1.053621e-14, 1.17597e-14, 
    1.194732e-14, 1.367114e-14, 1.482415e-14, 1.802428e-14, 2.094809e-14, 
    2.348285e-14, 2.287594e-14, 2.015179e-14, 1.579141e-14, 1.229693e-14, 
    1.301274e-14, 1.071756e-14, 1.747353e-14, 1.4371e-14, 1.552186e-14, 
    1.264334e-14, 1.948882e-14, 1.353535e-14, 2.125188e-14, 2.047993e-14, 
    1.821231e-14, 1.417485e-14, 1.337192e-14, 1.254819e-14, 1.305241e-14, 
    1.568996e-14, 1.615372e-14, 1.826542e-14, 1.887934e-14, 2.06464e-14, 
    2.219108e-14, 2.077667e-14, 1.935818e-14, 1.568894e-14, 1.281057e-14, 
    1.010068e-14, 9.501699e-15, 6.964675e-15, 8.989521e-15, 5.825771e-15, 
    8.456168e-15, 4.292765e-15, 1.323441e-14, 8.54412e-15, 1.811351e-14, 
    1.684586e-14, 1.470666e-14, 1.050424e-14, 1.265596e-14, 1.016581e-14, 
    1.617211e-14, 2.006169e-14, 2.116245e-14, 2.332302e-14, 2.111471e-14, 
    2.128881e-14, 1.930121e-14, 1.992564e-14, 1.55759e-14, 1.782272e-14, 
    1.195197e-14, 1.018414e-14, 6.148757e-15, 4.299076e-15, 2.839554e-15, 
    2.317233e-15, 2.172036e-15, 2.113177e-15,
  1.51744e-19, 1.286883e-19, 1.329689e-19, 1.158245e-19, 1.251365e-19, 
    1.141967e-19, 1.468595e-19, 1.278251e-19, 1.397679e-19, 1.495626e-19, 
    8.694903e-20, 1.150971e-19, 6.305827e-20, 7.711833e-20, 4.52239e-20, 
    6.5122e-20, 4.177787e-20, 4.573304e-20, 3.452882e-20, 3.752786e-20, 
    2.536346e-20, 3.319971e-20, 2.023541e-20, 2.711047e-20, 2.594689e-20, 
    3.348203e-20, 1.090012e-19, 9.016607e-20, 1.101934e-19, 1.073377e-19, 
    1.086133e-19, 1.249384e-19, 1.337632e-19, 1.536161e-19, 1.498718e-19, 
    1.353601e-19, 1.060701e-19, 1.154727e-19, 9.279489e-20, 9.327051e-20, 
    7.17163e-20, 8.096442e-20, 5.013672e-20, 5.79105e-20, 3.739939e-20, 
    4.200702e-20, 3.760778e-20, 3.890801e-20, 3.759104e-20, 4.449381e-20, 
    4.1442e-20, 4.786722e-20, 7.917452e-20, 6.887269e-20, 1.02565e-19, 
    1.273979e-19, 1.45986e-19, 1.602466e-19, 1.58175e-19, 1.542763e-19, 
    1.352781e-19, 1.189373e-19, 1.07426e-19, 1.001629e-19, 9.333902e-20, 
    7.46002e-20, 6.579534e-20, 4.865364e-20, 5.149666e-20, 4.674369e-20, 
    4.248494e-20, 3.592489e-20, 3.695517e-20, 3.424037e-20, 4.686596e-20, 
    3.818504e-20, 5.316406e-20, 4.873868e-20, 9.153326e-20, 1.128829e-19, 
    1.228906e-19, 1.321384e-19, 1.565945e-19, 1.394028e-19, 1.460165e-19, 
    1.306241e-19, 1.214412e-19, 1.259263e-19, 9.996909e-20, 1.095789e-19, 
    6.529649e-20, 8.249594e-20, 4.296785e-20, 5.090447e-20, 4.119615e-20, 
    4.598033e-20, 3.799196e-20, 4.513571e-20, 3.326487e-20, 3.098844e-20, 
    3.25325e-20, 2.686695e-20, 4.555567e-20, 3.760746e-20, 1.260531e-19, 
    1.253135e-19, 1.219077e-19, 1.373626e-19, 1.383498e-19, 1.537192e-19, 
    1.399902e-19, 1.344072e-19, 1.209235e-19, 1.133969e-19, 1.065438e-19, 
    9.247343e-20, 7.830494e-20, 6.104909e-20, 5.03627e-20, 4.394462e-20, 
    4.781151e-20, 4.438641e-20, 4.822627e-20, 5.009953e-20, 3.182876e-20, 
    4.1414e-20, 2.763832e-20, 2.830697e-20, 3.417734e-20, 2.82311e-20, 
    1.247961e-19, 1.290807e-19, 1.447328e-19, 1.3238e-19, 1.554606e-19, 
    1.422277e-19, 1.349789e-19, 1.093703e-19, 1.04227e-19, 9.960429e-20, 
    9.088701e-20, 8.047265e-20, 6.41941e-20, 5.196138e-20, 4.224557e-20, 
    4.291276e-20, 4.267706e-20, 4.067155e-20, 4.575674e-20, 3.987427e-20, 
    3.893857e-20, 4.141568e-20, 2.83973e-20, 3.179015e-20, 2.832129e-20, 
    3.049805e-20, 1.276773e-19, 1.205782e-19, 1.243798e-19, 1.172968e-19, 
    1.222567e-19, 1.012483e-19, 9.546307e-20, 7.133464e-20, 8.066915e-20, 
    6.617111e-20, 7.910826e-20, 7.670196e-20, 6.572798e-20, 7.836958e-20, 
    5.259062e-20, 6.931118e-20, 4.059489e-20, 5.476495e-20, 3.979852e-20, 
    4.228476e-20, 3.822233e-20, 3.481001e-20, 3.08111e-20, 2.424814e-20, 
    2.567691e-20, 2.076581e-20, 1.105015e-19, 1.022118e-19, 1.029254e-19, 
    9.467374e-20, 8.886684e-20, 7.71153e-20, 6.052066e-20, 6.644712e-20, 
    5.584834e-20, 5.386641e-20, 7.008557e-20, 5.978962e-20, 9.69067e-20, 
    9.008081e-20, 9.410525e-20, 1.098308e-19, 6.504722e-20, 8.606501e-20, 
    5.019728e-20, 5.940381e-20, 3.528364e-20, 4.624293e-20, 2.648634e-20, 
    2.011576e-20, 1.512521e-20, 1.041016e-20, 9.787181e-20, 1.032962e-19, 
    9.372361e-20, 8.149104e-20, 7.114896e-20, 5.881232e-20, 5.763807e-20, 
    5.552751e-20, 5.030199e-20, 4.616949e-20, 5.48702e-20, 4.517018e-20, 
    8.854313e-20, 6.340549e-20, 1.053977e-19, 9.12292e-20, 8.21809e-20, 
    8.607301e-20, 6.714842e-20, 6.313615e-20, 4.847614e-20, 5.57331e-20, 
    2.158187e-20, 3.411507e-20, 7.552855e-21, 1.253041e-20, 1.052381e-19, 
    9.789076e-20, 7.502142e-20, 8.53929e-20, 5.804454e-20, 5.235739e-20, 
    4.80177e-20, 4.282547e-20, 4.228878e-20, 3.941975e-20, 4.419142e-20, 
    3.960171e-20, 5.878772e-20, 4.959293e-20, 7.743227e-20, 6.98851e-20, 
    7.329304e-20, 7.715656e-20, 6.565404e-20, 5.47252e-20, 5.450743e-20, 
    5.128758e-20, 4.289649e-20, 5.79478e-20, 2.022785e-20, 4.045018e-20, 
    9.028293e-20, 7.783406e-20, 7.615827e-20, 8.076588e-20, 5.291e-20, 
    6.210154e-20, 3.948826e-20, 4.494046e-20, 3.624719e-20, 4.041271e-20, 
    4.105094e-20, 4.69087e-20, 5.082094e-20, 6.16581e-20, 7.153755e-20, 
    8.008654e-20, 7.804086e-20, 6.884892e-20, 5.409961e-20, 4.223986e-20, 
    4.467268e-20, 3.6865e-20, 5.979473e-20, 4.928391e-20, 5.318624e-20, 
    4.341743e-20, 6.660932e-20, 4.644765e-20, 7.256289e-20, 6.995705e-20, 
    6.229406e-20, 4.861839e-20, 4.589269e-20, 4.309403e-20, 4.480743e-20, 
    5.375586e-20, 5.532698e-20, 6.247368e-20, 6.45495e-20, 7.051909e-20, 
    7.573153e-20, 7.095891e-20, 6.616788e-20, 5.375243e-20, 4.398573e-20, 
    3.476279e-20, 3.271989e-20, 2.40463e-20, 3.097167e-20, 2.013967e-20, 
    2.914974e-20, 1.4865e-20, 4.542566e-20, 2.945029e-20, 6.19599e-20, 
    5.767061e-20, 5.042249e-20, 3.613822e-20, 4.346034e-20, 3.498482e-20, 
    5.538925e-20, 6.854463e-20, 7.226106e-20, 7.954787e-20, 7.209993e-20, 
    7.268751e-20, 6.597538e-20, 6.808507e-20, 5.336936e-20, 6.097623e-20, 
    4.106675e-20, 3.504732e-20, 2.12485e-20, 1.488676e-20, 9.842769e-21, 
    8.030605e-21, 7.526016e-21, 7.321354e-21,
  1.114151e-25, 9.456576e-26, 9.769499e-26, 8.515911e-26, 9.196894e-26, 
    8.396845e-26, 1.078464e-25, 9.393464e-26, 1.026644e-25, 1.098214e-25, 
    6.402566e-26, 8.462706e-26, 4.651485e-26, 5.682357e-26, 3.341952e-26, 
    4.802864e-26, 3.088625e-26, 3.379371e-26, 2.555337e-26, 2.776036e-26, 
    1.880127e-26, 2.457494e-26, 1.501728e-26, 2.008926e-26, 1.923146e-26, 
    2.47828e-26, 8.016771e-26, 6.638163e-26, 8.104e-26, 7.895063e-26, 
    7.988392e-26, 9.182406e-26, 9.827558e-26, 1.127828e-25, 1.100473e-25, 
    9.944279e-26, 7.802315e-26, 8.490182e-26, 6.830651e-26, 6.865475e-26, 
    5.286408e-26, 5.964178e-26, 3.702929e-26, 4.273748e-26, 2.766584e-26, 
    3.105474e-26, 2.781916e-26, 2.877567e-26, 2.780684e-26, 3.28829e-26, 
    3.063929e-26, 3.536199e-26, 5.833032e-26, 5.077922e-26, 7.545821e-26, 
    9.362236e-26, 1.072082e-25, 1.176261e-25, 1.161129e-25, 1.13265e-25, 
    9.938287e-26, 8.74358e-26, 7.901525e-26, 7.370017e-26, 6.87049e-26, 
    5.497806e-26, 4.852249e-26, 3.593978e-26, 3.802819e-26, 3.453642e-26, 
    3.140612e-26, 2.658087e-26, 2.733899e-26, 2.534105e-26, 3.462627e-26, 
    2.824384e-26, 3.925274e-26, 3.600226e-26, 6.738275e-26, 8.300746e-26, 
    9.032672e-26, 9.708786e-26, 1.149585e-25, 1.023975e-25, 1.072305e-25, 
    9.598093e-26, 8.92669e-26, 9.254638e-26, 7.355834e-26, 8.059041e-26, 
    4.815662e-26, 6.07638e-26, 3.176116e-26, 3.759323e-26, 3.04585e-26, 
    3.397545e-26, 2.81018e-26, 3.33547e-26, 2.462292e-26, 2.294661e-26, 
    2.408369e-26, 1.990976e-26, 3.366336e-26, 2.781892e-26, 9.263916e-26, 
    9.209839e-26, 8.9608e-26, 1.009065e-25, 1.016279e-25, 1.128581e-25, 
    1.028268e-25, 9.874628e-26, 8.888826e-26, 8.338348e-26, 7.83698e-26, 
    6.807115e-26, 5.769313e-26, 4.504083e-26, 3.719529e-26, 3.247922e-26, 
    3.532105e-26, 3.280396e-26, 3.56258e-26, 3.700198e-26, 2.356548e-26, 
    3.061869e-26, 2.047833e-26, 2.09711e-26, 2.529465e-26, 2.09152e-26, 
    9.172006e-26, 9.485261e-26, 1.062925e-25, 9.726448e-26, 1.141302e-25, 
    1.044619e-25, 9.916422e-26, 8.043782e-26, 7.667445e-26, 7.329133e-26, 
    6.690955e-26, 5.928147e-26, 4.734804e-26, 3.836951e-26, 3.123013e-26, 
    3.172066e-26, 3.154737e-26, 3.007272e-26, 3.381113e-26, 2.948638e-26, 
    2.879814e-26, 3.061993e-26, 2.103767e-26, 2.353705e-26, 2.098166e-26, 
    2.25854e-26, 9.382664e-26, 8.863577e-26, 9.141565e-26, 8.623598e-26, 
    8.986323e-26, 7.449461e-26, 7.025996e-26, 5.258428e-26, 5.942545e-26, 
    4.879809e-26, 5.828176e-26, 5.651844e-26, 4.84731e-26, 5.77405e-26, 
    3.883162e-26, 5.110074e-26, 3.001635e-26, 4.042825e-26, 2.943066e-26, 
    3.125894e-26, 2.827127e-26, 2.576035e-26, 2.281599e-26, 1.797871e-26, 
    1.90324e-26, 1.540892e-26, 8.126538e-26, 7.519972e-26, 7.572198e-26, 
    6.968209e-26, 6.54302e-26, 5.682135e-26, 4.465311e-26, 4.900051e-26, 
    4.122367e-26, 3.976848e-26, 5.166853e-26, 4.411667e-26, 7.131676e-26, 
    6.631919e-26, 6.926589e-26, 8.077469e-26, 4.797379e-26, 6.337819e-26, 
    3.707378e-26, 4.383353e-26, 2.610894e-26, 3.416844e-26, 1.962918e-26, 
    1.492893e-26, 1.124038e-26, 7.747884e-27, 7.202323e-26, 7.599336e-26, 
    6.898648e-26, 6.002759e-26, 5.244816e-26, 4.33994e-26, 4.253751e-26, 
    4.098812e-26, 3.715069e-26, 3.411447e-26, 4.050553e-26, 3.338004e-26, 
    6.519314e-26, 4.676956e-26, 7.753115e-26, 6.716011e-26, 6.0533e-26, 
    6.338405e-26, 4.951482e-26, 4.657198e-26, 3.580937e-26, 4.113907e-26, 
    1.601136e-26, 2.524882e-26, 5.626279e-27, 9.319528e-27, 7.741438e-26, 
    7.203711e-26, 5.528679e-26, 6.28859e-26, 4.283587e-26, 3.866034e-26, 
    3.547255e-26, 3.165648e-26, 3.126191e-26, 2.915208e-26, 3.266063e-26, 
    2.928591e-26, 4.338135e-26, 3.662983e-26, 5.705364e-26, 5.152155e-26, 
    5.401993e-26, 5.685159e-26, 4.841886e-26, 4.039907e-26, 4.023917e-26, 
    3.787463e-26, 3.17087e-26, 4.276485e-26, 1.50117e-26, 2.990993e-26, 
    6.64672e-26, 5.734807e-26, 5.611999e-26, 5.949631e-26, 3.906617e-26, 
    4.581299e-26, 2.920247e-26, 3.32112e-26, 2.681804e-26, 2.988237e-26, 
    3.035172e-26, 3.465768e-26, 3.753188e-26, 4.548765e-26, 5.273304e-26, 
    5.899857e-26, 5.749962e-26, 5.07618e-26, 3.993972e-26, 3.122593e-26, 
    3.301437e-26, 2.727265e-26, 4.412043e-26, 3.640282e-26, 3.926902e-26, 
    3.209167e-26, 4.911947e-26, 3.431888e-26, 5.34847e-26, 5.157429e-26, 
    4.595422e-26, 3.591388e-26, 3.391104e-26, 3.185392e-26, 3.311342e-26, 
    3.968731e-26, 4.08409e-26, 4.6086e-26, 4.760872e-26, 5.198637e-26, 
    5.580724e-26, 5.230882e-26, 4.879572e-26, 3.968479e-26, 3.250944e-26, 
    2.572559e-26, 2.422167e-26, 1.782982e-26, 2.293425e-26, 1.494658e-26, 
    2.15921e-26, 1.104787e-26, 3.356781e-26, 2.181354e-26, 4.570907e-26, 
    4.256139e-26, 3.723921e-26, 2.673785e-26, 3.212321e-26, 2.588901e-26, 
    4.088662e-26, 5.053867e-26, 5.326344e-26, 5.860389e-26, 5.314532e-26, 
    5.357605e-26, 4.865454e-26, 5.020168e-26, 3.94035e-26, 4.498737e-26, 
    3.036335e-26, 2.593501e-26, 1.576527e-26, 1.106397e-26, 7.326945e-27, 
    5.981358e-27, 5.606326e-27, 5.454163e-27,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.004725856, 0.004725883, 0.00472588, 0.004725895, 0.004725889, 
    0.004725897, 0.004725865, 0.004725881, 0.004725873, 0.004725862, 
    0.004725908, 0.004725896, 0.004725928, 0.004725928, 0.004725925, 
    0.004725925, 0.004725925, 0.004725931, 0.004725923, 0.004725927, 
    0.004712287, 0.004725921, 0.004712235, 0.004712311, 0.004712296, 
    0.004725921, 0.004725905, 0.004725905, 0.004725903, 0.004725904, 
    0.004725905, 0.004725887, 0.004725873, 0.004725858, 0.004725862, 
    0.004725875, 0.004725904, 0.004725899, 0.004725921, 0.004725921, 
    0.004725931, 0.004725927, 0.004725933, 0.004725935, 0.004725927, 
    0.004725929, 0.004725926, 0.004725927, 0.004725926, 0.00472593, 
    0.004725928, 0.004725933, 0.004725927, 0.00472593, 0.004725909, 
    0.004725877, 0.004725864, 0.004725849, 0.004725852, 0.004725854, 
    0.004725875, 0.004725896, 0.004725908, 0.004725914, 0.00472592, 
    0.004725919, 0.004725927, 0.004725929, 0.004725934, 0.004725929, 
    0.00472593, 0.004725923, 0.004725925, 0.004725921, 0.004725933, 
    0.004725924, 0.004725936, 0.004725933, 0.004725903, 0.004725901, 
    0.004725883, 0.00472588, 0.004725853, 0.004725871, 0.004725864, 
    0.004725884, 0.004725893, 0.004725889, 0.004725914, 0.004725905, 
    0.004725928, 0.004725924, 0.00472593, 0.004725934, 0.004725929, 
    0.004725933, 0.004725925, 0.004725932, 0.004725921, 0.004712364, 
    0.004725918, 0.00471231, 0.004725932, 0.004725924, 0.004725888, 
    0.004725889, 0.004725893, 0.004725873, 0.004725873, 0.004725857, 
    0.004725873, 0.004725877, 0.004725895, 0.004725901, 0.004725907, 
    0.004725919, 0.004725925, 0.004725931, 0.004725933, 0.004725932, 
    0.004725934, 0.004725932, 0.004725934, 0.004725935, 0.004712381, 
    0.004725927, 0.004712319, 0.004712328, 0.00472592, 0.004712327, 
    0.004725889, 0.004725886, 0.004725866, 0.004725882, 0.004725855, 
    0.004725868, 0.004725874, 0.004725901, 0.00472591, 0.004725913, 
    0.004725921, 0.004725928, 0.004725931, 0.004725932, 0.004725931, 
    0.004725931, 0.004725931, 0.004725928, 0.004725932, 0.004725928, 
    0.004725925, 0.004725929, 0.004712329, 0.004712381, 0.004712328, 
    0.004712358, 0.004725887, 0.004725894, 0.00472589, 0.004725896, 
    0.004725891, 0.004725907, 0.004725911, 0.004725926, 0.004725927, 
    0.00472593, 0.004725929, 0.004725928, 0.004725922, 0.00472593, 
    0.004725928, 0.004725925, 0.004725928, 0.004725924, 0.004725928, 
    0.004725931, 0.004725927, 0.004725922, 0.004712363, 0.004712279, 
    0.004712296, 0.004712243, 0.004725904, 0.004725909, 0.004725912, 
    0.004725918, 0.004725921, 0.00472593, 0.004725933, 0.004725934, 
    0.004725935, 0.004725934, 0.004725934, 0.004725932, 0.004725914, 
    0.004725916, 0.004725917, 0.004725902, 0.004725929, 0.004725919, 
    0.004725933, 0.004725934, 0.004725922, 0.004725927, 0.004712305, 
    0.00471223, 0.004712182, 0.004712114, 0.004725915, 0.004725912, 
    0.00472592, 0.004725922, 0.004725931, 0.004725934, 0.004725935, 
    0.004725934, 0.004725935, 0.004725933, 0.00472593, 0.004725933, 
    0.004725909, 0.004725931, 0.004725907, 0.004725914, 0.004725924, 
    0.004725923, 0.004725935, 0.004725935, 0.00472593, 0.004725935, 
    0.004712245, 0.004725915, 0.004712072, 0.004712144, 0.00472591, 
    0.004725916, 0.004725927, 0.004725924, 0.004725935, 0.004725934, 
    0.004725934, 0.004725928, 0.00472593, 0.004725927, 0.004725932, 
    0.004725928, 0.004725934, 0.004725934, 0.004725931, 0.004725932, 
    0.004725933, 0.004725931, 0.004725935, 0.004725929, 0.004725935, 
    0.004725932, 0.00472591, 0.004725935, 0.004712222, 0.00472591, 
    0.004725922, 0.004725923, 0.00472593, 0.004725929, 0.004725934, 
    0.004725934, 0.004725927, 0.004725932, 0.004725925, 0.004725928, 
    0.004725929, 0.004725933, 0.004725934, 0.004725933, 0.004725931, 
    0.00472593, 0.004725931, 0.004725931, 0.00472593, 0.004725928, 
    0.004725928, 0.004725926, 0.004725935, 0.004725931, 0.004725931, 
    0.00472593, 0.004725933, 0.004725915, 0.004725933, 0.004725934, 
    0.004725934, 0.004725927, 0.004725933, 0.004725928, 0.004725932, 
    0.004725931, 0.004725934, 0.004725935, 0.004725933, 0.004725934, 
    0.004725932, 0.004725933, 0.004725931, 0.004725934, 0.004725929, 
    0.004725921, 0.004725921, 0.00471227, 0.00471236, 0.00471222, 
    0.004712324, 0.004712166, 0.004725921, 0.004712335, 0.004725935, 
    0.004725936, 0.004725928, 0.004725917, 0.00472593, 0.004725917, 
    0.004725934, 0.004725928, 0.004725933, 0.004725929, 0.004725933, 
    0.004725933, 0.004725935, 0.004725935, 0.004725934, 0.004725935, 
    0.004725927, 0.004725919, 0.004712247, 0.004712174, 0.004712112, 
    0.004712082, 0.004712074, 0.00471207,
  9.42269e-06, 9.431394e-06, 9.429709e-06, 9.436701e-06, 9.432834e-06, 
    9.437402e-06, 9.424468e-06, 9.431728e-06, 9.427102e-06, 9.42349e-06, 
    9.450187e-06, 9.437015e-06, 9.465286e-06, 9.455782e-06, 9.479638e-06, 
    9.463793e-06, 9.482828e-06, 9.479209e-06, 9.490155e-06, 9.487025e-06, 
    9.461159e-06, 9.491599e-06, 9.468216e-06, 9.459006e-06, 9.460434e-06, 
    9.491287e-06, 9.439696e-06, 9.448543e-06, 9.439165e-06, 9.44043e-06, 
    9.439868e-06, 9.432905e-06, 9.429373e-06, 9.422041e-06, 9.423378e-06, 
    9.428773e-06, 9.441e-06, 9.436872e-06, 9.447314e-06, 9.44708e-06, 
    9.459299e-06, 9.453435e-06, 9.47539e-06, 9.469158e-06, 9.487157e-06, 
    9.482636e-06, 9.486939e-06, 9.485639e-06, 9.486957e-06, 9.480324e-06, 
    9.483167e-06, 9.477333e-06, 9.454489e-06, 9.461211e-06, 9.442616e-06, 
    9.431873e-06, 9.424782e-06, 9.41972e-06, 9.420436e-06, 9.421796e-06, 
    9.428803e-06, 9.4354e-06, 9.44041e-06, 9.443752e-06, 9.447045e-06, 
    9.45735e-06, 9.46333e-06, 9.476636e-06, 9.474261e-06, 9.4783e-06, 
    9.482186e-06, 9.488669e-06, 9.487607e-06, 9.490454e-06, 9.47821e-06, 
    9.486344e-06, 9.472903e-06, 9.476582e-06, 9.44785e-06, 9.43799e-06, 
    9.433712e-06, 9.430029e-06, 9.420984e-06, 9.427229e-06, 9.424767e-06, 
    9.430641e-06, 9.434353e-06, 9.432521e-06, 9.443844e-06, 9.439444e-06, 
    9.463683e-06, 9.452596e-06, 9.481733e-06, 9.47475e-06, 9.483409e-06, 
    9.478998e-06, 9.486544e-06, 9.479753e-06, 9.49152e-06, 9.454519e-06, 
    9.492324e-06, 9.459318e-06, 9.479374e-06, 9.48693e-06, 9.432466e-06, 
    9.432764e-06, 9.434164e-06, 9.428003e-06, 9.427631e-06, 9.422e-06, 
    9.427019e-06, 9.429146e-06, 9.434576e-06, 9.437766e-06, 9.440801e-06, 
    9.447464e-06, 9.455021e-06, 9.466772e-06, 9.475202e-06, 9.480837e-06, 
    9.47739e-06, 9.480433e-06, 9.477027e-06, 9.475433e-06, 9.453612e-06, 
    9.483187e-06, 9.458381e-06, 9.457587e-06, 9.490518e-06, 9.457676e-06, 
    9.432975e-06, 9.431255e-06, 9.425246e-06, 9.429949e-06, 9.421387e-06, 
    9.426172e-06, 9.428913e-06, 9.439516e-06, 9.441862e-06, 9.444007e-06, 
    9.448262e-06, 9.453702e-06, 9.464486e-06, 9.473865e-06, 9.482416e-06, 
    9.481792e-06, 9.482011e-06, 9.483909e-06, 9.479193e-06, 9.484684e-06, 
    9.485595e-06, 9.483197e-06, 9.45748e-06, 9.453664e-06, 9.45757e-06, 
    9.455075e-06, 9.431817e-06, 9.434713e-06, 9.433147e-06, 9.436088e-06, 
    9.434009e-06, 9.443214e-06, 9.445967e-06, 9.459529e-06, 9.45359e-06, 
    9.463079e-06, 9.454538e-06, 9.456047e-06, 9.46335e-06, 9.455006e-06, 
    9.47333e-06, 9.460883e-06, 9.483983e-06, 9.471557e-06, 9.484757e-06, 
    9.482379e-06, 9.486325e-06, 9.489846e-06, 9.454725e-06, 9.462626e-06, 
    9.46079e-06, 9.467449e-06, 9.439036e-06, 9.442776e-06, 9.442464e-06, 
    9.446385e-06, 9.449278e-06, 9.455796e-06, 9.467176e-06, 9.462907e-06, 
    9.470759e-06, 9.472326e-06, 9.460407e-06, 9.467714e-06, 9.44529e-06, 
    9.448638e-06, 9.446657e-06, 9.439322e-06, 9.463867e-06, 9.4507e-06, 
    9.475339e-06, 9.468017e-06, 9.489341e-06, 9.478737e-06, 9.459778e-06, 
    9.468371e-06, 9.476542e-06, 9.486003e-06, 9.444834e-06, 9.442293e-06, 
    9.446856e-06, 9.453127e-06, 9.45968e-06, 9.468461e-06, 9.469368e-06, 
    9.471004e-06, 9.475261e-06, 9.478828e-06, 9.471505e-06, 9.479723e-06, 
    9.44938e-06, 9.465052e-06, 9.441316e-06, 9.448056e-06, 9.452765e-06, 
    9.450717e-06, 9.462423e-06, 9.465268e-06, 9.476793e-06, 9.47085e-06, 
    9.466235e-06, 9.490564e-06, 9.493251e-06, 9.481454e-06, 9.4414e-06, 
    9.444833e-06, 9.45712e-06, 9.451075e-06, 9.469056e-06, 9.473548e-06, 
    9.47721e-06, 9.481858e-06, 9.482373e-06, 9.485125e-06, 9.480611e-06, 
    9.484953e-06, 9.468479e-06, 9.475854e-06, 9.455601e-06, 9.460531e-06, 
    9.45827e-06, 9.455774e-06, 9.463468e-06, 9.471616e-06, 9.471818e-06, 
    9.474421e-06, 9.481695e-06, 9.46913e-06, 9.46815e-06, 9.484032e-06, 
    9.448569e-06, 9.455306e-06, 9.456402e-06, 9.45355e-06, 9.473097e-06, 
    9.466012e-06, 9.485061e-06, 9.479931e-06, 9.488341e-06, 9.484162e-06, 
    9.483545e-06, 9.478175e-06, 9.47482e-06, 9.466332e-06, 9.459417e-06, 
    9.453938e-06, 9.455215e-06, 9.461232e-06, 9.47212e-06, 9.482406e-06, 
    9.480152e-06, 9.487702e-06, 9.467727e-06, 9.476104e-06, 9.47286e-06, 
    9.481318e-06, 9.462788e-06, 9.478489e-06, 9.458751e-06, 9.460493e-06, 
    9.465872e-06, 9.476653e-06, 9.479075e-06, 9.481608e-06, 9.480051e-06, 
    9.472401e-06, 9.471159e-06, 9.465748e-06, 9.464238e-06, 9.460116e-06, 
    9.456686e-06, 9.459813e-06, 9.463088e-06, 9.472416e-06, 9.480784e-06, 
    9.489891e-06, 9.492127e-06, 9.462849e-06, 9.454512e-06, 9.468276e-06, 
    9.456508e-06, 9.476938e-06, 9.479437e-06, 9.456207e-06, 9.466125e-06, 
    9.469344e-06, 9.475128e-06, 9.488414e-06, 9.481278e-06, 9.489636e-06, 
    9.471112e-06, 9.461425e-06, 9.458949e-06, 9.454267e-06, 9.459056e-06, 
    9.458668e-06, 9.463243e-06, 9.461775e-06, 9.472726e-06, 9.466849e-06, 
    9.483522e-06, 9.489577e-06, 9.466741e-06, 9.476943e-06, 9.487362e-06, 
    9.491943e-06, 9.493339e-06, 9.493921e-06,
  1.94896e-10, 1.951702e-10, 1.951171e-10, 1.953381e-10, 1.952158e-10, 
    1.953603e-10, 1.949519e-10, 1.951808e-10, 1.950349e-10, 1.949212e-10, 
    1.957668e-10, 1.95348e-10, 1.962441e-10, 1.959445e-10, 1.966989e-10, 
    1.961969e-10, 1.968003e-10, 1.966852e-10, 1.970339e-10, 1.96934e-10, 
    1.965435e-10, 1.9708e-10, 1.967717e-10, 1.964739e-10, 1.9652e-10, 
    1.9707e-10, 1.95433e-10, 1.957144e-10, 1.954162e-10, 1.954563e-10, 
    1.954385e-10, 1.95218e-10, 1.951065e-10, 1.948757e-10, 1.949177e-10, 
    1.950875e-10, 1.954744e-10, 1.953435e-10, 1.956752e-10, 1.956677e-10, 
    1.960552e-10, 1.958705e-10, 1.965639e-10, 1.963665e-10, 1.969382e-10, 
    1.967942e-10, 1.969313e-10, 1.968898e-10, 1.969318e-10, 1.967207e-10, 
    1.968111e-10, 1.966256e-10, 1.959038e-10, 1.961155e-10, 1.955257e-10, 
    1.951854e-10, 1.949618e-10, 1.948028e-10, 1.948253e-10, 1.948679e-10, 
    1.950885e-10, 1.952969e-10, 1.954557e-10, 1.955618e-10, 1.956666e-10, 
    1.959938e-10, 1.961823e-10, 1.966035e-10, 1.965281e-10, 1.966563e-10, 
    1.967799e-10, 1.969865e-10, 1.969526e-10, 1.970434e-10, 1.966535e-10, 
    1.969123e-10, 1.964851e-10, 1.966018e-10, 1.956923e-10, 1.953789e-10, 
    1.952435e-10, 1.951272e-10, 1.948425e-10, 1.950389e-10, 1.949614e-10, 
    1.951465e-10, 1.952638e-10, 1.952059e-10, 1.955647e-10, 1.95425e-10, 
    1.961935e-10, 1.958437e-10, 1.967655e-10, 1.965437e-10, 1.968188e-10, 
    1.966785e-10, 1.969187e-10, 1.967025e-10, 1.970775e-10, 1.963286e-10, 
    1.971032e-10, 1.96484e-10, 1.966905e-10, 1.96931e-10, 1.952041e-10, 
    1.952135e-10, 1.952578e-10, 1.950633e-10, 1.950515e-10, 1.948744e-10, 
    1.950323e-10, 1.950993e-10, 1.952708e-10, 1.953718e-10, 1.954681e-10, 
    1.9568e-10, 1.959205e-10, 1.96291e-10, 1.96558e-10, 1.96737e-10, 
    1.966274e-10, 1.967241e-10, 1.966159e-10, 1.965653e-10, 1.962991e-10, 
    1.968117e-10, 1.964537e-10, 1.96428e-10, 1.970455e-10, 1.964309e-10, 
    1.952202e-10, 1.951659e-10, 1.949764e-10, 1.951247e-10, 1.948551e-10, 
    1.950056e-10, 1.95092e-10, 1.954273e-10, 1.955018e-10, 1.955699e-10, 
    1.957054e-10, 1.95879e-10, 1.962188e-10, 1.965156e-10, 1.967872e-10, 
    1.967673e-10, 1.967743e-10, 1.968347e-10, 1.966847e-10, 1.968594e-10, 
    1.968884e-10, 1.968121e-10, 1.964246e-10, 1.963009e-10, 1.964275e-10, 
    1.963467e-10, 1.951836e-10, 1.952752e-10, 1.952256e-10, 1.953187e-10, 
    1.952529e-10, 1.955447e-10, 1.956323e-10, 1.960625e-10, 1.958754e-10, 
    1.961744e-10, 1.959053e-10, 1.959528e-10, 1.96183e-10, 1.9592e-10, 
    1.964986e-10, 1.961051e-10, 1.968371e-10, 1.964425e-10, 1.968617e-10, 
    1.96786e-10, 1.969117e-10, 1.97024e-10, 1.963353e-10, 1.965909e-10, 
    1.965316e-10, 1.967469e-10, 1.954121e-10, 1.955308e-10, 1.955209e-10, 
    1.956456e-10, 1.957378e-10, 1.959449e-10, 1.963038e-10, 1.96169e-10, 
    1.964171e-10, 1.964668e-10, 1.960901e-10, 1.963208e-10, 1.956107e-10, 
    1.957174e-10, 1.956543e-10, 1.954211e-10, 1.961993e-10, 1.957831e-10, 
    1.965623e-10, 1.963304e-10, 1.970079e-10, 1.966702e-10, 1.964989e-10, 
    1.967767e-10, 1.970415e-10, 1.973491e-10, 1.955962e-10, 1.955154e-10, 
    1.956606e-10, 1.958606e-10, 1.960672e-10, 1.963444e-10, 1.963731e-10, 
    1.964249e-10, 1.965599e-10, 1.966731e-10, 1.964408e-10, 1.967015e-10, 
    1.95741e-10, 1.962367e-10, 1.954844e-10, 1.956988e-10, 1.958491e-10, 
    1.957837e-10, 1.961537e-10, 1.962435e-10, 1.966085e-10, 1.9642e-10, 
    1.967076e-10, 1.97047e-10, 1.975855e-10, 1.972011e-10, 1.954871e-10, 
    1.955962e-10, 1.959866e-10, 1.957951e-10, 1.963632e-10, 1.965055e-10, 
    1.966217e-10, 1.967694e-10, 1.967858e-10, 1.968734e-10, 1.967298e-10, 
    1.96868e-10, 1.96345e-10, 1.965787e-10, 1.959388e-10, 1.96094e-10, 
    1.960228e-10, 1.959442e-10, 1.961867e-10, 1.964443e-10, 1.964507e-10, 
    1.965332e-10, 1.967643e-10, 1.963656e-10, 1.967696e-10, 1.968387e-10, 
    1.957152e-10, 1.959295e-10, 1.95964e-10, 1.958742e-10, 1.964912e-10, 
    1.96267e-10, 1.968714e-10, 1.967081e-10, 1.96976e-10, 1.968428e-10, 
    1.968231e-10, 1.966524e-10, 1.965458e-10, 1.962771e-10, 1.960589e-10, 
    1.958865e-10, 1.959266e-10, 1.961161e-10, 1.964603e-10, 1.967869e-10, 
    1.967152e-10, 1.969556e-10, 1.963212e-10, 1.965866e-10, 1.964837e-10, 
    1.967522e-10, 1.961652e-10, 1.966624e-10, 1.960379e-10, 1.960928e-10, 
    1.962626e-10, 1.96604e-10, 1.966809e-10, 1.967615e-10, 1.96712e-10, 
    1.964692e-10, 1.964298e-10, 1.962586e-10, 1.96211e-10, 1.960809e-10, 
    1.959729e-10, 1.960714e-10, 1.961747e-10, 1.964696e-10, 1.967353e-10, 
    1.970255e-10, 1.970969e-10, 1.965981e-10, 1.963283e-10, 1.967736e-10, 
    1.963929e-10, 1.970544e-10, 1.966925e-10, 1.963833e-10, 1.962706e-10, 
    1.963724e-10, 1.965556e-10, 1.969784e-10, 1.96751e-10, 1.970173e-10, 
    1.964283e-10, 1.961222e-10, 1.960442e-10, 1.958968e-10, 1.960475e-10, 
    1.960353e-10, 1.961796e-10, 1.961332e-10, 1.964795e-10, 1.962935e-10, 
    1.968224e-10, 1.970154e-10, 1.96724e-10, 1.970546e-10, 1.973934e-10, 
    1.975428e-10, 1.975883e-10, 1.976073e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  2.450342, 2.427233, 2.431731, 2.413054, 2.423421, 2.411183, 2.445663, 
    2.426313, 2.438672, 2.448266, 2.376692, 2.412221, 2.339646, 2.362414, 
    2.305115, 2.343192, 2.29742, 2.306219, 2.279717, 2.287317, 2.253425, 
    2.276208, 2.235767, 2.258894, 2.255279, 2.276961, 2.405085, 2.381123, 
    2.406502, 2.40309, 2.404621, 2.423206, 2.432554, 2.452108, 2.448562, 
    2.4342, 2.401555, 2.412652, 2.384662, 2.385296, 2.354031, 2.368141, 
    2.315432, 2.330445, 2.287, 2.297944, 2.287514, 2.290678, 2.287473, 
    2.303519, 2.296647, 2.310755, 2.3655, 2.349444, 2.397243, 2.425857, 
    2.444815, 2.458241, 2.456344, 2.452727, 2.434115, 2.416582, 2.403196, 
    2.39423, 2.385386, 2.358558, 2.344332, 2.312392, 2.318167, 2.308384, 
    2.299032, 2.283308, 2.285898, 2.278963, 2.308644, 2.288928, 2.321454, 
    2.312568, 2.382972, 2.40966, 2.420971, 2.430866, 2.454885, 2.438305, 
    2.444845, 2.42928, 2.419374, 2.424275, 2.393984, 2.405773, 2.343488, 
    2.37037, 2.300124, 2.316982, 2.296079, 2.306751, 2.288456, 2.304924, 
    2.276382, 2.270246, 2.27441, 2.258146, 2.305835, 2.287513, 2.424412, 
    2.423612, 2.419889, 2.436244, 2.437244, 2.452204, 2.438895, 2.433219, 
    2.4188, 2.410257, 2.40213, 2.384233, 2.364202, 2.336118, 2.31589, 
    2.302306, 2.310639, 2.303282, 2.311505, 2.315357, 2.272579, 2.296582, 
    2.2605, 2.262506, 2.278798, 2.26228, 2.423051, 2.427649, 2.443592, 
    2.431118, 2.453832, 2.441124, 2.433808, 2.405525, 2.3993, 2.393522, 
    2.3821, 2.367419, 2.341607, 2.31909, 2.298489, 2.3, 2.299468, 2.294859, 
    2.30627, 2.292984, 2.290752, 2.296586, 2.262774, 2.272472, 2.262548, 
    2.268864, 2.426155, 2.418416, 2.422599, 2.414731, 2.420274, 2.395598, 
    2.388186, 2.353423, 2.367708, 2.344965, 2.365401, 2.361783, 2.344218, 
    2.364299, 2.320332, 2.35016, 2.29468, 2.324545, 2.292805, 2.298578, 
    2.289019, 2.280448, 2.269748, 2.249802, 2.254425, 2.237722, 2.406866, 
    2.396803, 2.397691, 2.387151, 2.379346, 2.36241, 2.335177, 2.345428, 
    2.326602, 2.322818, 2.351416, 2.333866, 2.390064, 2.381006, 2.386401, 
    2.406072, 2.343065, 2.375455, 2.315555, 2.333169, 2.28167, 2.307315, 
    2.256968, 2.235321, 2.214913, 2.191003, 2.391308, 2.398151, 2.385897, 
    2.368911, 2.353126, 2.332096, 2.329942, 2.325996, 2.315767, 2.307158, 
    2.324746, 2.304999, 2.378901, 2.340248, 2.400735, 2.382562, 2.369914, 
    2.375466, 2.346599, 2.339782, 2.312025, 2.326385, 2.240667, 2.278635, 
    2.172766, 2.202488, 2.40054, 2.391333, 2.35921, 2.374508, 2.330691, 
    2.319873, 2.31107, 2.299803, 2.298587, 2.291904, 2.302852, 2.292338, 
    2.332051, 2.314325, 2.362889, 2.351092, 2.356521, 2.362472, 2.344093, 
    2.324469, 2.324052, 2.31775, 2.299963, 2.330513, 2.235739, 2.294341, 
    2.381281, 2.363495, 2.360955, 2.36785, 2.320958, 2.337976, 2.292068, 
    2.304498, 2.284123, 2.294253, 2.295742, 2.308735, 2.316814, 2.337196, 
    2.353746, 2.366851, 2.363806, 2.349405, 2.323268, 2.298476, 2.303912, 
    2.285673, 2.333875, 2.313692, 2.321497, 2.301132, 2.3457, 2.307753, 
    2.355373, 2.351208, 2.338313, 2.31232, 2.306563, 2.300408, 2.304207, 
    2.322604, 2.325616, 2.338628, 2.342216, 2.352115, 2.360301, 2.352822, 
    2.344959, 2.322597, 2.302397, 2.280326, 2.274918, 2.249134, 2.270199, 
    2.23541, 2.264989, 2.213734, 2.305554, 2.265863, 2.337727, 2.330002, 
    2.316011, 2.283848, 2.301228, 2.2809, 2.325734, 2.348907, 2.354896, 
    2.366054, 2.35464, 2.355569, 2.344635, 2.34815, 2.321854, 2.335989, 
    2.295779, 2.281062, 2.239473, 2.213833, 2.187672, 2.1761, 2.172575, 
    2.171101,
  1.699012, 1.675992, 1.68047, 1.661885, 1.672198, 1.660024, 1.694349, 
    1.675076, 1.687382, 1.696943, 1.625765, 1.661056, 1.589066, 1.611612, 
    1.554947, 1.592574, 1.547356, 1.556037, 1.529911, 1.537398, 1.503955, 
    1.526456, 1.486617, 1.509331, 1.505777, 1.527197, 1.653962, 1.630161, 
    1.655371, 1.651979, 1.653502, 1.671984, 1.681289, 1.700773, 1.697238, 
    1.682928, 1.650453, 1.661485, 1.633678, 1.634306, 1.603307, 1.617289, 
    1.565133, 1.579967, 1.537086, 1.547874, 1.537592, 1.54071, 1.537551, 
    1.553373, 1.546595, 1.560515, 1.61467, 1.598764, 1.64617, 1.67462, 
    1.693503, 1.706888, 1.704996, 1.701389, 1.682844, 1.665395, 1.652085, 
    1.643177, 1.634397, 1.607789, 1.593703, 1.56213, 1.567834, 1.558174, 
    1.548947, 1.533447, 1.536, 1.529168, 1.558431, 1.538984, 1.571081, 
    1.562305, 1.631996, 1.65851, 1.669759, 1.679609, 1.703542, 1.687017, 
    1.693533, 1.67803, 1.668171, 1.673048, 1.642933, 1.654646, 1.592867, 
    1.619498, 1.550024, 1.566664, 1.546035, 1.556563, 1.53852, 1.554759, 
    1.526627, 1.520496, 1.524686, 1.508597, 1.555659, 1.537591, 1.673185, 
    1.672389, 1.668684, 1.684964, 1.68596, 1.700869, 1.687605, 1.681952, 
    1.667601, 1.659104, 1.651025, 1.633252, 1.613383, 1.585577, 1.565585, 
    1.552177, 1.5604, 1.55314, 1.561255, 1.565059, 1.522792, 1.546531, 
    1.510911, 1.512883, 1.529006, 1.512661, 1.671831, 1.676407, 1.692284, 
    1.67986, 1.702492, 1.689826, 1.682538, 1.654399, 1.648214, 1.642474, 
    1.631135, 1.616573, 1.591007, 1.568745, 1.548411, 1.549902, 1.549377, 
    1.544831, 1.556088, 1.542983, 1.540782, 1.546535, 1.513147, 1.522688, 
    1.512925, 1.519138, 1.67492, 1.667219, 1.67138, 1.663553, 1.669067, 
    1.644535, 1.637174, 1.602703, 1.616859, 1.59433, 1.614573, 1.610986, 
    1.593589, 1.61348, 1.569971, 1.599471, 1.544655, 1.574133, 1.542806, 
    1.548499, 1.539075, 1.530631, 1.520007, 1.500396, 1.504938, 1.488536, 
    1.655733, 1.645733, 1.646616, 1.636147, 1.628402, 1.611608, 1.584646, 
    1.594789, 1.576169, 1.572428, 1.600717, 1.583349, 1.639039, 1.630048, 
    1.635404, 1.654943, 1.592449, 1.62454, 1.565254, 1.582661, 1.531834, 
    1.557118, 1.507438, 1.486179, 1.466176, 1.442783, 1.640276, 1.647073, 
    1.634903, 1.61805, 1.60241, 1.581599, 1.579471, 1.575569, 1.565464, 
    1.556964, 1.574333, 1.554833, 1.627957, 1.589662, 1.649639, 1.631592, 
    1.619045, 1.624552, 1.595949, 1.589202, 1.561767, 1.575954, 1.491424, 
    1.528844, 1.424978, 1.454013, 1.649446, 1.6403, 1.608436, 1.623603, 
    1.580211, 1.569518, 1.560826, 1.549707, 1.548508, 1.541918, 1.552716, 
    1.542346, 1.581555, 1.564039, 1.612083, 1.600396, 1.605774, 1.61167, 
    1.593468, 1.574059, 1.573648, 1.567421, 1.549861, 1.580035, 1.486586, 
    1.544317, 1.630322, 1.612682, 1.610166, 1.617, 1.57059, 1.587415, 
    1.54208, 1.554339, 1.534251, 1.544234, 1.545702, 1.558521, 1.566498, 
    1.586643, 1.603025, 1.61601, 1.612991, 1.598726, 1.572872, 1.548398, 
    1.55376, 1.535778, 1.583359, 1.563414, 1.571123, 1.551018, 1.595058, 
    1.557548, 1.604636, 1.600512, 1.587749, 1.562058, 1.556377, 1.550303, 
    1.554052, 1.572216, 1.575193, 1.58806, 1.59161, 1.60141, 1.609519, 
    1.602109, 1.594324, 1.57221, 1.552266, 1.53051, 1.525186, 1.499738, 
    1.520448, 1.486264, 1.51532, 1.465018, 1.555379, 1.516182, 1.587169, 
    1.57953, 1.565703, 1.533978, 1.551113, 1.531075, 1.57531, 1.598231, 
    1.604164, 1.61522, 1.603911, 1.604831, 1.594005, 1.597484, 1.571476, 
    1.58545, 1.545738, 1.531235, 1.490254, 1.465117, 1.43953, 1.428231, 
    1.424792, 1.423354,
  0.7766946, 0.7627776, 0.7654802, 0.7542791, 0.7604898, 0.7531599, 
    0.7738705, 0.7622251, 0.7696564, 0.7754412, 0.7326248, 0.7537803, 
    0.7107803, 0.7241812, 0.6906163, 0.7128611, 0.6861491, 0.6912581, 
    0.6759107, 0.6803001, 0.660747, 0.6738869, 0.6506647, 0.6638809, 
    0.6618087, 0.674321, 0.7495161, 0.7352519, 0.7503623, 0.7483249, 
    0.7492394, 0.7603607, 0.7659746, 0.7777615, 0.7756197, 0.7669645, 
    0.7474091, 0.7540386, 0.7373553, 0.7377313, 0.7192376, 0.7275648, 
    0.6966211, 0.7053889, 0.6801168, 0.6864539, 0.6804138, 0.6822444, 
    0.6803899, 0.6896892, 0.6857015, 0.6938971, 0.7260035, 0.716537, 
    0.744839, 0.7619504, 0.7733588, 0.7814701, 0.7803226, 0.7781352, 
    0.7669139, 0.7563912, 0.7483889, 0.7430443, 0.7377854, 0.7219047, 
    0.7135311, 0.6948498, 0.6982155, 0.6925172, 0.6870851, 0.677983, 
    0.6794797, 0.6754755, 0.6926687, 0.6812311, 0.7001337, 0.6949527, 
    0.7363496, 0.7522494, 0.7590198, 0.7649603, 0.7794402, 0.7694353, 
    0.7733765, 0.7640073, 0.7580633, 0.7610024, 0.7428982, 0.749927, 
    0.7130355, 0.7288826, 0.6877182, 0.6975246, 0.6853724, 0.6915681, 
    0.6809587, 0.6905056, 0.6739872, 0.6704009, 0.672851, 0.6634524, 
    0.6910354, 0.6804131, 0.7610844, 0.7606049, 0.7583724, 0.7681944, 
    0.7687964, 0.7778199, 0.7697906, 0.7663751, 0.7577195, 0.7526066, 
    0.7477525, 0.7371002, 0.7252363, 0.7087115, 0.696888, 0.6889852, 
    0.6938293, 0.6895522, 0.6943336, 0.6965774, 0.6717437, 0.685664, 
    0.6648025, 0.6659534, 0.6753801, 0.6658237, 0.7602683, 0.7630281, 
    0.7726212, 0.765112, 0.7788037, 0.7711337, 0.7667289, 0.7497784, 
    0.7460651, 0.7426226, 0.735834, 0.7271381, 0.7119315, 0.6987538, 
    0.6867697, 0.6876464, 0.6873376, 0.6846652, 0.691288, 0.6835793, 
    0.6822866, 0.6856665, 0.6661075, 0.6716829, 0.6659778, 0.6696069, 
    0.762131, 0.7574896, 0.7599969, 0.7552828, 0.7586028, 0.7438582, 
    0.7394478, 0.7188787, 0.7273087, 0.7139033, 0.7259454, 0.7238083, 
    0.7134638, 0.7252941, 0.6994777, 0.7169574, 0.6845614, 0.7019377, 
    0.6834754, 0.6868214, 0.6812841, 0.6763322, 0.6701149, 0.6586742, 
    0.6613199, 0.6517788, 0.7505801, 0.7445768, 0.7451063, 0.7388333, 
    0.7342001, 0.7241787, 0.7081602, 0.714176, 0.7031413, 0.7009298, 
    0.717698, 0.7073919, 0.7405649, 0.7351843, 0.738388, 0.7501054, 0.712787, 
    0.731893, 0.6966926, 0.7069842, 0.6770376, 0.6918953, 0.6627769, 
    0.6504103, 0.6388266, 0.6253446, 0.7413055, 0.7453803, 0.7380884, 
    0.7280194, 0.7187045, 0.7063553, 0.705095, 0.7027867, 0.6968166, 
    0.6918043, 0.7020559, 0.6905492, 0.7339346, 0.7111338, 0.7469206, 
    0.7361076, 0.7286127, 0.7319001, 0.7148646, 0.7108604, 0.6946357, 
    0.7030142, 0.6534564, 0.6752853, 0.6151302, 0.6318076, 0.7468047, 
    0.7413202, 0.7222897, 0.7313329, 0.7055332, 0.6992105, 0.6940804, 
    0.6875319, 0.6868266, 0.6829538, 0.6893024, 0.6832049, 0.7063291, 
    0.6959758, 0.7244618, 0.7175068, 0.7207052, 0.7242157, 0.7133918, 
    0.7018939, 0.7016509, 0.6979719, 0.6876227, 0.7054291, 0.6506468, 
    0.6843631, 0.7353481, 0.7248185, 0.7233196, 0.7273929, 0.6998438, 
    0.7098011, 0.6830485, 0.6902581, 0.6784543, 0.6843143, 0.6851771, 
    0.6927216, 0.6974267, 0.7093435, 0.7190698, 0.7268022, 0.7250029, 
    0.7165142, 0.7011923, 0.6867618, 0.6899172, 0.6793499, 0.7073976, 
    0.6956068, 0.7001585, 0.6883036, 0.7143355, 0.6921486, 0.7200283, 
    0.7175756, 0.709999, 0.6948071, 0.6914585, 0.6878828, 0.6900892, 
    0.7008047, 0.7025644, 0.7101835, 0.712289, 0.7181096, 0.7229345, 
    0.7185254, 0.7139003, 0.700801, 0.6890377, 0.6762614, 0.6731435, 
    0.6582915, 0.6703731, 0.6504596, 0.6673768, 0.6381576, 0.6908706, 
    0.6678802, 0.7096554, 0.7051302, 0.6969579, 0.6782945, 0.6883593, 
    0.6765928, 0.7026336, 0.7162206, 0.7197471, 0.7263312, 0.7195967, 
    0.7201441, 0.7137104, 0.7157767, 0.700367, 0.7086362, 0.6851982, 
    0.676686, 0.6527765, 0.6382148, 0.623475, 0.6169931, 0.6150236, 0.6142007,
  0.1898269, 0.184835, 0.185801, 0.181808, 0.1840185, 0.1814106, 0.1888104, 
    0.1846378, 0.1872969, 0.1893755, 0.174169, 0.1816309, 0.1665713, 
    0.1712191, 0.1596566, 0.1672903, 0.1581376, 0.1598752, 0.1546741, 
    0.1561559, 0.1495906, 0.1539924, 0.1462413, 0.1506367, 0.1499447, 
    0.1541386, 0.1801186, 0.1750901, 0.1804184, 0.1796969, 0.1800206, 
    0.1839725, 0.185978, 0.1902113, 0.1894398, 0.1863323, 0.1793729, 
    0.1817226, 0.1758285, 0.1759607, 0.1694996, 0.1723992, 0.1617057, 
    0.164713, 0.1560939, 0.158241, 0.1561943, 0.1568137, 0.1561863, 
    0.1593409, 0.1579856, 0.1607751, 0.1718543, 0.1685628, 0.1784647, 
    0.1845398, 0.1886264, 0.1915497, 0.1911352, 0.190346, 0.1863142, 
    0.1825587, 0.1797195, 0.1778313, 0.1759797, 0.1704267, 0.167522, 
    0.1611004, 0.1622513, 0.1603043, 0.1584554, 0.1553731, 0.1558786, 
    0.1545274, 0.160356, 0.1564708, 0.1629084, 0.1611355, 0.1754755, 
    0.1810874, 0.1834946, 0.1856151, 0.1908167, 0.1872177, 0.1886328, 
    0.1852743, 0.1831538, 0.1842013, 0.1777798, 0.1802641, 0.1673505, 
    0.1728595, 0.1586705, 0.1620148, 0.1578739, 0.1599808, 0.1563786, 
    0.1596188, 0.1540262, 0.1528206, 0.1536439, 0.1504935, 0.1597993, 
    0.1561941, 0.1842306, 0.1840596, 0.1832639, 0.1867729, 0.1869886, 
    0.1902323, 0.1873451, 0.1861213, 0.1830314, 0.1812142, 0.1794944, 
    0.1757389, 0.1715868, 0.1658574, 0.161797, 0.1591013, 0.1607519, 
    0.1592942, 0.1609241, 0.1616907, 0.1532716, 0.1579729, 0.1509447, 
    0.1513297, 0.1544953, 0.1512863, 0.1839395, 0.1849245, 0.1883613, 
    0.1856693, 0.1905871, 0.1878271, 0.1862479, 0.1802115, 0.1788977, 
    0.1776826, 0.1752942, 0.1722502, 0.1669689, 0.1624356, 0.1583482, 
    0.1586461, 0.1585412, 0.157634, 0.1598853, 0.1572659, 0.156828, 
    0.1579737, 0.1513813, 0.1532512, 0.1513379, 0.152554, 0.1846041, 
    0.1829496, 0.1838428, 0.1821646, 0.183346, 0.1781185, 0.1765644, 
    0.1693751, 0.1723098, 0.1676507, 0.171834, 0.1710892, 0.1674987, 
    0.1716069, 0.1626836, 0.1687086, 0.1575988, 0.1635273, 0.1572307, 
    0.1583658, 0.1564887, 0.1548162, 0.1527245, 0.1489, 0.1497816, 0.1466102, 
    0.1804955, 0.1783721, 0.178559, 0.1763481, 0.174721, 0.1712182, 
    0.1656674, 0.167745, 0.1639404, 0.1631813, 0.1689653, 0.1654026, 
    0.1769576, 0.1750662, 0.1761916, 0.1803274, 0.1672646, 0.1739126, 
    0.1617302, 0.1652622, 0.1550541, 0.1600923, 0.1502679, 0.1461572, 
    0.1423403, 0.1379398, 0.1772184, 0.1786558, 0.1760862, 0.1725579, 
    0.1693145, 0.1650456, 0.164612, 0.1638186, 0.1617725, 0.1600613, 
    0.1635678, 0.1596337, 0.174628, 0.1666933, 0.1792002, 0.1753904, 
    0.1727652, 0.173915, 0.1679833, 0.1665989, 0.1610273, 0.1638967, 
    0.1471663, 0.1544634, 0.1346359, 0.1400438, 0.1791591, 0.1772235, 
    0.1705606, 0.1737164, 0.1647627, 0.162592, 0.1608376, 0.1586072, 
    0.1583676, 0.157054, 0.1592092, 0.157139, 0.1650366, 0.1614851, 
    0.1713168, 0.168899, 0.1700095, 0.1712311, 0.1674737, 0.1635122, 
    0.1634287, 0.1621679, 0.1586383, 0.1647269, 0.1462356, 0.1575318, 
    0.1751237, 0.1714412, 0.170919, 0.1723391, 0.162809, 0.1662332, 0.157086, 
    0.1595345, 0.1555322, 0.157515, 0.1578077, 0.160374, 0.1619813, 
    0.1660754, 0.1694414, 0.1721329, 0.1715054, 0.1685548, 0.1632714, 
    0.1583456, 0.1594185, 0.1558347, 0.1654046, 0.161359, 0.1629169, 
    0.1588695, 0.1678002, 0.1601788, 0.1697742, 0.1689228, 0.1663015, 
    0.1610858, 0.1599434, 0.1587265, 0.159477, 0.1631384, 0.1637423, 
    0.1663652, 0.1670924, 0.1691081, 0.1707849, 0.1692524, 0.1676496, 
    0.1631372, 0.1591192, 0.1547923, 0.1537423, 0.1487727, 0.1528113, 
    0.1461736, 0.1518066, 0.1421211, 0.1597432, 0.1519751, 0.1661829, 
    0.1646241, 0.161821, 0.1554783, 0.1588885, 0.1549041, 0.163766, 
    0.1684531, 0.1696766, 0.1719686, 0.1696243, 0.1698145, 0.1675839, 
    0.1682993, 0.1629883, 0.1658314, 0.1578149, 0.1549355, 0.1469408, 
    0.1421397, 0.1373331, 0.1352364, 0.1346015, 0.1343365,
  0.01657276, 0.01593613, 0.0160587, 0.015554, 0.01583276, 0.01550405, 
    0.01644248, 0.01591114, 0.0162491, 0.01651487, 0.014603, 0.01553172, 
    0.01367639, 0.01424091, 0.0128502, 0.01376325, 0.01267092, 0.01287605, 
    0.01226515, 0.01243823, 0.01167734, 0.01218579, 0.0112951, 0.01179754, 
    0.01171798, 0.01220279, 0.01534201, 0.01471665, 0.01537956, 0.01528925, 
    0.01532975, 0.01582694, 0.01608119, 0.01662212, 0.0165231, 0.01612624, 
    0.01524875, 0.01554324, 0.01480794, 0.0148243, 0.01403121, 0.0143854, 
    0.01309331, 0.01345274, 0.01243098, 0.01268309, 0.01244273, 0.01251532, 
    0.01244179, 0.01281287, 0.01265302, 0.01298271, 0.01431863, 0.01391738, 
    0.0151354, 0.01589873, 0.01641893, 0.01679433, 0.01674094, 0.01663943, 
    0.01612393, 0.01564849, 0.01529207, 0.01505651, 0.01482665, 0.01414416, 
    0.01379127, 0.01302135, 0.01315828, 0.01292689, 0.01270835, 0.01234671, 
    0.01240578, 0.01224807, 0.012933, 0.01247512, 0.01323667, 0.01302551, 
    0.01476428, 0.01546346, 0.01576656, 0.01603508, 0.01669995, 0.016239, 
    0.01641975, 0.01599183, 0.01572352, 0.01585588, 0.0150501, 0.01536024, 
    0.01377053, 0.01444189, 0.01273372, 0.01313011, 0.01263987, 0.01288855, 
    0.01246432, 0.01284572, 0.01218972, 0.01204976, 0.01214529, 0.01178105, 
    0.01286707, 0.01244271, 0.01585959, 0.01583795, 0.01573741, 0.01618232, 
    0.0162098, 0.01662482, 0.01625524, 0.0160994, 0.01570808, 0.01547938, 
    0.01526393, 0.01479685, 0.01428589, 0.01359034, 0.01310417, 0.01278456, 
    0.01297996, 0.01280735, 0.0130004, 0.01309153, 0.01210207, 0.01265152, 
    0.011833, 0.01187739, 0.01224433, 0.01187238, 0.01582277, 0.01594746, 
    0.01638502, 0.01604196, 0.01667042, 0.01631676, 0.01611551, 0.01535366, 
    0.01518941, 0.01503801, 0.01474185, 0.01436713, 0.0137244, 0.01318026, 
    0.01269572, 0.01273084, 0.01271847, 0.01261166, 0.01287725, 0.01256839, 
    0.012517, 0.01265162, 0.01188334, 0.01209969, 0.01187833, 0.01201888, 
    0.01590687, 0.01569775, 0.01581053, 0.01559886, 0.01574778, 0.01509227, 
    0.01489913, 0.01401607, 0.01437444, 0.01380684, 0.01431614, 0.01422503, 
    0.01378846, 0.01428834, 0.01320985, 0.01393508, 0.01260752, 0.01331066, 
    0.01256426, 0.01269779, 0.01247721, 0.01228172, 0.01203863, 0.01159818, 
    0.01169925, 0.01133699, 0.01538923, 0.01512386, 0.01514716, 0.0148723, 
    0.01467105, 0.0142408, 0.01356745, 0.01381826, 0.0133601, 0.01326929, 
    0.01396625, 0.0135356, 0.01494791, 0.01471368, 0.0148529, 0.01536816, 
    0.01376014, 0.01457139, 0.01309622, 0.01351871, 0.01230947, 0.01290177, 
    0.01175511, 0.01128556, 0.01085507, 0.01036544, 0.0149803, 0.01515923, 
    0.01483984, 0.01440488, 0.0140087, 0.01349269, 0.01344061, 0.01334552, 
    0.01310126, 0.01289809, 0.0133155, 0.01284747, 0.0146596, 0.01369112, 
    0.01522717, 0.01475374, 0.01443032, 0.01457169, 0.01384712, 0.01367971, 
    0.01301266, 0.01335487, 0.01140026, 0.01224062, 0.01000258, 0.01059864, 
    0.01522204, 0.01498094, 0.01416048, 0.01454724, 0.0134587, 0.01319891, 
    0.01299013, 0.01272625, 0.01269801, 0.01254351, 0.01279731, 0.01255349, 
    0.0134916, 0.01306706, 0.01425285, 0.0139582, 0.01409328, 0.01424237, 
    0.01378542, 0.01330885, 0.01329886, 0.01314835, 0.01272994, 0.0134544, 
    0.01129447, 0.01259966, 0.01472077, 0.01426808, 0.01420424, 0.01437803, 
    0.01322481, 0.01363561, 0.01254727, 0.01283575, 0.01236529, 0.01259766, 
    0.01263208, 0.01293514, 0.01312612, 0.01361659, 0.01402413, 0.01435276, 
    0.01427592, 0.01391642, 0.01328006, 0.01269542, 0.01282204, 0.01240065, 
    0.01353583, 0.01305207, 0.0132377, 0.0127572, 0.01382494, 0.01291203, 
    0.01406463, 0.01396109, 0.01364385, 0.01301962, 0.01288413, 0.01274032, 
    0.01282895, 0.01326416, 0.01333638, 0.01365152, 0.01373932, 0.0139836, 
    0.01418786, 0.01400114, 0.01380671, 0.01326401, 0.01278668, 0.01227894, 
    0.01215671, 0.01158362, 0.0120487, 0.01128744, 0.01193246, 0.01083052, 
    0.01286045, 0.01195193, 0.01362955, 0.01344206, 0.01310703, 0.012359, 
    0.01275943, 0.01229198, 0.01333922, 0.01390408, 0.01405274, 0.01433262, 
    0.01404639, 0.01406953, 0.01379875, 0.01388541, 0.01324623, 0.0135872, 
    0.01263293, 0.01229564, 0.01137459, 0.01083259, 0.01029849, 0.01006823, 
    0.009998826, 0.009969902,
  0.0004566624, 0.0004320031, 0.0004367211, 0.0004173861, 0.0004280352, 
    0.0004154858, 0.000451585, 0.0004310432, 0.0004440784, 0.000454404, 
    0.0003816249, 0.0004165384, 0.0003476543, 0.0003682451, 0.0003181235, 
    0.000350801, 0.0003118128, 0.0003190363, 0.0002976614, 0.0003036752, 
    0.0002774913, 0.0002949153, 0.0002645903, 0.0002815835, 0.0002788731, 
    0.000295503, 0.0004093378, 0.0003858515, 0.0004107601, 0.0004073414, 
    0.0004088735, 0.0004278123, 0.0004375888, 0.0004585896, 0.0004547251, 
    0.0004393271, 0.0004058109, 0.0004169767, 0.0003892554, 0.0003898664, 
    0.000360558, 0.0003735682, 0.0003267369, 0.0003395882, 0.0003034224, 
    0.0003122402, 0.0003038321, 0.0003063644, 0.0003037992, 0.0003168064, 
    0.0003111848, 0.0003228103, 0.0003711057, 0.0003564039, 0.0004015354, 
    0.0004305669, 0.0004506692, 0.0004653326, 0.0004632392, 0.0004592665, 
    0.0004392381, 0.0004209873, 0.000407448, 0.0003985673, 0.0003899543, 
    0.0003646933, 0.0003518177, 0.0003241806, 0.0003290496, 0.0003208336, 
    0.0003131276, 0.000300491, 0.0003025452, 0.0002970698, 0.00032105, 
    0.0003049614, 0.0003318462, 0.0003243283, 0.0003876269, 0.0004139434, 
    0.0004254998, 0.000435811, 0.000461634, 0.0004436872, 0.0004507011, 
    0.0004341454, 0.0004238533, 0.0004289219, 0.0003983264, 0.0004100279, 
    0.000351065, 0.0003756552, 0.0003140194, 0.0003280461, 0.0003107235, 
    0.000319478, 0.0003045846, 0.0003179652, 0.0002950511, 0.0002902248, 
    0.0002935165, 0.0002810212, 0.000318719, 0.0003038314, 0.0004290641, 
    0.0004282342, 0.0004243844, 0.000441494, 0.000442557, 0.0004586954, 
    0.0004443162, 0.0004382911, 0.0004232629, 0.0004145479, 0.0004063841, 
    0.0003888416, 0.0003699001, 0.0003445444, 0.0003271232, 0.0003158088, 
    0.0003227129, 0.0003166118, 0.0003234374, 0.0003266734, 0.0002920259, 
    0.0003111323, 0.0002827941, 0.0002843112, 0.0002969402, 0.00028414, 
    0.0004276524, 0.0004324387, 0.000449351, 0.0004360762, 0.000460478, 
    0.0004467008, 0.0004389131, 0.0004097788, 0.0004035709, 0.0003978724, 
    0.00038679, 0.0003728941, 0.0003493922, 0.0003298331, 0.0003126838, 
    0.000313918, 0.000313483, 0.0003097345, 0.0003190788, 0.0003082198, 
    0.0003064233, 0.0003111355, 0.0002845148, 0.0002919438, 0.0002843435, 
    0.0002891628, 0.0004308789, 0.0004228685, 0.0004271835, 0.0004190948, 
    0.000424781, 0.0003999122, 0.0003926646, 0.0003600047, 0.0003731636, 
    0.0003523831, 0.0003710141, 0.0003676616, 0.000351716, 0.0003699901, 
    0.0003308888, 0.0003570493, 0.0003095895, 0.0003344919, 0.0003080751, 
    0.0003127565, 0.0003050342, 0.0002982357, 0.0002898418, 0.0002748056, 
    0.0002782358, 0.0002659957, 0.0004111266, 0.0004011009, 0.0004019783, 
    0.0003916609, 0.0003841537, 0.000368241, 0.0003437187, 0.0003527975, 
    0.0003362627, 0.0003330116, 0.0003581854, 0.0003425704, 0.0003944916, 
    0.0003857409, 0.0003909353, 0.0004103282, 0.000350688, 0.0003804515, 
    0.0003268405, 0.0003419619, 0.000299198, 0.0003199453, 0.0002801371, 
    0.0002642705, 0.000249954, 0.000233947, 0.000395706, 0.000402433, 
    0.0003904472, 0.0003742877, 0.0003597354, 0.000341025, 0.0003391521, 
    0.0003357401, 0.0003270196, 0.0003198149, 0.0003346649, 0.0003180272, 
    0.0003837281, 0.0003481873, 0.0004049959, 0.0003872336, 0.0003752274, 
    0.0003804624, 0.0003538465, 0.0003477743, 0.0003238722, 0.0003360751, 
    0.0002681226, 0.0002968119, 0.0002222784, 0.0002415337, 0.0004048022, 
    0.0003957299, 0.0003652916, 0.0003795556, 0.0003398024, 0.0003304984, 
    0.0003230734, 0.0003137569, 0.000312764, 0.0003073497, 0.0003162579, 
    0.0003076986, 0.0003409859, 0.0003258039, 0.0003686843, 0.0003578919, 
    0.0003628286, 0.0003682988, 0.0003516052, 0.0003344269, 0.0003340692, 
    0.0003286958, 0.0003138871, 0.0003396478, 0.0002645694, 0.0003093146, 
    0.0003860046, 0.0003692446, 0.0003668976, 0.0003732964, 0.0003314226, 
    0.0003461795, 0.0003074812, 0.0003176136, 0.0003011367, 0.0003092444, 
    0.0003104504, 0.0003211255, 0.0003279041, 0.0003454922, 0.0003602991, 
    0.0003723637, 0.000369533, 0.0003563689, 0.0003333968, 0.0003126731, 
    0.00031713, 0.0003023666, 0.0003425786, 0.0003252714, 0.0003318828, 
    0.0003148454, 0.0003530406, 0.0003203084, 0.00036178, 0.0003579973, 
    0.0003464772, 0.0003241193, 0.0003193216, 0.0003142516, 0.0003173736, 
    0.0003328285, 0.0003354127, 0.0003467546, 0.0003499331, 0.0003588187, 
    0.0003662962, 0.0003594592, 0.0003523783, 0.0003328229, 0.0003158835, 
    0.0002981393, 0.0002939108, 0.0002743126, 0.0002901883, 0.0002643339, 
    0.0002861974, 0.0002491447, 0.0003184855, 0.0002868644, 0.0003459603, 
    0.0003392043, 0.0003272251, 0.0003009184, 0.000314924, 0.0002985914, 
    0.0003355144, 0.0003559195, 0.0003613451, 0.0003716215, 0.0003611126, 
    0.0003619593, 0.0003520891, 0.0003552396, 0.0003321875, 0.000344431, 
    0.00031048, 0.0002987185, 0.0002672588, 0.000249213, 0.0002317813, 
    0.000224377, 0.0002221585, 0.0002212358,
  3.51061e-06, 3.237437e-06, 3.28925e-06, 3.078303e-06, 3.194029e-06, 
    3.057771e-06, 3.453889e-06, 3.226922e-06, 3.370477e-06, 3.48535e-06, 
    2.698163e-06, 3.06914e-06, 2.349834e-06, 2.559429e-06, 2.057902e-06, 
    2.381551e-06, 1.996902e-06, 2.066767e-06, 1.861957e-06, 1.918986e-06, 
    1.6742e-06, 1.836073e-06, 1.557054e-06, 1.711845e-06, 1.686885e-06, 
    1.841604e-06, 2.991595e-06, 2.742392e-06, 3.00687e-06, 2.97019e-06, 
    2.986613e-06, 3.191596e-06, 3.298804e-06, 3.532201e-06, 3.488939e-06, 
    3.317962e-06, 2.953807e-06, 3.073875e-06, 2.778147e-06, 2.784579e-06, 
    2.480618e-06, 2.614387e-06, 2.141961e-06, 2.269057e-06, 1.91658e-06, 
    2.001016e-06, 1.920481e-06, 1.94464e-06, 1.920168e-06, 2.045129e-06, 
    1.990858e-06, 2.103527e-06, 2.588924e-06, 2.438307e-06, 2.908169e-06, 
    3.221709e-06, 3.443684e-06, 3.608022e-06, 3.584438e-06, 3.539794e-06, 
    3.31698e-06, 3.117311e-06, 2.97133e-06, 2.876596e-06, 2.785504e-06, 
    2.522935e-06, 2.391823e-06, 2.116919e-06, 2.164686e-06, 2.084252e-06, 
    2.009568e-06, 1.888732e-06, 1.908235e-06, 1.856372e-06, 2.086358e-06, 
    1.931245e-06, 2.192252e-06, 2.118363e-06, 2.761027e-06, 3.041132e-06, 
    3.166376e-06, 3.279238e-06, 3.566382e-06, 3.366146e-06, 3.44404e-06, 
    3.260936e-06, 3.148449e-06, 3.203715e-06, 2.874038e-06, 2.999004e-06, 
    2.384217e-06, 2.636021e-06, 2.018173e-06, 2.154818e-06, 1.986422e-06, 
    2.071059e-06, 1.927652e-06, 2.056365e-06, 1.837351e-06, 1.792093e-06, 
    1.822927e-06, 1.706658e-06, 2.063683e-06, 1.920474e-06, 3.205269e-06, 
    3.196202e-06, 3.154227e-06, 3.341886e-06, 3.353638e-06, 3.533388e-06, 
    3.373111e-06, 3.306539e-06, 3.142027e-06, 3.04765e-06, 2.959938e-06, 
    2.773793e-06, 2.576482e-06, 2.3186e-06, 2.145753e-06, 2.035468e-06, 
    2.102576e-06, 2.043244e-06, 2.109652e-06, 2.141337e-06, 1.808946e-06, 
    1.990353e-06, 1.723025e-06, 1.737066e-06, 1.855149e-06, 1.73548e-06, 
    3.189849e-06, 3.24221e-06, 3.429009e-06, 3.282153e-06, 3.553393e-06, 
    3.399556e-06, 3.313396e-06, 2.996329e-06, 2.929872e-06, 2.869218e-06, 
    2.752235e-06, 2.60741e-06, 2.367336e-06, 2.1724e-06, 2.00529e-06, 
    2.017194e-06, 2.012996e-06, 1.976922e-06, 2.067178e-06, 1.962394e-06, 
    1.945203e-06, 1.990383e-06, 1.738952e-06, 1.808177e-06, 1.737365e-06, 
    1.782176e-06, 3.225122e-06, 3.13774e-06, 3.184731e-06, 3.096795e-06, 
    3.158545e-06, 2.890893e-06, 2.814086e-06, 2.474972e-06, 2.610199e-06, 
    2.39754e-06, 2.587978e-06, 2.553424e-06, 2.390796e-06, 2.57741e-06, 
    2.182806e-06, 2.444869e-06, 1.975529e-06, 2.218421e-06, 1.961008e-06, 
    2.005991e-06, 1.931939e-06, 1.867382e-06, 1.788514e-06, 1.649619e-06, 
    1.681031e-06, 1.5697e-06, 3.010809e-06, 2.903541e-06, 2.912886e-06, 
    2.803491e-06, 2.724599e-06, 2.559386e-06, 2.310325e-06, 2.401733e-06, 
    2.235978e-06, 2.203768e-06, 2.456428e-06, 2.298833e-06, 2.833394e-06, 
    2.74123e-06, 2.79584e-06, 3.002229e-06, 2.380409e-06, 2.685916e-06, 
    2.142978e-06, 2.292748e-06, 1.876484e-06, 2.075605e-06, 1.698512e-06, 
    1.554181e-06, 1.427069e-06, 1.288627e-06, 2.846248e-06, 2.917733e-06, 
    2.790696e-06, 2.62184e-06, 2.472224e-06, 2.28339e-06, 2.264712e-06, 
    2.230792e-06, 2.144735e-06, 2.074336e-06, 2.220133e-06, 2.056967e-06, 
    2.720147e-06, 2.355197e-06, 2.945092e-06, 2.756894e-06, 2.631581e-06, 
    2.686028e-06, 2.412355e-06, 2.351039e-06, 2.113903e-06, 2.234117e-06, 
    1.588895e-06, 1.85394e-06, 1.190268e-06, 1.353748e-06, 2.943021e-06, 
    2.846501e-06, 2.52907e-06, 2.676575e-06, 2.271193e-06, 2.178955e-06, 
    2.106097e-06, 2.01564e-06, 2.006063e-06, 1.954063e-06, 2.039816e-06, 
    1.957403e-06, 2.283e-06, 2.132811e-06, 2.56395e-06, 2.45344e-06, 
    2.503828e-06, 2.559981e-06, 2.389673e-06, 2.217776e-06, 2.214233e-06, 
    2.161206e-06, 2.016899e-06, 2.269652e-06, 1.556869e-06, 1.972895e-06, 
    2.743993e-06, 2.569725e-06, 2.545566e-06, 2.611572e-06, 2.188072e-06, 
    2.335007e-06, 1.955322e-06, 2.052954e-06, 1.894856e-06, 1.972217e-06, 
    1.983797e-06, 2.087094e-06, 2.153422e-06, 2.328106e-06, 2.477976e-06, 
    2.601923e-06, 2.572696e-06, 2.437951e-06, 2.207579e-06, 2.005187e-06, 
    2.048265e-06, 1.906537e-06, 2.298915e-06, 2.127595e-06, 2.192615e-06, 
    2.026152e-06, 2.404193e-06, 2.079141e-06, 2.493102e-06, 2.454513e-06, 
    2.337997e-06, 2.11632e-06, 2.069539e-06, 2.020415e-06, 2.050626e-06, 
    2.201959e-06, 2.227546e-06, 2.340785e-06, 2.37279e-06, 2.462878e-06, 
    2.539384e-06, 2.469407e-06, 2.397491e-06, 2.201903e-06, 2.036193e-06, 
    1.866472e-06, 1.82663e-06, 1.645119e-06, 1.791753e-06, 1.554753e-06, 
    1.75457e-06, 1.419977e-06, 2.061418e-06, 1.760768e-06, 2.332805e-06, 
    2.265232e-06, 2.146754e-06, 1.892786e-06, 2.026912e-06, 1.870746e-06, 
    2.228554e-06, 2.433386e-06, 2.488657e-06, 2.594252e-06, 2.486282e-06, 
    2.494935e-06, 2.394566e-06, 2.426482e-06, 2.195623e-06, 2.317462e-06, 
    1.984082e-06, 1.871948e-06, 1.581091e-06, 1.420574e-06, 1.270204e-06, 
    1.207793e-06, 1.189268e-06, 1.181587e-06,
  4.241074e-09, 3.589786e-09, 3.710587e-09, 3.227115e-09, 3.489595e-09, 
    3.181262e-09, 4.102966e-09, 3.565431e-09, 3.902573e-09, 4.179387e-09, 
    2.415208e-09, 3.206625e-09, 1.746218e-09, 2.139585e-09, 1.248865e-09, 
    1.80389e-09, 1.153027e-09, 1.263033e-09, 9.51759e-10, 1.034968e-09, 
    6.980488e-10, 9.149106e-10, 5.565537e-10, 7.463336e-10, 7.141696e-10, 
    9.227362e-10, 3.034975e-09, 2.505498e-09, 3.068537e-09, 2.988158e-09, 
    3.024057e-09, 3.484007e-09, 3.733008e-09, 4.294027e-09, 4.188133e-09, 
    3.778091e-09, 2.95249e-09, 3.217206e-09, 2.579312e-09, 2.59267e-09, 
    1.988326e-09, 2.247364e-09, 1.385657e-09, 1.602459e-09, 1.031402e-09, 
    1.159397e-09, 1.037187e-09, 1.073289e-09, 1.036722e-09, 1.228553e-09, 
    1.143692e-09, 1.322443e-09, 2.197197e-09, 1.908764e-09, 2.853891e-09, 
    3.553381e-09, 4.078276e-09, 4.481642e-09, 4.42301e-09, 4.312701e-09, 
    3.775776e-09, 3.314826e-09, 2.990643e-09, 2.786347e-09, 2.594594e-09, 
    2.069058e-09, 1.822711e-09, 1.344343e-09, 1.423554e-09, 1.291163e-09, 
    1.172684e-09, 9.904828e-10, 1.019072e-09, 9.437605e-10, 1.294566e-09, 
    1.053213e-09, 1.470037e-09, 1.346712e-09, 2.543883e-09, 3.144262e-09, 
    3.426263e-09, 3.687143e-09, 4.378289e-09, 3.89226e-09, 4.079137e-09, 
    3.644408e-09, 3.385401e-09, 3.511869e-09, 2.780899e-09, 3.051238e-09, 
    1.808767e-09, 2.290302e-09, 1.186111e-09, 1.40705e-09, 1.136859e-09, 
    1.269915e-09, 1.047853e-09, 1.246412e-09, 9.167166e-10, 8.536455e-10, 
    8.964196e-10, 7.396008e-10, 1.258097e-09, 1.037178e-09, 3.515448e-09, 
    3.494588e-09, 3.398552e-09, 3.834638e-09, 3.862516e-09, 4.296943e-09, 
    3.908852e-09, 3.751187e-09, 3.370805e-09, 3.158739e-09, 2.96582e-09, 
    2.570284e-09, 2.17283e-09, 1.690095e-09, 1.391953e-09, 1.213276e-09, 
    1.320892e-09, 1.225565e-09, 1.332441e-09, 1.384621e-09, 8.769213e-10, 
    1.142913e-09, 7.6093e-10, 7.794247e-10, 9.420128e-10, 7.773261e-10, 
    3.479995e-09, 3.600856e-09, 4.042856e-09, 3.693962e-09, 4.346207e-09, 
    3.972066e-09, 3.76733e-09, 3.045367e-09, 2.900637e-09, 2.770643e-09, 
    2.525738e-09, 2.233579e-09, 1.777956e-09, 1.436508e-09, 1.166029e-09, 
    1.184579e-09, 1.178025e-09, 1.12228e-09, 1.263693e-09, 1.100129e-09, 
    1.074138e-09, 1.14296e-09, 7.819237e-10, 8.758517e-10, 7.79821e-10, 
    8.40066e-10, 3.561264e-09, 3.361073e-09, 3.468255e-09, 3.268597e-09, 
    3.408392e-09, 2.816866e-09, 2.654261e-09, 1.977645e-09, 2.239087e-09, 
    1.833217e-09, 2.19534e-09, 2.127921e-09, 1.820829e-09, 2.174641e-09, 
    1.454049e-09, 1.92103e-09, 1.12015e-09, 1.514684e-09, 1.098024e-09, 
    1.167118e-09, 1.054249e-09, 9.595571e-10, 8.487346e-10, 6.672433e-10, 
    7.067092e-10, 5.711711e-10, 3.07721e-09, 2.843958e-09, 2.864028e-09, 
    2.632085e-09, 2.469028e-09, 2.1395e-09, 1.675338e-09, 1.840933e-09, 
    1.544908e-09, 1.489623e-09, 1.942695e-09, 1.654925e-09, 2.694823e-09, 
    2.503104e-09, 2.616116e-09, 3.058328e-09, 1.801799e-09, 2.390404e-09, 
    1.387344e-09, 1.644151e-09, 9.726936e-10, 1.277224e-09, 7.290792e-10, 
    5.53257e-10, 4.159632e-10, 2.867027e-10, 2.721946e-09, 2.874458e-09, 
    2.605396e-09, 2.262127e-09, 1.972449e-09, 1.627635e-09, 1.594854e-09, 
    1.535957e-09, 1.390262e-09, 1.27518e-09, 1.51762e-09, 1.247371e-09, 
    2.459942e-09, 1.75592e-09, 2.933572e-09, 2.535346e-09, 2.281468e-09, 
    2.390629e-09, 1.860542e-09, 1.748394e-09, 1.3394e-09, 1.541693e-09, 
    5.936692e-10, 9.402864e-10, 2.086518e-10, 3.447674e-10, 2.929082e-09, 
    2.722479e-09, 2.080853e-09, 2.371549e-09, 1.606201e-09, 1.447547e-09, 
    1.326633e-09, 1.182152e-09, 1.16723e-09, 1.087503e-09, 1.220141e-09, 
    1.092557e-09, 1.626948e-09, 1.370507e-09, 2.14838e-09, 1.937086e-09, 
    2.03246e-09, 2.140656e-09, 1.818762e-09, 1.513575e-09, 1.507501e-09, 
    1.417727e-09, 1.184127e-09, 1.6035e-09, 5.563454e-10, 1.116129e-09, 
    2.508778e-09, 2.159637e-09, 2.112692e-09, 2.241799e-09, 1.462953e-09, 
    1.719491e-09, 1.089406e-09, 1.240979e-09, 9.994252e-10, 1.115088e-09, 
    1.132823e-09, 1.295756e-09, 1.404722e-09, 1.707104e-09, 1.983324e-09, 
    2.222757e-09, 2.165431e-09, 1.9081e-09, 1.496126e-09, 1.16587e-09, 
    1.233529e-09, 1.01657e-09, 1.655068e-09, 1.361898e-09, 1.470656e-09, 
    1.198613e-09, 1.845468e-09, 1.282922e-09, 2.012021e-09, 1.939099e-09, 
    1.724869e-09, 1.343362e-09, 1.267476e-09, 1.18962e-09, 1.237278e-09, 
    1.48654e-09, 1.530362e-09, 1.729886e-09, 1.787889e-09, 1.954824e-09, 
    2.10074e-09, 1.967131e-09, 1.833126e-09, 1.486444e-09, 1.21442e-09, 
    9.582476e-10, 9.016126e-10, 6.616702e-10, 8.531811e-10, 5.539156e-10, 
    8.027432e-10, 4.088173e-10, 1.25448e-09, 8.110609e-10, 1.715534e-09, 
    1.595763e-09, 1.393619e-09, 9.964017e-10, 1.199807e-09, 9.644052e-10, 
    1.5321e-09, 1.899588e-09, 2.003573e-09, 2.20766e-09, 1.999063e-09, 
    2.01551e-09, 1.827745e-09, 1.886735e-09, 1.475762e-09, 1.68806e-09, 
    1.133263e-09, 9.661388e-10, 5.844773e-10, 4.094148e-10, 2.711841e-10, 
    2.216841e-10, 2.079199e-10, 2.023397e-10,
  4.175727e-13, 4.150125e-13, 4.154877e-13, 4.135849e-13, 4.146183e-13, 
    4.134043e-13, 4.170302e-13, 4.149167e-13, 4.162426e-13, 4.173304e-13, 
    4.10383e-13, 4.135042e-13, 4.077376e-13, 4.09294e-13, 4.05766e-13, 
    4.07966e-13, 4.053854e-13, 4.058222e-13, 4.045855e-13, 4.049164e-13, 
    4.035756e-13, 4.04439e-13, 4.030114e-13, 4.037679e-13, 4.036398e-13, 
    4.044701e-13, 4.128279e-13, 4.107395e-13, 4.129602e-13, 4.126434e-13, 
    4.127849e-13, 4.145963e-13, 4.155759e-13, 4.177807e-13, 4.173647e-13, 
    4.157532e-13, 4.125028e-13, 4.135459e-13, 4.110309e-13, 4.110836e-13, 
    4.086958e-13, 4.0972e-13, 4.063087e-13, 4.071682e-13, 4.049022e-13, 
    4.054108e-13, 4.049252e-13, 4.050687e-13, 4.049233e-13, 4.056854e-13, 
    4.053484e-13, 4.06058e-13, 4.095217e-13, 4.08381e-13, 4.121141e-13, 
    4.148693e-13, 4.169331e-13, 4.185173e-13, 4.182871e-13, 4.17854e-13, 
    4.157441e-13, 4.139303e-13, 4.126532e-13, 4.118477e-13, 4.110912e-13, 
    4.090151e-13, 4.080405e-13, 4.061449e-13, 4.06459e-13, 4.059339e-13, 
    4.054635e-13, 4.047395e-13, 4.048532e-13, 4.045537e-13, 4.059474e-13, 
    4.049889e-13, 4.066434e-13, 4.061543e-13, 4.108911e-13, 4.132585e-13, 
    4.14369e-13, 4.153955e-13, 4.181115e-13, 4.162021e-13, 4.169365e-13, 
    4.152274e-13, 4.142082e-13, 4.147059e-13, 4.118263e-13, 4.12892e-13, 
    4.079853e-13, 4.098896e-13, 4.055168e-13, 4.063936e-13, 4.053212e-13, 
    4.058495e-13, 4.049676e-13, 4.057562e-13, 4.044461e-13, 4.041952e-13, 
    4.043654e-13, 4.037411e-13, 4.058026e-13, 4.049251e-13, 4.1472e-13, 
    4.146379e-13, 4.142599e-13, 4.159755e-13, 4.160851e-13, 4.177921e-13, 
    4.162673e-13, 4.156474e-13, 4.141507e-13, 4.133156e-13, 4.125554e-13, 
    4.109953e-13, 4.094254e-13, 4.075153e-13, 4.063337e-13, 4.056247e-13, 
    4.060518e-13, 4.056735e-13, 4.060977e-13, 4.063047e-13, 4.042878e-13, 
    4.053453e-13, 4.038261e-13, 4.038997e-13, 4.045468e-13, 4.038914e-13, 
    4.145805e-13, 4.150561e-13, 4.16794e-13, 4.154223e-13, 4.179856e-13, 
    4.165158e-13, 4.157109e-13, 4.128689e-13, 4.122984e-13, 4.117858e-13, 
    4.108194e-13, 4.096655e-13, 4.078633e-13, 4.065104e-13, 4.054371e-13, 
    4.055107e-13, 4.054847e-13, 4.052633e-13, 4.058248e-13, 4.051753e-13, 
    4.05072e-13, 4.053455e-13, 4.039097e-13, 4.042836e-13, 4.039013e-13, 
    4.041411e-13, 4.149003e-13, 4.141124e-13, 4.145343e-13, 4.137482e-13, 
    4.142987e-13, 4.119681e-13, 4.113267e-13, 4.086536e-13, 4.096873e-13, 
    4.08082e-13, 4.095144e-13, 4.092479e-13, 4.08033e-13, 4.094326e-13, 
    4.0658e-13, 4.084296e-13, 4.052548e-13, 4.068203e-13, 4.051669e-13, 
    4.054414e-13, 4.04993e-13, 4.046166e-13, 4.041756e-13, 4.034528e-13, 
    4.036101e-13, 4.030697e-13, 4.129943e-13, 4.120749e-13, 4.121541e-13, 
    4.112392e-13, 4.105955e-13, 4.092936e-13, 4.074569e-13, 4.081126e-13, 
    4.069401e-13, 4.06721e-13, 4.085153e-13, 4.07376e-13, 4.114867e-13, 
    4.107301e-13, 4.111761e-13, 4.129199e-13, 4.079577e-13, 4.102851e-13, 
    4.063154e-13, 4.073333e-13, 4.046688e-13, 4.058785e-13, 4.036992e-13, 
    4.029982e-13, 4.024501e-13, 4.019333e-13, 4.115937e-13, 4.121952e-13, 
    4.111339e-13, 4.097783e-13, 4.08633e-13, 4.072679e-13, 4.07138e-13, 
    4.069047e-13, 4.06327e-13, 4.058704e-13, 4.06832e-13, 4.057601e-13, 
    4.105597e-13, 4.07776e-13, 4.124283e-13, 4.108574e-13, 4.098547e-13, 
    4.10286e-13, 4.081902e-13, 4.077462e-13, 4.061253e-13, 4.069274e-13, 
    4.031594e-13, 4.045399e-13, 4.016209e-13, 4.021656e-13, 4.124106e-13, 
    4.115958e-13, 4.090618e-13, 4.102106e-13, 4.07183e-13, 4.065542e-13, 
    4.060746e-13, 4.055011e-13, 4.054418e-13, 4.051252e-13, 4.05652e-13, 
    4.051452e-13, 4.072652e-13, 4.062487e-13, 4.093287e-13, 4.084931e-13, 
    4.088704e-13, 4.092982e-13, 4.080248e-13, 4.068159e-13, 4.067919e-13, 
    4.06436e-13, 4.05509e-13, 4.071723e-13, 4.030106e-13, 4.052389e-13, 
    4.107525e-13, 4.093732e-13, 4.091877e-13, 4.09698e-13, 4.066153e-13, 
    4.076317e-13, 4.051327e-13, 4.057347e-13, 4.047751e-13, 4.052347e-13, 
    4.053052e-13, 4.059521e-13, 4.063844e-13, 4.075827e-13, 4.08676e-13, 
    4.096227e-13, 4.093961e-13, 4.083784e-13, 4.067468e-13, 4.054365e-13, 
    4.057051e-13, 4.048432e-13, 4.073766e-13, 4.062145e-13, 4.066458e-13, 
    4.055665e-13, 4.081305e-13, 4.059012e-13, 4.087895e-13, 4.085011e-13, 
    4.076531e-13, 4.06141e-13, 4.058399e-13, 4.055308e-13, 4.0572e-13, 
    4.067088e-13, 4.068825e-13, 4.076729e-13, 4.079026e-13, 4.085633e-13, 
    4.091404e-13, 4.08612e-13, 4.080817e-13, 4.067084e-13, 4.056293e-13, 
    4.046113e-13, 4.043861e-13, 4.034306e-13, 4.041933e-13, 4.030009e-13, 
    4.039926e-13, 4.024215e-13, 4.057883e-13, 4.040257e-13, 4.076161e-13, 
    4.071416e-13, 4.063403e-13, 4.047631e-13, 4.055712e-13, 4.046358e-13, 
    4.068894e-13, 4.083447e-13, 4.087561e-13, 4.095631e-13, 4.087383e-13, 
    4.088033e-13, 4.080604e-13, 4.082939e-13, 4.06666e-13, 4.075073e-13, 
    4.053069e-13, 4.046427e-13, 4.031228e-13, 4.024239e-13, 4.018712e-13, 
    4.016731e-13, 4.01618e-13, 4.015957e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 
    8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949652e-07, 
    8.949654e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949652e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949654e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 
    8.949653e-07, 8.949653e-07, 8.949654e-07, 8.949653e-07, 8.949655e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.94965e-07, 8.94965e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949651e-07, 8.949652e-07, 8.94965e-07, 8.94965e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949653e-07, 8.949652e-07, 8.949653e-07, 8.949651e-07, 8.949652e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949654e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.94965e-07, 8.949652e-07, 8.949652e-07, 8.949654e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.94965e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.787388e-16, 6.805754e-16, 6.802186e-16, 6.816986e-16, 6.80878e-16, 
    6.818466e-16, 6.791115e-16, 6.80648e-16, 6.796675e-16, 6.789045e-16, 
    6.845663e-16, 6.817646e-16, 6.874738e-16, 6.856903e-16, 6.901676e-16, 
    6.87196e-16, 6.907663e-16, 6.900826e-16, 6.921408e-16, 6.915515e-16, 
    6.9418e-16, 6.924128e-16, 6.955418e-16, 6.937585e-16, 6.940374e-16, 
    6.923544e-16, 6.823293e-16, 6.842175e-16, 6.822173e-16, 6.824867e-16, 
    6.823659e-16, 6.808947e-16, 6.801525e-16, 6.785987e-16, 6.78881e-16, 
    6.800224e-16, 6.826079e-16, 6.81731e-16, 6.839411e-16, 6.838912e-16, 
    6.86348e-16, 6.852408e-16, 6.89365e-16, 6.88194e-16, 6.915761e-16, 
    6.907261e-16, 6.915361e-16, 6.912906e-16, 6.915393e-16, 6.902926e-16, 
    6.908268e-16, 6.897295e-16, 6.854481e-16, 6.867073e-16, 6.829485e-16, 
    6.806835e-16, 6.791789e-16, 6.781099e-16, 6.782611e-16, 6.785491e-16, 
    6.800291e-16, 6.814198e-16, 6.824789e-16, 6.831868e-16, 6.838841e-16, 
    6.859915e-16, 6.871071e-16, 6.896014e-16, 6.89152e-16, 6.899136e-16, 
    6.906416e-16, 6.918623e-16, 6.916615e-16, 6.921989e-16, 6.898939e-16, 
    6.914261e-16, 6.888959e-16, 6.895883e-16, 6.840717e-16, 6.819677e-16, 
    6.81071e-16, 6.802872e-16, 6.783773e-16, 6.796963e-16, 6.791764e-16, 
    6.804134e-16, 6.811988e-16, 6.808105e-16, 6.832061e-16, 6.822751e-16, 
    6.871733e-16, 6.850652e-16, 6.905567e-16, 6.892444e-16, 6.908711e-16, 
    6.900413e-16, 6.914627e-16, 6.901836e-16, 6.923991e-16, 6.928809e-16, 
    6.925516e-16, 6.938168e-16, 6.901126e-16, 6.915359e-16, 6.807995e-16, 
    6.808628e-16, 6.81158e-16, 6.7986e-16, 6.797807e-16, 6.785909e-16, 
    6.796498e-16, 6.801004e-16, 6.812444e-16, 6.819204e-16, 6.825629e-16, 
    6.839747e-16, 6.855497e-16, 6.877501e-16, 6.893294e-16, 6.903872e-16, 
    6.897388e-16, 6.903113e-16, 6.896712e-16, 6.893713e-16, 6.927003e-16, 
    6.908317e-16, 6.936349e-16, 6.9348e-16, 6.922116e-16, 6.934974e-16, 
    6.809073e-16, 6.805429e-16, 6.792762e-16, 6.802676e-16, 6.784613e-16, 
    6.794723e-16, 6.800533e-16, 6.822941e-16, 6.827865e-16, 6.832424e-16, 
    6.841428e-16, 6.852975e-16, 6.873209e-16, 6.890797e-16, 6.90684e-16, 
    6.905666e-16, 6.906079e-16, 6.909659e-16, 6.900787e-16, 6.911115e-16, 
    6.912846e-16, 6.908317e-16, 6.934592e-16, 6.92709e-16, 6.934767e-16, 
    6.929883e-16, 6.806614e-16, 6.812746e-16, 6.809432e-16, 6.815663e-16, 
    6.811272e-16, 6.83078e-16, 6.836625e-16, 6.863951e-16, 6.852746e-16, 
    6.87058e-16, 6.85456e-16, 6.857399e-16, 6.871153e-16, 6.855427e-16, 
    6.889824e-16, 6.866505e-16, 6.909798e-16, 6.886531e-16, 6.911254e-16, 
    6.906771e-16, 6.914195e-16, 6.920839e-16, 6.929199e-16, 6.944604e-16, 
    6.941038e-16, 6.953917e-16, 6.821886e-16, 6.829832e-16, 6.829136e-16, 
    6.83745e-16, 6.843594e-16, 6.85691e-16, 6.878239e-16, 6.870223e-16, 
    6.884941e-16, 6.887893e-16, 6.865533e-16, 6.879262e-16, 6.83515e-16, 
    6.842281e-16, 6.838038e-16, 6.822512e-16, 6.872066e-16, 6.84665e-16, 
    6.893554e-16, 6.87981e-16, 6.919892e-16, 6.899967e-16, 6.939075e-16, 
    6.955754e-16, 6.971451e-16, 6.989756e-16, 6.83417e-16, 6.828773e-16, 
    6.838439e-16, 6.851796e-16, 6.86419e-16, 6.880648e-16, 6.882333e-16, 
    6.885413e-16, 6.893392e-16, 6.900097e-16, 6.886383e-16, 6.901777e-16, 
    6.843927e-16, 6.874272e-16, 6.826729e-16, 6.841054e-16, 6.851011e-16, 
    6.846648e-16, 6.869308e-16, 6.874642e-16, 6.896302e-16, 6.885111e-16, 
    6.951635e-16, 6.922238e-16, 7.00369e-16, 6.980969e-16, 6.826886e-16, 
    6.834154e-16, 6.859416e-16, 6.847402e-16, 6.881748e-16, 6.89019e-16, 
    6.897052e-16, 6.905815e-16, 6.906763e-16, 6.911952e-16, 6.903447e-16, 
    6.911618e-16, 6.880683e-16, 6.894515e-16, 6.856535e-16, 6.865785e-16, 
    6.861531e-16, 6.856862e-16, 6.871269e-16, 6.886598e-16, 6.886931e-16, 
    6.891842e-16, 6.905664e-16, 6.881887e-16, 6.955415e-16, 6.910037e-16, 
    6.842074e-16, 6.856049e-16, 6.858051e-16, 6.852638e-16, 6.889343e-16, 
    6.876053e-16, 6.911826e-16, 6.902167e-16, 6.917992e-16, 6.91013e-16, 
    6.908972e-16, 6.898869e-16, 6.892574e-16, 6.876661e-16, 6.863703e-16, 
    6.853424e-16, 6.855815e-16, 6.867105e-16, 6.887537e-16, 6.906846e-16, 
    6.902618e-16, 6.91679e-16, 6.87926e-16, 6.895004e-16, 6.888919e-16, 
    6.904783e-16, 6.870009e-16, 6.899608e-16, 6.862432e-16, 6.865696e-16, 
    6.875788e-16, 6.896068e-16, 6.90056e-16, 6.905345e-16, 6.902394e-16, 
    6.888056e-16, 6.885708e-16, 6.875545e-16, 6.872734e-16, 6.864986e-16, 
    6.858566e-16, 6.864431e-16, 6.870586e-16, 6.888065e-16, 6.903797e-16, 
    6.920933e-16, 6.925126e-16, 6.945105e-16, 6.928836e-16, 6.955666e-16, 
    6.932846e-16, 6.972334e-16, 6.901331e-16, 6.932186e-16, 6.876249e-16, 
    6.882286e-16, 6.893193e-16, 6.918195e-16, 6.904709e-16, 6.920482e-16, 
    6.885617e-16, 6.867492e-16, 6.862806e-16, 6.854048e-16, 6.863006e-16, 
    6.862278e-16, 6.870845e-16, 6.868093e-16, 6.888644e-16, 6.877608e-16, 
    6.908942e-16, 6.920359e-16, 6.952565e-16, 6.972271e-16, 6.992314e-16, 
    7.001151e-16, 7.00384e-16, 7.004964e-16 ;

 CWDC_TO_LITR2C =
  5.158415e-16, 5.172373e-16, 5.169662e-16, 5.180909e-16, 5.174673e-16, 
    5.182035e-16, 5.161248e-16, 5.172925e-16, 5.165473e-16, 5.159674e-16, 
    5.202703e-16, 5.181411e-16, 5.224801e-16, 5.211246e-16, 5.245274e-16, 
    5.22269e-16, 5.249823e-16, 5.244628e-16, 5.26027e-16, 5.255791e-16, 
    5.275768e-16, 5.262337e-16, 5.286118e-16, 5.272565e-16, 5.274684e-16, 
    5.261893e-16, 5.185703e-16, 5.200053e-16, 5.184851e-16, 5.186899e-16, 
    5.185981e-16, 5.1748e-16, 5.169159e-16, 5.15735e-16, 5.159496e-16, 
    5.16817e-16, 5.18782e-16, 5.181155e-16, 5.197953e-16, 5.197574e-16, 
    5.216245e-16, 5.20783e-16, 5.239174e-16, 5.230274e-16, 5.255978e-16, 
    5.249519e-16, 5.255674e-16, 5.253809e-16, 5.255699e-16, 5.246223e-16, 
    5.250284e-16, 5.241944e-16, 5.209406e-16, 5.218976e-16, 5.190409e-16, 
    5.173195e-16, 5.161759e-16, 5.153635e-16, 5.154784e-16, 5.156973e-16, 
    5.168221e-16, 5.178791e-16, 5.186839e-16, 5.192219e-16, 5.197519e-16, 
    5.213536e-16, 5.222014e-16, 5.240971e-16, 5.237556e-16, 5.243344e-16, 
    5.248876e-16, 5.258153e-16, 5.256627e-16, 5.260712e-16, 5.243194e-16, 
    5.254838e-16, 5.235609e-16, 5.240871e-16, 5.198945e-16, 5.182954e-16, 
    5.176139e-16, 5.170182e-16, 5.155667e-16, 5.165692e-16, 5.16174e-16, 
    5.171142e-16, 5.17711e-16, 5.17416e-16, 5.192366e-16, 5.185291e-16, 
    5.222517e-16, 5.206496e-16, 5.248231e-16, 5.238257e-16, 5.250621e-16, 
    5.244314e-16, 5.255117e-16, 5.245395e-16, 5.262233e-16, 5.265895e-16, 
    5.263392e-16, 5.273007e-16, 5.244856e-16, 5.255673e-16, 5.174076e-16, 
    5.174558e-16, 5.176801e-16, 5.166936e-16, 5.166333e-16, 5.15729e-16, 
    5.165338e-16, 5.168763e-16, 5.177458e-16, 5.182595e-16, 5.187478e-16, 
    5.198207e-16, 5.210177e-16, 5.226901e-16, 5.238904e-16, 5.246942e-16, 
    5.242015e-16, 5.246365e-16, 5.241501e-16, 5.239222e-16, 5.264522e-16, 
    5.250321e-16, 5.271625e-16, 5.270448e-16, 5.260808e-16, 5.27058e-16, 
    5.174895e-16, 5.172126e-16, 5.1625e-16, 5.170033e-16, 5.156306e-16, 
    5.16399e-16, 5.168405e-16, 5.185435e-16, 5.189177e-16, 5.192642e-16, 
    5.199485e-16, 5.208261e-16, 5.223638e-16, 5.237006e-16, 5.249199e-16, 
    5.248306e-16, 5.24862e-16, 5.251341e-16, 5.244598e-16, 5.252447e-16, 
    5.253763e-16, 5.250321e-16, 5.27029e-16, 5.264589e-16, 5.270423e-16, 
    5.266711e-16, 5.173027e-16, 5.177687e-16, 5.175169e-16, 5.179903e-16, 
    5.176567e-16, 5.191393e-16, 5.195835e-16, 5.216602e-16, 5.208087e-16, 
    5.22164e-16, 5.209465e-16, 5.211623e-16, 5.222077e-16, 5.210125e-16, 
    5.236267e-16, 5.218544e-16, 5.251447e-16, 5.233764e-16, 5.252553e-16, 
    5.249146e-16, 5.254788e-16, 5.259838e-16, 5.266191e-16, 5.277899e-16, 
    5.275189e-16, 5.284976e-16, 5.184634e-16, 5.190672e-16, 5.190143e-16, 
    5.196461e-16, 5.201132e-16, 5.211252e-16, 5.227462e-16, 5.221369e-16, 
    5.232555e-16, 5.234799e-16, 5.217806e-16, 5.228239e-16, 5.194714e-16, 
    5.200133e-16, 5.196909e-16, 5.185108e-16, 5.22277e-16, 5.203454e-16, 
    5.239102e-16, 5.228656e-16, 5.259118e-16, 5.243975e-16, 5.273697e-16, 
    5.286373e-16, 5.298303e-16, 5.312214e-16, 5.19397e-16, 5.189868e-16, 
    5.197214e-16, 5.207365e-16, 5.216785e-16, 5.229292e-16, 5.230573e-16, 
    5.232913e-16, 5.238978e-16, 5.244073e-16, 5.233651e-16, 5.245351e-16, 
    5.201385e-16, 5.224446e-16, 5.188314e-16, 5.199202e-16, 5.206768e-16, 
    5.203452e-16, 5.220674e-16, 5.224728e-16, 5.24119e-16, 5.232684e-16, 
    5.283243e-16, 5.2609e-16, 5.322805e-16, 5.305536e-16, 5.188434e-16, 
    5.193957e-16, 5.213156e-16, 5.204025e-16, 5.230128e-16, 5.236544e-16, 
    5.241759e-16, 5.248419e-16, 5.24914e-16, 5.253083e-16, 5.24662e-16, 
    5.252829e-16, 5.229319e-16, 5.239831e-16, 5.210966e-16, 5.217997e-16, 
    5.214764e-16, 5.211215e-16, 5.222164e-16, 5.233814e-16, 5.234068e-16, 
    5.2378e-16, 5.248305e-16, 5.230234e-16, 5.286116e-16, 5.251628e-16, 
    5.199976e-16, 5.210597e-16, 5.212119e-16, 5.208005e-16, 5.235901e-16, 
    5.2258e-16, 5.252988e-16, 5.245647e-16, 5.257674e-16, 5.251699e-16, 
    5.250819e-16, 5.24314e-16, 5.238356e-16, 5.226262e-16, 5.216414e-16, 
    5.208602e-16, 5.210419e-16, 5.219e-16, 5.234528e-16, 5.249203e-16, 
    5.24599e-16, 5.256761e-16, 5.228237e-16, 5.240203e-16, 5.235578e-16, 
    5.247635e-16, 5.221206e-16, 5.243702e-16, 5.215449e-16, 5.217929e-16, 
    5.225599e-16, 5.241012e-16, 5.244426e-16, 5.248062e-16, 5.245819e-16, 
    5.234922e-16, 5.233138e-16, 5.225414e-16, 5.223278e-16, 5.217389e-16, 
    5.21251e-16, 5.216967e-16, 5.221645e-16, 5.234929e-16, 5.246886e-16, 
    5.259909e-16, 5.263096e-16, 5.27828e-16, 5.265915e-16, 5.286306e-16, 
    5.268963e-16, 5.298974e-16, 5.245011e-16, 5.268462e-16, 5.22595e-16, 
    5.230538e-16, 5.238827e-16, 5.257828e-16, 5.247579e-16, 5.259566e-16, 
    5.233069e-16, 5.219294e-16, 5.215732e-16, 5.209076e-16, 5.215884e-16, 
    5.215331e-16, 5.221842e-16, 5.219751e-16, 5.23537e-16, 5.226983e-16, 
    5.250796e-16, 5.259473e-16, 5.283949e-16, 5.298926e-16, 5.314159e-16, 
    5.320875e-16, 5.322919e-16, 5.323773e-16 ;

 CWDC_TO_LITR3C =
  1.628973e-16, 1.633381e-16, 1.632525e-16, 1.636077e-16, 1.634107e-16, 
    1.636432e-16, 1.629868e-16, 1.633555e-16, 1.631202e-16, 1.629371e-16, 
    1.642959e-16, 1.636235e-16, 1.649937e-16, 1.645657e-16, 1.656402e-16, 
    1.649271e-16, 1.657839e-16, 1.656198e-16, 1.661138e-16, 1.659724e-16, 
    1.666032e-16, 1.661791e-16, 1.6693e-16, 1.66502e-16, 1.66569e-16, 
    1.66165e-16, 1.637591e-16, 1.642122e-16, 1.637321e-16, 1.637968e-16, 
    1.637678e-16, 1.634147e-16, 1.632366e-16, 1.628637e-16, 1.629314e-16, 
    1.632054e-16, 1.638259e-16, 1.636154e-16, 1.641459e-16, 1.641339e-16, 
    1.647235e-16, 1.644578e-16, 1.654476e-16, 1.651666e-16, 1.659783e-16, 
    1.657743e-16, 1.659687e-16, 1.659097e-16, 1.659694e-16, 1.656702e-16, 
    1.657984e-16, 1.655351e-16, 1.645075e-16, 1.648098e-16, 1.639077e-16, 
    1.633641e-16, 1.630029e-16, 1.627464e-16, 1.627827e-16, 1.628518e-16, 
    1.63207e-16, 1.635408e-16, 1.637949e-16, 1.639648e-16, 1.641322e-16, 
    1.64638e-16, 1.649057e-16, 1.655043e-16, 1.653965e-16, 1.655793e-16, 
    1.65754e-16, 1.66047e-16, 1.659988e-16, 1.661278e-16, 1.655745e-16, 
    1.659423e-16, 1.65335e-16, 1.655012e-16, 1.641772e-16, 1.636722e-16, 
    1.63457e-16, 1.632689e-16, 1.628105e-16, 1.631271e-16, 1.630023e-16, 
    1.632992e-16, 1.634877e-16, 1.633945e-16, 1.639695e-16, 1.63746e-16, 
    1.649216e-16, 1.644157e-16, 1.657336e-16, 1.654186e-16, 1.658091e-16, 
    1.656099e-16, 1.659511e-16, 1.656441e-16, 1.661758e-16, 1.662914e-16, 
    1.662124e-16, 1.66516e-16, 1.65627e-16, 1.659686e-16, 1.633919e-16, 
    1.634071e-16, 1.634779e-16, 1.631664e-16, 1.631474e-16, 1.628618e-16, 
    1.63116e-16, 1.632241e-16, 1.634987e-16, 1.636609e-16, 1.638151e-16, 
    1.641539e-16, 1.645319e-16, 1.6506e-16, 1.654391e-16, 1.656929e-16, 
    1.655373e-16, 1.656747e-16, 1.655211e-16, 1.654491e-16, 1.662481e-16, 
    1.657996e-16, 1.664724e-16, 1.664352e-16, 1.661308e-16, 1.664394e-16, 
    1.634177e-16, 1.633303e-16, 1.630263e-16, 1.632642e-16, 1.628307e-16, 
    1.630734e-16, 1.632128e-16, 1.637506e-16, 1.638688e-16, 1.639782e-16, 
    1.641943e-16, 1.644714e-16, 1.64957e-16, 1.653791e-16, 1.657642e-16, 
    1.65736e-16, 1.657459e-16, 1.658318e-16, 1.656189e-16, 1.658668e-16, 
    1.659083e-16, 1.657996e-16, 1.664302e-16, 1.662502e-16, 1.664344e-16, 
    1.663172e-16, 1.633587e-16, 1.635059e-16, 1.634264e-16, 1.635759e-16, 
    1.634705e-16, 1.639387e-16, 1.64079e-16, 1.647348e-16, 1.644659e-16, 
    1.648939e-16, 1.645094e-16, 1.645776e-16, 1.649077e-16, 1.645303e-16, 
    1.653558e-16, 1.647961e-16, 1.658351e-16, 1.652767e-16, 1.658701e-16, 
    1.657625e-16, 1.659407e-16, 1.661001e-16, 1.663008e-16, 1.666705e-16, 
    1.665849e-16, 1.66894e-16, 1.637253e-16, 1.63916e-16, 1.638993e-16, 
    1.640988e-16, 1.642463e-16, 1.645658e-16, 1.650777e-16, 1.648854e-16, 
    1.652386e-16, 1.653094e-16, 1.647728e-16, 1.651023e-16, 1.640436e-16, 
    1.642147e-16, 1.641129e-16, 1.637403e-16, 1.649296e-16, 1.643196e-16, 
    1.654453e-16, 1.651154e-16, 1.660774e-16, 1.655992e-16, 1.665378e-16, 
    1.669381e-16, 1.673148e-16, 1.677541e-16, 1.640201e-16, 1.638906e-16, 
    1.641225e-16, 1.644431e-16, 1.647406e-16, 1.651355e-16, 1.65176e-16, 
    1.652499e-16, 1.654414e-16, 1.656023e-16, 1.652732e-16, 1.656427e-16, 
    1.642542e-16, 1.649825e-16, 1.638415e-16, 1.641853e-16, 1.644243e-16, 
    1.643195e-16, 1.648634e-16, 1.649914e-16, 1.655113e-16, 1.652427e-16, 
    1.668393e-16, 1.661337e-16, 1.680886e-16, 1.675433e-16, 1.638453e-16, 
    1.640197e-16, 1.64626e-16, 1.643376e-16, 1.651619e-16, 1.653645e-16, 
    1.655292e-16, 1.657395e-16, 1.657623e-16, 1.658868e-16, 1.656827e-16, 
    1.658788e-16, 1.651364e-16, 1.654683e-16, 1.645568e-16, 1.647788e-16, 
    1.646768e-16, 1.645647e-16, 1.649104e-16, 1.652783e-16, 1.652863e-16, 
    1.654042e-16, 1.657359e-16, 1.651653e-16, 1.6693e-16, 1.658409e-16, 
    1.642098e-16, 1.645452e-16, 1.645932e-16, 1.644633e-16, 1.653442e-16, 
    1.650253e-16, 1.658838e-16, 1.65652e-16, 1.660318e-16, 1.658431e-16, 
    1.658153e-16, 1.655729e-16, 1.654218e-16, 1.650399e-16, 1.647289e-16, 
    1.644822e-16, 1.645396e-16, 1.648105e-16, 1.653009e-16, 1.657643e-16, 
    1.656628e-16, 1.66003e-16, 1.651022e-16, 1.654801e-16, 1.653341e-16, 
    1.657148e-16, 1.648802e-16, 1.655906e-16, 1.646984e-16, 1.647767e-16, 
    1.650189e-16, 1.655056e-16, 1.656134e-16, 1.657283e-16, 1.656574e-16, 
    1.653133e-16, 1.65257e-16, 1.650131e-16, 1.649456e-16, 1.647597e-16, 
    1.646056e-16, 1.647463e-16, 1.648941e-16, 1.653135e-16, 1.656911e-16, 
    1.661024e-16, 1.66203e-16, 1.666825e-16, 1.662921e-16, 1.66936e-16, 
    1.663883e-16, 1.67336e-16, 1.656319e-16, 1.663725e-16, 1.6503e-16, 
    1.651749e-16, 1.654366e-16, 1.660367e-16, 1.65713e-16, 1.660916e-16, 
    1.652548e-16, 1.648198e-16, 1.647073e-16, 1.644972e-16, 1.647121e-16, 
    1.646947e-16, 1.649003e-16, 1.648342e-16, 1.653275e-16, 1.650626e-16, 
    1.658146e-16, 1.660886e-16, 1.668616e-16, 1.673345e-16, 1.678155e-16, 
    1.680276e-16, 1.680922e-16, 1.681191e-16 ;

 CWDC_vr =
  5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110344e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110343e-05, 5.110344e-05, 5.110342e-05, 5.110343e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110343e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  1.031683e-18, 1.034475e-18, 1.033932e-18, 1.036182e-18, 1.034935e-18, 
    1.036407e-18, 1.03225e-18, 1.034585e-18, 1.033095e-18, 1.031935e-18, 
    1.040541e-18, 1.036282e-18, 1.04496e-18, 1.042249e-18, 1.049055e-18, 
    1.044538e-18, 1.049965e-18, 1.048926e-18, 1.052054e-18, 1.051158e-18, 
    1.055154e-18, 1.052467e-18, 1.057223e-18, 1.054513e-18, 1.054937e-18, 
    1.052379e-18, 1.037141e-18, 1.040011e-18, 1.03697e-18, 1.03738e-18, 
    1.037196e-18, 1.03496e-18, 1.033832e-18, 1.03147e-18, 1.031899e-18, 
    1.033634e-18, 1.037564e-18, 1.036231e-18, 1.03959e-18, 1.039515e-18, 
    1.043249e-18, 1.041566e-18, 1.047835e-18, 1.046055e-18, 1.051196e-18, 
    1.049904e-18, 1.051135e-18, 1.050762e-18, 1.05114e-18, 1.049245e-18, 
    1.050057e-18, 1.048389e-18, 1.041881e-18, 1.043795e-18, 1.038082e-18, 
    1.034639e-18, 1.032352e-18, 1.030727e-18, 1.030957e-18, 1.031395e-18, 
    1.033644e-18, 1.035758e-18, 1.037368e-18, 1.038444e-18, 1.039504e-18, 
    1.042707e-18, 1.044403e-18, 1.048194e-18, 1.047511e-18, 1.048669e-18, 
    1.049775e-18, 1.051631e-18, 1.051325e-18, 1.052142e-18, 1.048639e-18, 
    1.050968e-18, 1.047122e-18, 1.048174e-18, 1.039789e-18, 1.036591e-18, 
    1.035228e-18, 1.034036e-18, 1.031133e-18, 1.033138e-18, 1.032348e-18, 
    1.034228e-18, 1.035422e-18, 1.034832e-18, 1.038473e-18, 1.037058e-18, 
    1.044503e-18, 1.041299e-18, 1.049646e-18, 1.047651e-18, 1.050124e-18, 
    1.048863e-18, 1.051023e-18, 1.049079e-18, 1.052447e-18, 1.053179e-18, 
    1.052678e-18, 1.054602e-18, 1.048971e-18, 1.051135e-18, 1.034815e-18, 
    1.034912e-18, 1.03536e-18, 1.033387e-18, 1.033267e-18, 1.031458e-18, 
    1.033068e-18, 1.033753e-18, 1.035491e-18, 1.036519e-18, 1.037496e-18, 
    1.039641e-18, 1.042036e-18, 1.04538e-18, 1.047781e-18, 1.049389e-18, 
    1.048403e-18, 1.049273e-18, 1.0483e-18, 1.047844e-18, 1.052904e-18, 
    1.050064e-18, 1.054325e-18, 1.054089e-18, 1.052162e-18, 1.054116e-18, 
    1.034979e-18, 1.034425e-18, 1.0325e-18, 1.034007e-18, 1.031261e-18, 
    1.032798e-18, 1.033681e-18, 1.037087e-18, 1.037835e-18, 1.038528e-18, 
    1.039897e-18, 1.041652e-18, 1.044728e-18, 1.047401e-18, 1.04984e-18, 
    1.049661e-18, 1.049724e-18, 1.050268e-18, 1.04892e-18, 1.050489e-18, 
    1.050753e-18, 1.050064e-18, 1.054058e-18, 1.052918e-18, 1.054085e-18, 
    1.053342e-18, 1.034605e-18, 1.035537e-18, 1.035034e-18, 1.035981e-18, 
    1.035313e-18, 1.038279e-18, 1.039167e-18, 1.043321e-18, 1.041617e-18, 
    1.044328e-18, 1.041893e-18, 1.042325e-18, 1.044415e-18, 1.042025e-18, 
    1.047253e-18, 1.043709e-18, 1.050289e-18, 1.046753e-18, 1.050511e-18, 
    1.049829e-18, 1.050958e-18, 1.051968e-18, 1.053238e-18, 1.05558e-18, 
    1.055038e-18, 1.056995e-18, 1.036927e-18, 1.038134e-18, 1.038029e-18, 
    1.039292e-18, 1.040226e-18, 1.04225e-18, 1.045492e-18, 1.044274e-18, 
    1.046511e-18, 1.04696e-18, 1.043561e-18, 1.045648e-18, 1.038943e-18, 
    1.040027e-18, 1.039382e-18, 1.037022e-18, 1.044554e-18, 1.040691e-18, 
    1.04782e-18, 1.045731e-18, 1.051824e-18, 1.048795e-18, 1.054739e-18, 
    1.057275e-18, 1.059661e-18, 1.062443e-18, 1.038794e-18, 1.037974e-18, 
    1.039443e-18, 1.041473e-18, 1.043357e-18, 1.045858e-18, 1.046115e-18, 
    1.046583e-18, 1.047796e-18, 1.048815e-18, 1.04673e-18, 1.04907e-18, 
    1.040277e-18, 1.044889e-18, 1.037663e-18, 1.03984e-18, 1.041354e-18, 
    1.04069e-18, 1.044135e-18, 1.044946e-18, 1.048238e-18, 1.046537e-18, 
    1.056649e-18, 1.05218e-18, 1.064561e-18, 1.061107e-18, 1.037687e-18, 
    1.038791e-18, 1.042631e-18, 1.040805e-18, 1.046026e-18, 1.047309e-18, 
    1.048352e-18, 1.049684e-18, 1.049828e-18, 1.050617e-18, 1.049324e-18, 
    1.050566e-18, 1.045864e-18, 1.047966e-18, 1.042193e-18, 1.043599e-18, 
    1.042953e-18, 1.042243e-18, 1.044433e-18, 1.046763e-18, 1.046814e-18, 
    1.04756e-18, 1.049661e-18, 1.046047e-18, 1.057223e-18, 1.050326e-18, 
    1.039995e-18, 1.042119e-18, 1.042424e-18, 1.041601e-18, 1.04718e-18, 
    1.04516e-18, 1.050598e-18, 1.049129e-18, 1.051535e-18, 1.05034e-18, 
    1.050164e-18, 1.048628e-18, 1.047671e-18, 1.045252e-18, 1.043283e-18, 
    1.04172e-18, 1.042084e-18, 1.0438e-18, 1.046906e-18, 1.049841e-18, 
    1.049198e-18, 1.051352e-18, 1.045647e-18, 1.048041e-18, 1.047116e-18, 
    1.049527e-18, 1.044241e-18, 1.04874e-18, 1.04309e-18, 1.043586e-18, 
    1.04512e-18, 1.048202e-18, 1.048885e-18, 1.049612e-18, 1.049164e-18, 
    1.046985e-18, 1.046628e-18, 1.045083e-18, 1.044656e-18, 1.043478e-18, 
    1.042502e-18, 1.043393e-18, 1.044329e-18, 1.046986e-18, 1.049377e-18, 
    1.051982e-18, 1.052619e-18, 1.055656e-18, 1.053183e-18, 1.057261e-18, 
    1.053793e-18, 1.059795e-18, 1.049002e-18, 1.053692e-18, 1.04519e-18, 
    1.046108e-18, 1.047765e-18, 1.051566e-18, 1.049516e-18, 1.051913e-18, 
    1.046614e-18, 1.043859e-18, 1.043147e-18, 1.041815e-18, 1.043177e-18, 
    1.043066e-18, 1.044368e-18, 1.04395e-18, 1.047074e-18, 1.045396e-18, 
    1.050159e-18, 1.051895e-18, 1.05679e-18, 1.059785e-18, 1.062832e-18, 
    1.064175e-18, 1.064584e-18, 1.064755e-18 ;

 CWDN_TO_LITR3N =
  3.257946e-19, 3.266762e-19, 3.265049e-19, 3.272153e-19, 3.268214e-19, 
    3.272864e-19, 3.259735e-19, 3.267111e-19, 3.262404e-19, 3.258742e-19, 
    3.285918e-19, 3.27247e-19, 3.299874e-19, 3.291313e-19, 3.312805e-19, 
    3.298541e-19, 3.315678e-19, 3.312396e-19, 3.322276e-19, 3.319447e-19, 
    3.332064e-19, 3.323581e-19, 3.3386e-19, 3.330041e-19, 3.331379e-19, 
    3.323301e-19, 3.275181e-19, 3.284244e-19, 3.274643e-19, 3.275936e-19, 
    3.275357e-19, 3.268295e-19, 3.264732e-19, 3.257274e-19, 3.258629e-19, 
    3.264107e-19, 3.276518e-19, 3.272309e-19, 3.282917e-19, 3.282678e-19, 
    3.294471e-19, 3.289156e-19, 3.308952e-19, 3.303331e-19, 3.319565e-19, 
    3.315485e-19, 3.319373e-19, 3.318195e-19, 3.319389e-19, 3.313404e-19, 
    3.315969e-19, 3.310701e-19, 3.290151e-19, 3.296195e-19, 3.278153e-19, 
    3.267281e-19, 3.260058e-19, 3.254928e-19, 3.255653e-19, 3.257036e-19, 
    3.264139e-19, 3.270815e-19, 3.275898e-19, 3.279297e-19, 3.282644e-19, 
    3.292759e-19, 3.298114e-19, 3.310087e-19, 3.30793e-19, 3.311586e-19, 
    3.31508e-19, 3.320939e-19, 3.319975e-19, 3.322555e-19, 3.311491e-19, 
    3.318845e-19, 3.306701e-19, 3.310024e-19, 3.283544e-19, 3.273445e-19, 
    3.269141e-19, 3.265378e-19, 3.256211e-19, 3.262542e-19, 3.260047e-19, 
    3.265985e-19, 3.269754e-19, 3.26789e-19, 3.279389e-19, 3.27492e-19, 
    3.298432e-19, 3.288313e-19, 3.314672e-19, 3.308373e-19, 3.316182e-19, 
    3.312198e-19, 3.319021e-19, 3.312881e-19, 3.323516e-19, 3.325829e-19, 
    3.324248e-19, 3.33032e-19, 3.31254e-19, 3.319372e-19, 3.267837e-19, 
    3.268141e-19, 3.269559e-19, 3.263328e-19, 3.262947e-19, 3.257236e-19, 
    3.262319e-19, 3.264482e-19, 3.269973e-19, 3.273218e-19, 3.276302e-19, 
    3.283078e-19, 3.290638e-19, 3.301201e-19, 3.308781e-19, 3.313858e-19, 
    3.310746e-19, 3.313494e-19, 3.310422e-19, 3.308982e-19, 3.324961e-19, 
    3.315992e-19, 3.329447e-19, 3.328704e-19, 3.322616e-19, 3.328788e-19, 
    3.268355e-19, 3.266606e-19, 3.260526e-19, 3.265284e-19, 3.256614e-19, 
    3.261467e-19, 3.264256e-19, 3.275012e-19, 3.277375e-19, 3.279564e-19, 
    3.283886e-19, 3.289428e-19, 3.29914e-19, 3.307583e-19, 3.315283e-19, 
    3.31472e-19, 3.314918e-19, 3.316636e-19, 3.312378e-19, 3.317335e-19, 
    3.318166e-19, 3.315992e-19, 3.328604e-19, 3.325003e-19, 3.328688e-19, 
    3.326344e-19, 3.267175e-19, 3.270118e-19, 3.268528e-19, 3.271518e-19, 
    3.269411e-19, 3.278774e-19, 3.28158e-19, 3.294696e-19, 3.289318e-19, 
    3.297878e-19, 3.290189e-19, 3.291551e-19, 3.298154e-19, 3.290605e-19, 
    3.307116e-19, 3.295922e-19, 3.316703e-19, 3.305535e-19, 3.317402e-19, 
    3.31525e-19, 3.318814e-19, 3.322003e-19, 3.326015e-19, 3.33341e-19, 
    3.331699e-19, 3.33788e-19, 3.274506e-19, 3.278319e-19, 3.277985e-19, 
    3.281976e-19, 3.284925e-19, 3.291317e-19, 3.301555e-19, 3.297707e-19, 
    3.304772e-19, 3.306189e-19, 3.295456e-19, 3.302046e-19, 3.280872e-19, 
    3.284295e-19, 3.282258e-19, 3.274805e-19, 3.298592e-19, 3.286392e-19, 
    3.308906e-19, 3.302309e-19, 3.321548e-19, 3.311984e-19, 3.330756e-19, 
    3.338762e-19, 3.346297e-19, 3.355083e-19, 3.280402e-19, 3.277811e-19, 
    3.282451e-19, 3.288862e-19, 3.294811e-19, 3.302711e-19, 3.30352e-19, 
    3.304998e-19, 3.308828e-19, 3.312046e-19, 3.305464e-19, 3.312853e-19, 
    3.285085e-19, 3.29965e-19, 3.27683e-19, 3.283706e-19, 3.288485e-19, 
    3.286391e-19, 3.297268e-19, 3.299828e-19, 3.310225e-19, 3.304853e-19, 
    3.336785e-19, 3.322674e-19, 3.361771e-19, 3.350865e-19, 3.276905e-19, 
    3.280394e-19, 3.29252e-19, 3.286753e-19, 3.303239e-19, 3.307291e-19, 
    3.310585e-19, 3.314791e-19, 3.315246e-19, 3.317737e-19, 3.313655e-19, 
    3.317576e-19, 3.302728e-19, 3.309367e-19, 3.291137e-19, 3.295577e-19, 
    3.293535e-19, 3.291294e-19, 3.298209e-19, 3.305567e-19, 3.305727e-19, 
    3.308084e-19, 3.314718e-19, 3.303306e-19, 3.338599e-19, 3.316817e-19, 
    3.284196e-19, 3.290903e-19, 3.291864e-19, 3.289266e-19, 3.306885e-19, 
    3.300505e-19, 3.317677e-19, 3.31304e-19, 3.320636e-19, 3.316862e-19, 
    3.316307e-19, 3.311457e-19, 3.308436e-19, 3.300797e-19, 3.294578e-19, 
    3.289644e-19, 3.290791e-19, 3.29621e-19, 3.306018e-19, 3.315286e-19, 
    3.313256e-19, 3.320059e-19, 3.302045e-19, 3.309602e-19, 3.306681e-19, 
    3.314296e-19, 3.297604e-19, 3.311812e-19, 3.293968e-19, 3.295534e-19, 
    3.300379e-19, 3.310112e-19, 3.312269e-19, 3.314565e-19, 3.313149e-19, 
    3.306267e-19, 3.30514e-19, 3.300261e-19, 3.298913e-19, 3.295193e-19, 
    3.292112e-19, 3.294927e-19, 3.297881e-19, 3.306271e-19, 3.313823e-19, 
    3.322048e-19, 3.324061e-19, 3.333651e-19, 3.325841e-19, 3.33872e-19, 
    3.327766e-19, 3.34672e-19, 3.312639e-19, 3.327449e-19, 3.3006e-19, 
    3.303498e-19, 3.308733e-19, 3.320733e-19, 3.31426e-19, 3.321831e-19, 
    3.305096e-19, 3.296396e-19, 3.294147e-19, 3.289943e-19, 3.294243e-19, 
    3.293893e-19, 3.298006e-19, 3.296684e-19, 3.306549e-19, 3.301252e-19, 
    3.316292e-19, 3.321773e-19, 3.337231e-19, 3.34669e-19, 3.356311e-19, 
    3.360553e-19, 3.361843e-19, 3.362383e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_LH_TOT_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.215762e-08, 6.243169e-08, 6.237841e-08, 6.259947e-08, 6.247685e-08, 
    6.26216e-08, 6.221319e-08, 6.244257e-08, 6.229614e-08, 6.21823e-08, 
    6.302847e-08, 6.260934e-08, 6.346394e-08, 6.319659e-08, 6.386823e-08, 
    6.342233e-08, 6.395815e-08, 6.385538e-08, 6.416472e-08, 6.40761e-08, 
    6.447177e-08, 6.420563e-08, 6.46769e-08, 6.440823e-08, 6.445025e-08, 
    6.419685e-08, 6.269369e-08, 6.297628e-08, 6.267695e-08, 6.271725e-08, 
    6.269916e-08, 6.247938e-08, 6.236861e-08, 6.213668e-08, 6.217878e-08, 
    6.234914e-08, 6.273537e-08, 6.260426e-08, 6.29347e-08, 6.292724e-08, 
    6.329513e-08, 6.312926e-08, 6.374764e-08, 6.357188e-08, 6.40798e-08, 
    6.395206e-08, 6.40738e-08, 6.403688e-08, 6.407428e-08, 6.388693e-08, 
    6.39672e-08, 6.380235e-08, 6.316031e-08, 6.334899e-08, 6.278628e-08, 
    6.244793e-08, 6.222324e-08, 6.20638e-08, 6.208634e-08, 6.212931e-08, 
    6.235014e-08, 6.255778e-08, 6.271602e-08, 6.282187e-08, 6.292617e-08, 
    6.324185e-08, 6.340898e-08, 6.378317e-08, 6.371565e-08, 6.383004e-08, 
    6.393935e-08, 6.412285e-08, 6.409265e-08, 6.417349e-08, 6.382704e-08, 
    6.405729e-08, 6.367719e-08, 6.378114e-08, 6.295448e-08, 6.263964e-08, 
    6.250578e-08, 6.238865e-08, 6.210367e-08, 6.230047e-08, 6.222289e-08, 
    6.240747e-08, 6.252476e-08, 6.246675e-08, 6.282476e-08, 6.268557e-08, 
    6.341888e-08, 6.310301e-08, 6.39266e-08, 6.372951e-08, 6.397384e-08, 
    6.384917e-08, 6.406279e-08, 6.387053e-08, 6.420358e-08, 6.427612e-08, 
    6.422655e-08, 6.441695e-08, 6.385987e-08, 6.40738e-08, 6.246512e-08, 
    6.247458e-08, 6.251866e-08, 6.232491e-08, 6.231306e-08, 6.213552e-08, 
    6.229349e-08, 6.236077e-08, 6.253156e-08, 6.263257e-08, 6.27286e-08, 
    6.293975e-08, 6.317556e-08, 6.350534e-08, 6.374228e-08, 6.390112e-08, 
    6.380372e-08, 6.388971e-08, 6.379359e-08, 6.374854e-08, 6.424895e-08, 
    6.396795e-08, 6.438957e-08, 6.436624e-08, 6.417542e-08, 6.436887e-08, 
    6.248122e-08, 6.242679e-08, 6.223777e-08, 6.238569e-08, 6.211619e-08, 
    6.226703e-08, 6.235377e-08, 6.268847e-08, 6.276202e-08, 6.283021e-08, 
    6.296489e-08, 6.313774e-08, 6.344097e-08, 6.370482e-08, 6.394571e-08, 
    6.392806e-08, 6.393427e-08, 6.398808e-08, 6.385479e-08, 6.400997e-08, 
    6.403601e-08, 6.396792e-08, 6.436311e-08, 6.425022e-08, 6.436574e-08, 
    6.429224e-08, 6.244449e-08, 6.253608e-08, 6.248658e-08, 6.257967e-08, 
    6.251409e-08, 6.280568e-08, 6.289311e-08, 6.330224e-08, 6.313434e-08, 
    6.340156e-08, 6.316149e-08, 6.320403e-08, 6.341026e-08, 6.317446e-08, 
    6.369027e-08, 6.334054e-08, 6.399017e-08, 6.36409e-08, 6.401206e-08, 
    6.394467e-08, 6.405626e-08, 6.415619e-08, 6.428195e-08, 6.451393e-08, 
    6.446022e-08, 6.465423e-08, 6.267265e-08, 6.279146e-08, 6.278102e-08, 
    6.290536e-08, 6.299733e-08, 6.319667e-08, 6.35164e-08, 6.339616e-08, 
    6.361689e-08, 6.366121e-08, 6.332587e-08, 6.353175e-08, 6.2871e-08, 
    6.297773e-08, 6.291419e-08, 6.268202e-08, 6.342385e-08, 6.304312e-08, 
    6.37462e-08, 6.353994e-08, 6.414194e-08, 6.384253e-08, 6.443064e-08, 
    6.468203e-08, 6.491868e-08, 6.51952e-08, 6.285632e-08, 6.277559e-08, 
    6.292016e-08, 6.312016e-08, 6.330577e-08, 6.355251e-08, 6.357777e-08, 
    6.362399e-08, 6.374373e-08, 6.384442e-08, 6.363859e-08, 6.386966e-08, 
    6.300247e-08, 6.345691e-08, 6.274506e-08, 6.295939e-08, 6.310837e-08, 
    6.304303e-08, 6.338242e-08, 6.346242e-08, 6.378748e-08, 6.361945e-08, 
    6.461998e-08, 6.417729e-08, 6.540579e-08, 6.506244e-08, 6.274738e-08, 
    6.285605e-08, 6.323427e-08, 6.305431e-08, 6.356899e-08, 6.369568e-08, 
    6.379868e-08, 6.393034e-08, 6.394456e-08, 6.402257e-08, 6.389474e-08, 
    6.401752e-08, 6.355304e-08, 6.37606e-08, 6.319105e-08, 6.332966e-08, 
    6.326589e-08, 6.319594e-08, 6.341183e-08, 6.364183e-08, 6.364677e-08, 
    6.372051e-08, 6.392831e-08, 6.357108e-08, 6.467708e-08, 6.399399e-08, 
    6.297455e-08, 6.318386e-08, 6.321378e-08, 6.313269e-08, 6.368298e-08, 
    6.348358e-08, 6.402067e-08, 6.387551e-08, 6.411335e-08, 6.399516e-08, 
    6.397777e-08, 6.382598e-08, 6.373148e-08, 6.349272e-08, 6.329847e-08, 
    6.314445e-08, 6.318027e-08, 6.334945e-08, 6.365591e-08, 6.394584e-08, 
    6.388233e-08, 6.409527e-08, 6.353167e-08, 6.376798e-08, 6.367664e-08, 
    6.391483e-08, 6.339297e-08, 6.383731e-08, 6.327939e-08, 6.332831e-08, 
    6.347963e-08, 6.378401e-08, 6.385137e-08, 6.392327e-08, 6.387891e-08, 
    6.366369e-08, 6.362843e-08, 6.347595e-08, 6.343384e-08, 6.331766e-08, 
    6.322146e-08, 6.330935e-08, 6.340164e-08, 6.366378e-08, 6.390003e-08, 
    6.415761e-08, 6.422066e-08, 6.452161e-08, 6.427662e-08, 6.468089e-08, 
    6.433715e-08, 6.493221e-08, 6.386308e-08, 6.432707e-08, 6.348652e-08, 
    6.357706e-08, 6.374083e-08, 6.41165e-08, 6.39137e-08, 6.415087e-08, 
    6.362706e-08, 6.335529e-08, 6.328499e-08, 6.315381e-08, 6.328799e-08, 
    6.327708e-08, 6.340547e-08, 6.336422e-08, 6.367249e-08, 6.35069e-08, 
    6.397733e-08, 6.414901e-08, 6.463389e-08, 6.493114e-08, 6.523376e-08, 
    6.536735e-08, 6.540802e-08, 6.542501e-08 ;

 ERRH2O =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -1.359657e-14, -2.05645e-14, -8.889341e-15, -5.937103e-15, -1.236956e-14, 
    -7.10196e-15, -2.087441e-14, -1.100031e-14, -1.672329e-14, -2.499059e-14, 
    -6.839192e-15, -1.474107e-14, -1.659774e-14, -1.180052e-14, 
    -1.557504e-14, -1.091568e-14, -1.105728e-14, -1.111469e-14, 
    -1.273378e-14, -8.912497e-15, -1.529139e-14, -1.380104e-14, 
    -1.061199e-14, -1.290652e-14, -1.10362e-14, -9.975221e-15, -1.210517e-14, 
    -2.099237e-14, -1.718764e-14, -1.332296e-14, -1.749261e-14, 
    -1.096074e-14, -1.309865e-14, -1.004585e-14, -1.804299e-14, 
    -5.378532e-15, -9.852598e-15, -7.613499e-15, -2.011807e-14, 
    -8.351467e-15, -1.461984e-14, -1.833461e-14, -1.148414e-14, 
    -1.665345e-14, -8.193752e-15, -5.990749e-15, -1.883114e-14, 
    -1.044309e-14, -1.379712e-14, -2.208165e-14, -1.285503e-14, 
    -1.734834e-14, -1.284898e-14, -1.034721e-14, -5.035612e-15, 
    -1.561071e-14, -2.090988e-15, -2.443739e-15, -5.362058e-15, 
    -1.399363e-14, -1.182948e-14, -1.577987e-14, -1.494634e-14, 
    -1.200451e-14, -1.740924e-14, -1.478177e-14, -1.573175e-14, 
    -1.166343e-14, -1.092669e-14, -1.6887e-14, -1.594797e-14, -1.932333e-14, 
    -7.869626e-15, -1.182889e-14, -1.724011e-14, -1.373206e-14, 
    -1.781817e-14, -1.489905e-14, -8.081232e-15, -1.138609e-14, 
    -5.475304e-15, -1.302546e-14, -1.416642e-14, -1.414965e-14, 
    -1.199525e-14, -1.162625e-14, -1.479349e-14, -1.194572e-14, 
    -1.121486e-14, -1.193407e-14, -1.548725e-14, -1.562581e-14, 
    -8.246573e-15, -7.464023e-15, -1.194006e-14, -1.271416e-14, 
    -4.059896e-15, -1.192554e-14, -1.908284e-14, -1.27022e-14, -1.559229e-14, 
    -1.388135e-14, -1.156345e-14, -1.474368e-14, -1.496864e-14, 
    -1.265353e-14, -1.115267e-14, -1.920879e-14, -9.465302e-15, 
    -1.314363e-14, -1.09245e-14, -1.777368e-14, -1.255408e-14, -1.41414e-14, 
    -1.188004e-14, -1.58851e-14, -4.468805e-15, -1.536989e-14, -1.184827e-14, 
    -1.716859e-14, -1.680685e-14, -1.384382e-14, -1.583921e-14, 
    -1.308721e-14, -9.311751e-15, -1.448951e-14, -1.824822e-14, 
    -1.766307e-14, -1.283769e-14, -1.479284e-14, -1.011789e-14, 
    -1.627027e-14, -1.078418e-14, -1.364776e-14, -1.74615e-14, -7.379497e-15, 
    -1.819708e-14, -1.335433e-14, -1.794241e-14, 3.755253e-16, -8.732558e-15, 
    -1.449947e-14, -1.417087e-14, -1.478948e-14, -1.428588e-14, 
    -1.574871e-14, -9.026309e-15, -1.409236e-14, -1.309223e-14, 
    -1.498039e-14, -8.105934e-15, -1.84871e-14, -1.17872e-14, -9.531053e-15, 
    -1.042964e-14, -1.551181e-14, -1.759335e-14, -1.619122e-14, 
    -1.059845e-14, -1.415647e-14, -1.742397e-14, -1.151103e-14, 
    -1.204296e-14, -7.892252e-15, -1.712923e-14, -9.930629e-15, 
    -8.023749e-15, -1.244653e-14, -7.992316e-15, -1.871058e-14, 
    -9.590677e-15, -5.497096e-15, -9.314017e-15, -2.175076e-14, 
    -1.186341e-14, -1.345461e-14, -1.691409e-14, -2.044701e-14, 
    -1.116955e-14, -6.391656e-15, -8.426983e-15, -1.366767e-14, 
    -1.049668e-14, -1.637067e-14, -1.04249e-14, -1.767098e-14, -1.410203e-14, 
    -1.732808e-14, -1.229981e-14, -1.631929e-14, -1.741325e-14, -9.64665e-15, 
    -1.436283e-14, -2.573331e-14, -2.103501e-14, -1.432573e-14, 
    -1.241198e-14, -8.132364e-15, -1.23478e-14, -8.818249e-15, -6.967372e-15, 
    -1.058833e-14, -9.532313e-15, -1.67701e-14, -1.468112e-14, -1.470123e-14, 
    -6.98236e-15, -1.445864e-14, -6.228603e-15, -1.32845e-14, -1.273192e-14, 
    -1.494378e-14, -1.728911e-14, -1.006631e-14, -4.656007e-15, 
    -1.532875e-14, -1.158589e-14, -1.44792e-14, -6.341654e-15, -1.763612e-14, 
    -1.239283e-14, -1.334025e-14, -9.425975e-15, -1.603158e-14, 
    -1.674765e-14, -1.209307e-14, -1.224237e-14, -7.113998e-15, 
    -1.524367e-14, -1.523806e-14, -1.345929e-14, -6.839131e-15, 
    -1.575888e-14, -1.857821e-14, -1.68021e-14, -1.325122e-14, -1.01733e-14, 
    -6.490788e-15, -1.412503e-14, -1.584711e-14, -1.107061e-14, 
    -1.415666e-14, -1.035481e-14, -1.197011e-14, -1.147306e-14, 
    -1.482755e-14, -8.470465e-15, -1.407436e-14, -7.583732e-15, 
    -1.795312e-14, -1.105888e-14, -7.627765e-15, -1.625882e-14, 
    -8.460815e-15, -9.173724e-15, -6.86021e-15, -2.404625e-14, -5.692475e-15, 
    -1.270796e-14, -1.669822e-14, -1.428343e-14, -9.524771e-15, 
    -9.932942e-15, -1.115024e-14, -1.102507e-14, -1.331325e-14, 
    -1.694368e-14, -1.029779e-14, -2.048829e-14, -8.07185e-15, -1.022591e-14, 
    -1.911889e-14, -2.358672e-14, -1.544993e-14, -1.358969e-14, 
    -1.995404e-14, -1.178014e-14, -1.763536e-14, -1.519171e-14, -1.17405e-14, 
    -1.204197e-14, -1.266204e-14, -2.25833e-14, -1.535363e-14, -1.847866e-14, 
    -1.560926e-14, -1.122388e-14, -1.458277e-14, -1.503394e-14, 
    -4.962354e-15, -1.176647e-14, -1.252587e-14, -5.903448e-15, 
    -9.714803e-15, -2.08974e-14, -8.65237e-15, -1.076483e-14, -9.36798e-15, 
    -1.687698e-14, -1.5158e-14, -1.193936e-14, -1.503313e-14, -1.451596e-14, 
    -1.512126e-14, -9.148822e-15, -8.867466e-15, -1.840232e-14, 
    -8.367235e-15, -1.451465e-14, -6.067177e-15, -1.146112e-14, 
    -1.370285e-14, -1.467954e-14, -1.348211e-14, -1.650992e-14, 
    -2.074097e-14, -1.901881e-14, -5.734835e-15, -1.037728e-14, 
    -1.172074e-14, -1.535527e-14, -1.504782e-14, -8.638779e-15, -1.59938e-14, 
    -1.540104e-14, -6.356521e-15, -1.124811e-14, -1.269007e-14, 
    -2.151007e-14, -1.46394e-14, -1.282696e-14, -1.448593e-14, -1.152931e-14, 
    -4.606332e-15, -9.921382e-15, -8.419315e-15, -1.622662e-14, -1.710202e-14 ;

 ERRSOI =
  -4.090069e-10, -3.898483e-10, -4.426774e-10, -3.631617e-10, -3.275914e-10, 
    -2.659812e-10, -2.049339e-10, -2.853442e-10, -3.191629e-10, 
    -5.454376e-10, -3.663976e-10, -2.041492e-10, -3.567062e-10, 
    -1.940392e-10, -2.857709e-10, -1.981749e-10, -3.756453e-10, 
    -3.267113e-10, -2.548871e-10, -5.337828e-11, -3.641685e-10, 
    -2.829078e-10, -2.752846e-10, -3.705833e-10, -5.761821e-10, 
    -4.431324e-10, -2.474199e-10, -2.575608e-10, -3.623463e-10, 
    -2.181668e-10, -2.374137e-10, -2.337752e-10, -3.795294e-10, 
    -2.859855e-10, -5.106129e-10, -3.904322e-10, -1.818034e-10, 
    -1.091919e-10, -3.57283e-10, -2.472394e-10, -4.428087e-10, -3.68462e-10, 
    -2.8464e-10, -2.496582e-10, -2.218905e-10, -2.982186e-10, -1.12018e-10, 
    -1.946832e-10, -3.138196e-10, -5.511234e-10, -3.102172e-10, 
    -3.195665e-10, -2.98675e-10, -3.273972e-10, -1.920322e-10, -2.697638e-10, 
    -1.940249e-10, -1.960644e-10, -2.851906e-10, -4.704452e-10, 
    -4.540996e-10, -3.523034e-10, -3.056667e-10, -3.522986e-10, 
    -1.978839e-10, -4.723015e-10, -3.606656e-10, -2.973614e-10, 
    -3.879017e-10, -3.704048e-10, -2.987216e-10, -3.203088e-10, 
    -2.317156e-10, -4.922818e-10, -1.405869e-10, -2.601793e-10, -2.28922e-10, 
    -2.969314e-10, -2.712919e-10, -3.089227e-10, -3.706693e-10, 
    -3.568324e-10, -2.228819e-10, -4.195995e-10, -1.939456e-10, 
    -4.354856e-10, -3.966288e-10, -3.554353e-10, -4.004404e-10, 
    -4.141767e-10, -2.237782e-10, -2.970312e-10, -2.521501e-10, 
    -1.521138e-10, -1.348882e-10, -3.572693e-10, -3.059665e-10, 
    -4.331416e-10, -4.062593e-10, -4.474849e-10, -4.236446e-10, 
    -3.116747e-10, -4.532566e-10, -2.340301e-10, -3.685912e-10, 
    -1.976577e-10, -3.261841e-10, -3.013531e-10, -5.422167e-10, 
    -2.761114e-10, -3.871519e-10, -2.872281e-10, -3.546932e-10, 
    -4.049664e-10, -2.728576e-10, -3.494655e-10, -3.800174e-10, 
    -3.615168e-10, -1.885021e-10, -2.802115e-10, -2.666794e-10, 
    -3.440097e-10, -4.010284e-10, -2.429121e-10, -3.636759e-10, 
    -3.453511e-10, -4.287012e-10, -3.789999e-10, -3.890475e-10, 
    -3.126003e-10, -2.923249e-10, -4.644035e-10, -3.626139e-10, 
    -2.906828e-10, -4.087712e-10, -4.919711e-10, -4.268435e-10, 
    -2.143371e-10, -4.256277e-10, -2.64819e-10, -2.838791e-10, -2.374583e-10, 
    -3.776494e-10, -3.396826e-10, -3.839714e-10, -3.748729e-10, 
    -8.485006e-11, -2.650286e-10, -4.253197e-10, -2.787116e-10, 
    -2.684041e-10, -4.999602e-10, -4.038682e-10, -4.902626e-10, -3.55029e-10, 
    -3.486751e-10, -3.10243e-10, -4.214645e-10, -3.041278e-10, -3.530393e-10, 
    -2.767842e-10, -2.602485e-10, -4.471512e-10, -5.043579e-10, 
    -2.993119e-10, -4.036277e-10, -3.129637e-10, -4.329972e-10, 
    -3.129838e-10, -4.88828e-10, -1.763373e-10, -1.141654e-10, -3.7828e-10, 
    -4.38879e-10, -5.989764e-10, -1.306704e-10, -2.340363e-10, -3.309834e-10, 
    -2.771022e-10, -4.499786e-10, -5.771132e-10, -3.083215e-10, 
    -3.551021e-10, -3.641022e-10, -5.844025e-11, -3.223224e-10, 
    -3.176466e-10, -3.597219e-10, -4.171445e-10, -2.75516e-10, -2.664545e-10, 
    -3.950567e-10, -2.054976e-10, -1.923893e-10, -3.905596e-10, 
    -1.001603e-10, -2.190681e-10, -2.602136e-10, -2.801806e-10, 
    -3.533365e-10, -1.081927e-10, -3.279868e-10, -1.722972e-10, 
    -1.956542e-10, -4.556584e-10, -1.718141e-10, -2.513737e-10, 
    -4.761144e-10, -6.312376e-10, -1.940842e-10, -3.571246e-10, 
    -2.482719e-10, -4.709845e-10, -3.864384e-10, -2.676226e-10, 
    -2.666569e-10, -3.22581e-10, -3.624568e-10, -5.337827e-10, -1.839091e-10, 
    -7.587932e-11, -3.691848e-10, -2.877073e-10, -1.950624e-10, 
    -5.608478e-11, -3.740228e-10, -4.960943e-10, -2.710089e-10, 
    -4.314908e-10, -4.153904e-10, -6.358768e-11, -3.620816e-10, 
    -3.437907e-10, -2.231277e-10, -3.057277e-10, -4.183598e-10, 
    -2.690554e-10, -2.996225e-10, -3.836582e-10, -1.899995e-10, 
    -3.493895e-10, -4.678412e-10, -3.510833e-10, -3.513087e-10, 
    -3.373541e-10, -3.136235e-10, -3.325386e-10, -2.136128e-10, 
    -2.185538e-10, -1.862316e-10, -2.851678e-10, -5.239081e-10, 
    -3.915134e-10, -4.334493e-10, -2.444754e-10, -3.110148e-10, 
    -3.358647e-10, -4.017692e-10, -4.816988e-10, -4.382316e-10, 
    -3.284251e-10, -3.487875e-10, -6.44148e-10, -3.154539e-10, -3.066484e-10, 
    -2.765405e-10, -2.223551e-10, -4.066589e-10, -4.169383e-10, 
    -2.053551e-10, -3.204523e-10, -3.77725e-10, -2.627865e-10, -1.89181e-10, 
    -2.428815e-10, -1.601074e-10, -3.869128e-10, -2.246953e-10, 
    -2.177774e-10, -2.199507e-10, -4.157559e-10, -1.634023e-10, 
    -3.877103e-10, -2.093354e-10, -2.588384e-10, -3.000407e-10, 
    -4.251172e-10, -3.031199e-10, -4.147943e-10, -1.536809e-10, 
    -1.366941e-10, -3.141805e-10, -3.322523e-10, -4.098754e-10, 
    -5.315617e-10, -3.554208e-10, -3.179737e-10, -4.207278e-10, 
    -4.028863e-10, -2.253652e-10, -4.617216e-10, -4.81746e-10, -4.166097e-10, 
    -3.024842e-10, -2.611551e-10, -2.220818e-10, -3.736496e-10, 
    -2.991805e-10, -1.116245e-10, -2.379295e-10, -3.464306e-10, 
    -2.854753e-10, -4.241995e-10, -4.729001e-10, -3.399801e-10, 
    -1.336642e-10, -3.448125e-10, -1.2169e-10, -2.604267e-10, -2.667301e-10, 
    -3.050781e-10, -3.275528e-10, -2.271237e-10, -5.28892e-10, -3.47892e-10, 
    -9.287026e-11, -3.736881e-10, -3.857443e-10, -2.660092e-10, 
    -3.677911e-10, -2.883584e-10, -4.932516e-10, -3.474866e-10, 
    -2.697228e-10, -2.593776e-10, -3.861699e-10, -4.427788e-10, -3.631815e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4 =
  5.810961e-16, 5.748851e-16, 5.760943e-16, 5.710734e-16, 5.738605e-16, 
    5.705704e-16, 5.798389e-16, 5.746377e-16, 5.779598e-16, 5.805384e-16, 
    5.61294e-16, 5.708493e-16, 5.513279e-16, 5.574545e-16, 5.420333e-16, 
    5.522817e-16, 5.399614e-16, 5.423308e-16, 5.351949e-16, 5.372416e-16, 
    5.26468e-16, 5.342496e-16, 5.217193e-16, 5.279392e-16, 5.269666e-16, 
    5.344525e-16, 5.689309e-16, 5.624856e-16, 5.693119e-16, 5.683942e-16, 
    5.688063e-16, 5.738026e-16, 5.763151e-16, 5.815708e-16, 5.806178e-16, 
    5.767577e-16, 5.679814e-16, 5.709655e-16, 5.634392e-16, 5.636094e-16, 
    5.55199e-16, 5.589952e-16, 5.448113e-16, 5.488522e-16, 5.371562e-16, 
    5.401031e-16, 5.372945e-16, 5.381466e-16, 5.372834e-16, 5.416039e-16, 
    5.397537e-16, 5.435523e-16, 5.582845e-16, 5.539647e-16, 5.668223e-16, 
    5.745145e-16, 5.796108e-16, 5.832188e-16, 5.827091e-16, 5.817369e-16, 
    5.76735e-16, 5.720222e-16, 5.684232e-16, 5.660121e-16, 5.636339e-16, 
    5.564162e-16, 5.525888e-16, 5.439927e-16, 5.455475e-16, 5.429138e-16, 
    5.403961e-16, 5.361617e-16, 5.368593e-16, 5.349916e-16, 5.42984e-16, 
    5.37675e-16, 5.464323e-16, 5.440404e-16, 5.62983e-16, 5.70161e-16, 
    5.732013e-16, 5.758618e-16, 5.82317e-16, 5.778611e-16, 5.796187e-16, 
    5.754355e-16, 5.727726e-16, 5.740902e-16, 5.659461e-16, 5.691159e-16, 
    5.523617e-16, 5.595944e-16, 5.406899e-16, 5.452285e-16, 5.396008e-16, 
    5.424745e-16, 5.375481e-16, 5.419822e-16, 5.342965e-16, 5.309936e-16, 
    5.337654e-16, 5.277381e-16, 5.422277e-16, 5.372941e-16, 5.741269e-16, 
    5.739121e-16, 5.729112e-16, 5.773071e-16, 5.775759e-16, 5.815968e-16, 
    5.780197e-16, 5.764943e-16, 5.726184e-16, 5.703217e-16, 5.681363e-16, 
    5.633236e-16, 5.579351e-16, 5.503787e-16, 5.449346e-16, 5.412776e-16, 
    5.43521e-16, 5.415404e-16, 5.437542e-16, 5.447912e-16, 5.316221e-16, 
    5.397362e-16, 5.283713e-16, 5.289109e-16, 5.34947e-16, 5.2885e-16, 
    5.737613e-16, 5.749974e-16, 5.792822e-16, 5.759297e-16, 5.820342e-16, 
    5.786189e-16, 5.766523e-16, 5.690489e-16, 5.673756e-16, 5.658216e-16, 
    5.627499e-16, 5.58801e-16, 5.518559e-16, 5.457958e-16, 5.402497e-16, 
    5.406566e-16, 5.405133e-16, 5.392723e-16, 5.423447e-16, 5.387675e-16, 
    5.381662e-16, 5.397374e-16, 5.289831e-16, 5.315935e-16, 5.289223e-16, 
    5.306219e-16, 5.745958e-16, 5.725152e-16, 5.736396e-16, 5.715244e-16, 
    5.730145e-16, 5.663795e-16, 5.643861e-16, 5.55035e-16, 5.588786e-16, 
    5.527593e-16, 5.582581e-16, 5.572845e-16, 5.525578e-16, 5.579616e-16, 
    5.461296e-16, 5.541567e-16, 5.39224e-16, 5.472634e-16, 5.387192e-16, 
    5.402737e-16, 5.376997e-16, 5.353916e-16, 5.308596e-16, 5.254937e-16, 
    5.267371e-16, 5.222453e-16, 5.6941e-16, 5.667039e-16, 5.66943e-16, 
    5.641083e-16, 5.620092e-16, 5.574534e-16, 5.501257e-16, 5.528843e-16, 
    5.47818e-16, 5.467993e-16, 5.544956e-16, 5.497727e-16, 5.648915e-16, 
    5.624552e-16, 5.639066e-16, 5.691962e-16, 5.522479e-16, 5.609621e-16, 
    5.448443e-16, 5.495854e-16, 5.357207e-16, 5.426258e-16, 5.274212e-16, 
    5.215992e-16, 5.161114e-16, 5.096799e-16, 5.652264e-16, 5.670666e-16, 
    5.637711e-16, 5.592017e-16, 5.549556e-16, 5.492964e-16, 5.48717e-16, 
    5.476547e-16, 5.449016e-16, 5.425839e-16, 5.47318e-16, 5.420025e-16, 
    5.618884e-16, 5.514902e-16, 5.677613e-16, 5.628737e-16, 5.594717e-16, 
    5.609655e-16, 5.531995e-16, 5.513649e-16, 5.438937e-16, 5.477595e-16, 
    5.230367e-16, 5.349027e-16, 5.047744e-16, 5.127691e-16, 5.677091e-16, 
    5.652331e-16, 5.565921e-16, 5.607079e-16, 5.489185e-16, 5.460065e-16, 
    5.436371e-16, 5.406034e-16, 5.402762e-16, 5.384766e-16, 5.414246e-16, 
    5.385934e-16, 5.492843e-16, 5.445132e-16, 5.575824e-16, 5.544082e-16, 
    5.558693e-16, 5.574703e-16, 5.525252e-16, 5.472433e-16, 5.471316e-16, 
    5.45435e-16, 5.406449e-16, 5.488706e-16, 5.217108e-16, 5.391313e-16, 
    5.625297e-16, 5.577447e-16, 5.570618e-16, 5.58917e-16, 5.462986e-16, 
    5.508789e-16, 5.385207e-16, 5.418676e-16, 5.363814e-16, 5.391092e-16, 
    5.395101e-16, 5.430085e-16, 5.451833e-16, 5.506689e-16, 5.551225e-16, 
    5.586482e-16, 5.57829e-16, 5.539543e-16, 5.469201e-16, 5.402459e-16, 
    5.417094e-16, 5.367989e-16, 5.497754e-16, 5.443427e-16, 5.464436e-16, 
    5.409614e-16, 5.529573e-16, 5.427427e-16, 5.555603e-16, 5.544397e-16, 
    5.509697e-16, 5.439729e-16, 5.424236e-16, 5.407662e-16, 5.417893e-16, 
    5.467415e-16, 5.475523e-16, 5.510544e-16, 5.520198e-16, 5.546838e-16, 
    5.568863e-16, 5.548738e-16, 5.527579e-16, 5.467399e-16, 5.413018e-16, 
    5.353585e-16, 5.339022e-16, 5.253137e-16, 5.309808e-16, 5.216224e-16, 
    5.295781e-16, 5.157934e-16, 5.42151e-16, 5.298137e-16, 5.508121e-16, 
    5.487332e-16, 5.449667e-16, 5.363067e-16, 5.409872e-16, 5.35513e-16, 
    5.475841e-16, 5.538199e-16, 5.554318e-16, 5.584338e-16, 5.553632e-16, 
    5.556131e-16, 5.526711e-16, 5.53617e-16, 5.465398e-16, 5.503443e-16, 
    5.395199e-16, 5.355566e-16, 5.227159e-16, 5.158206e-16, 5.087843e-16, 
    5.056713e-16, 5.047231e-16, 5.043265e-16 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGR =
  -384.5455, -385.5921, -385.3889, -386.2325, -385.7648, -386.317, -384.758, 
    -385.6335, -385.0748, -384.6401, -387.8684, -386.2702, -389.53, 
    -388.5111, -391.0797, -389.3712, -391.4224, -391.0312, -392.2097, 
    -391.8722, -393.5343, -392.3654, -394.3158, -393.2928, -393.4526, 
    -392.332, -386.5925, -387.6693, -386.5286, -386.6822, -386.6134, 
    -385.7742, -385.3509, -384.4659, -384.6267, -385.2769, -386.7513, 
    -386.2513, -387.5124, -387.4839, -388.8869, -388.2544, -390.6118, 
    -389.9422, -391.8863, -391.3996, -391.8633, -391.7228, -391.8651, 
    -391.1514, -391.4572, -390.8204, -388.3728, -389.0921, -386.9457, 
    -385.6534, -384.7963, -384.1875, -384.2735, -384.4375, -385.2807, 
    -386.0738, -386.6779, -387.0818, -387.4798, -388.6827, -389.3205, 
    -390.7469, -390.4901, -390.9256, -391.3512, -392.0501, -391.9352, 
    -392.2429, -390.9145, -391.8002, -390.3436, -390.7396, -387.586, 
    -386.3862, -385.8744, -385.4279, -384.3397, -385.0911, -384.7948, -385.5, 
    -385.9477, -385.7263, -387.0928, -386.5616, -389.3582, -388.154, 
    -391.3026, -390.5428, -391.4827, -390.9989, -391.8213, -391.0891, 
    -392.3575, -392.7894, -392.4449, -393.3264, -391.0485, -391.8631, 
    -385.7201, -385.7561, -385.9245, -385.1844, -385.1392, -384.4614, 
    -385.0647, -385.3214, -385.9738, -386.3593, -386.7257, -387.5314, 
    -388.4307, -389.6881, -390.5915, -391.2057, -390.8258, -391.1622, 
    -390.7871, -390.6155, -392.6857, -391.4599, -393.222, -393.1332, 
    -392.2501, -393.1432, -385.7815, -385.5738, -384.8518, -385.4168, 
    -384.3876, -384.9635, -385.2944, -386.5722, -386.8534, -387.1135, 
    -387.6275, -388.2868, -389.4428, -390.4485, -391.3756, -391.3083, 
    -391.332, -391.5368, -391.0291, -391.6202, -391.7192, -391.4601, 
    -393.1213, -392.6909, -393.1313, -392.8512, -385.6414, -385.991, 
    -385.802, -386.1572, -385.9068, -387.0194, -387.3529, -388.9135, 
    -388.2737, -389.2925, -388.3774, -388.5394, -389.3249, -388.427, 
    -390.3927, -389.0594, -391.5448, -390.2042, -391.6282, -391.3716, 
    -391.7966, -392.177, -392.8119, -393.6954, -393.491, -394.2298, 
    -386.5123, -386.9655, -386.9259, -387.4004, -387.7511, -388.5116, 
    -389.7305, -389.2723, -390.1138, -390.2826, -389.0044, -389.7888, 
    -387.269, -387.6758, -387.4339, -386.5478, -389.3774, -387.9254, 
    -390.6064, -389.8203, -392.1227, -390.9731, -393.3783, -394.3348, 
    -395.2363, -396.2871, -387.2131, -386.9052, -387.4569, -388.2193, 
    -388.9275, -389.8682, -389.9646, -390.1407, -390.5972, -390.9807, 
    -390.196, -391.0858, -387.7694, -389.5035, -386.7885, -387.6058, 
    -388.1745, -387.9254, -389.2201, -389.525, -390.7635, -390.1235, 
    -394.0984, -392.2568, -397.0881, -395.7825, -386.7975, -387.2123, 
    -388.6546, -387.9685, -389.9312, -390.4139, -390.8066, -391.3167, 
    -391.3711, -391.6681, -391.1814, -391.649, -389.8702, -390.6613, 
    -388.4903, -389.0186, -388.7757, -388.5089, -389.3321, -390.2083, 
    -390.2276, -390.5083, -391.3071, -389.9391, -394.3147, -391.5576, 
    -387.6644, -388.4621, -388.5768, -388.2677, -390.3655, -389.6055, 
    -391.6609, -391.1081, -392.014, -391.5638, -391.4976, -390.9105, 
    -390.5503, -389.6402, -388.8996, -388.3126, -388.4492, -389.094, 
    -390.262, -391.3758, -391.1337, -391.9452, -389.7889, -390.6892, 
    -390.3411, -391.2578, -389.26, -390.9518, -388.8272, -389.0137, 
    -389.5904, -390.7498, -391.0161, -391.2898, -391.1211, -390.2917, 
    -390.1576, -389.5765, -389.4158, -388.9731, -388.6063, -388.9413, 
    -389.2929, -390.2923, -391.2012, -392.1823, -392.4226, -393.7236, 
    -392.7905, -394.329, -393.0198, -395.2861, -391.0597, -392.9826, 
    -389.6169, -389.962, -390.5855, -392.0252, -391.2535, -392.1563, 
    -390.1524, -389.1159, -388.8485, -388.3482, -388.8599, -388.8183, 
    -389.3079, -389.1506, -390.3255, -389.6945, -391.4958, -392.1494, 
    -394.1521, -395.283, -396.4345, -396.9423, -397.0969, -397.1614 ;

 FGR12 =
  -50.01731, -50.0848, -50.0717, -50.12616, -50.09598, -50.13163, -50.03103, 
    -50.08744, -50.05144, -50.02344, -50.23201, -50.12862, -50.34003, 
    -50.27389, -50.44043, -50.3297, -50.46284, -50.43734, -50.51439, 
    -50.49231, -50.59677, -50.5246, -50.64814, -50.58098, -50.59143, 
    -50.5224, -50.14949, -50.21909, -50.14534, -50.15527, -50.15083, 
    -50.09657, -50.06918, -50.01223, -50.02258, -50.06445, -50.15973, 
    -50.12742, -50.2091, -50.20726, -50.29829, -50.25726, -50.41056, 
    -50.36694, -50.49323, -50.46141, -50.49172, -50.48254, -50.49184, 
    -50.44519, -50.46516, -50.42418, -50.26492, -50.3116, -50.17233, 
    -50.0887, -50.03348, -49.9943, -49.99983, -50.01037, -50.0647, -50.11594, 
    -50.15503, -50.18118, -50.207, -50.28493, -50.32642, -50.41933, 
    -50.40264, -50.43101, -50.45825, -50.50393, -50.49642, -50.51654, 
    -50.43032, -50.48756, -50.3931, -50.4189, -50.21368, -50.13615, 
    -50.10297, -50.07421, -50.00409, -50.05247, -50.03338, -50.07888, 
    -50.1078, -50.09351, -50.1819, -50.1475, -50.32887, -50.25071, -50.45506, 
    -50.40607, -50.46683, -50.43584, -50.48895, -50.44114, -50.52406, 
    -50.54799, -50.52977, -50.58321, -50.43848, -50.49168, -50.0931, 
    -50.09542, -50.10629, -50.05849, -50.05557, -50.01193, -50.0508, 
    -50.06734, -50.1095, -50.1344, -50.15812, -50.21031, -50.26865, 
    -50.35035, -50.40924, -50.44874, -50.42454, -50.4459, -50.42201, 
    -50.41083, -50.54119, -50.46533, -50.57637, -50.57055, -50.51702, 
    -50.5712, -50.09706, -50.08366, -50.03707, -50.07352, -50.00718, 
    -50.04425, -50.06558, -50.14814, -50.16639, -50.18322, -50.21656, 
    -50.25935, -50.33441, -50.39989, -50.45984, -50.45545, -50.457, 
    -50.47037, -50.43721, -50.47581, -50.48228, -50.46536, -50.56977, 
    -50.54158, -50.57042, -50.55208, -50.08802, -50.11059, -50.09839, 
    -50.12133, -50.10515, -50.17708, -50.1987, -50.29996, -50.2585, 
    -50.32462, -50.26523, -50.27573, -50.32664, -50.26846, -50.39622, 
    -50.30943, -50.47088, -50.3839, -50.47634, -50.45958, -50.48737, 
    -50.51224, -50.5495, -50.60739, -50.594, -50.64252, -50.14431, -50.17361, 
    -50.17109, -50.20182, -50.22456, -50.27394, -50.35313, -50.32336, 
    -50.37811, -50.3891, -50.30595, -50.35691, -50.19329, -50.21963, 
    -50.20398, -50.14659, -50.33012, -50.23584, -50.4102, -50.35899, 
    -50.50868, -50.4341, -50.58661, -50.64935, -50.70879, -50.77805, 
    -50.18968, -50.16975, -50.20551, -50.25491, -50.30094, -50.36209, 
    -50.3684, -50.37986, -50.40963, -50.43465, -50.38343, -50.44091, 
    -50.22564, -50.33834, -50.16217, -50.21507, -50.25203, -50.23588, 
    -50.31997, -50.33979, -50.42043, -50.37875, -50.63379, -50.51741, 
    -50.83107, -50.74475, -50.16278, -50.18964, -50.28319, -50.23868, 
    -50.36622, -50.39765, -50.42329, -50.45597, -50.45955, -50.47894, 
    -50.44716, -50.4777, -50.36223, -50.41379, -50.27257, -50.30685, 
    -50.2911, -50.27378, -50.32726, -50.3842, -50.38553, -50.4038, -50.45515, 
    -50.36675, -50.6479, -50.47157, -50.21896, -50.27066, -50.27816, 
    -50.25813, -50.3945, -50.34501, -50.47848, -50.44238, -50.50158, 
    -50.47214, -50.4678, -50.43007, -50.40655, -50.34726, -50.29911, 
    -50.26105, -50.26991, -50.31174, -50.38773, -50.45982, -50.44401, 
    -50.49708, -50.35696, -50.4156, -50.39289, -50.45214, -50.32255, 
    -50.43257, -50.29445, -50.30655, -50.34403, -50.4195, -50.43637, 
    -50.45421, -50.44321, -50.38968, -50.38095, -50.34314, -50.33266, 
    -50.30392, -50.2801, -50.30184, -50.32467, -50.38973, -50.44843, 
    -50.51257, -50.52834, -50.60915, -50.54801, -50.64883, -50.56291, 
    -50.71191, -50.43911, -50.56055, -50.34577, -50.36823, -50.40881, 
    -50.50223, -50.45186, -50.51083, -50.38061, -50.31314, -50.29582, 
    -50.26335, -50.29656, -50.29387, -50.32568, -50.31546, -50.3919, 
    -50.35082, -50.46767, -50.5104, -50.6374, -50.7118, -50.78786, -50.82145, 
    -50.83168, -50.83596 ;

 FGR_R =
  -384.5455, -385.5921, -385.3889, -386.2325, -385.7648, -386.317, -384.758, 
    -385.6335, -385.0748, -384.6401, -387.8684, -386.2702, -389.53, 
    -388.5111, -391.0797, -389.3712, -391.4224, -391.0312, -392.2097, 
    -391.8722, -393.5343, -392.3654, -394.3158, -393.2928, -393.4526, 
    -392.332, -386.5925, -387.6693, -386.5286, -386.6822, -386.6134, 
    -385.7742, -385.3509, -384.4659, -384.6267, -385.2769, -386.7513, 
    -386.2513, -387.5124, -387.4839, -388.8869, -388.2544, -390.6118, 
    -389.9422, -391.8863, -391.3996, -391.8633, -391.7228, -391.8651, 
    -391.1514, -391.4572, -390.8204, -388.3728, -389.0921, -386.9457, 
    -385.6534, -384.7963, -384.1875, -384.2735, -384.4375, -385.2807, 
    -386.0738, -386.6779, -387.0818, -387.4798, -388.6827, -389.3205, 
    -390.7469, -390.4901, -390.9256, -391.3512, -392.0501, -391.9352, 
    -392.2429, -390.9145, -391.8002, -390.3436, -390.7396, -387.586, 
    -386.3862, -385.8744, -385.4279, -384.3397, -385.0911, -384.7948, -385.5, 
    -385.9477, -385.7263, -387.0928, -386.5616, -389.3582, -388.154, 
    -391.3026, -390.5428, -391.4827, -390.9989, -391.8213, -391.0891, 
    -392.3575, -392.7894, -392.4449, -393.3264, -391.0485, -391.8631, 
    -385.7201, -385.7561, -385.9245, -385.1844, -385.1392, -384.4614, 
    -385.0647, -385.3214, -385.9738, -386.3593, -386.7257, -387.5314, 
    -388.4307, -389.6881, -390.5915, -391.2057, -390.8258, -391.1622, 
    -390.7871, -390.6155, -392.6857, -391.4599, -393.222, -393.1332, 
    -392.2501, -393.1432, -385.7815, -385.5738, -384.8518, -385.4168, 
    -384.3876, -384.9635, -385.2944, -386.5722, -386.8534, -387.1135, 
    -387.6275, -388.2868, -389.4428, -390.4485, -391.3756, -391.3083, 
    -391.332, -391.5368, -391.0291, -391.6202, -391.7192, -391.4601, 
    -393.1213, -392.6909, -393.1313, -392.8512, -385.6414, -385.991, 
    -385.802, -386.1572, -385.9068, -387.0194, -387.3529, -388.9135, 
    -388.2737, -389.2925, -388.3774, -388.5394, -389.3249, -388.427, 
    -390.3927, -389.0594, -391.5448, -390.2042, -391.6282, -391.3716, 
    -391.7966, -392.177, -392.8119, -393.6954, -393.491, -394.2298, 
    -386.5123, -386.9655, -386.9259, -387.4004, -387.7511, -388.5116, 
    -389.7305, -389.2723, -390.1138, -390.2826, -389.0044, -389.7888, 
    -387.269, -387.6758, -387.4339, -386.5478, -389.3774, -387.9254, 
    -390.6064, -389.8203, -392.1227, -390.9731, -393.3783, -394.3348, 
    -395.2363, -396.2871, -387.2131, -386.9052, -387.4569, -388.2193, 
    -388.9275, -389.8682, -389.9646, -390.1407, -390.5972, -390.9807, 
    -390.196, -391.0858, -387.7694, -389.5035, -386.7885, -387.6058, 
    -388.1745, -387.9254, -389.2201, -389.525, -390.7635, -390.1235, 
    -394.0984, -392.2568, -397.0881, -395.7825, -386.7975, -387.2123, 
    -388.6546, -387.9685, -389.9312, -390.4139, -390.8066, -391.3167, 
    -391.3711, -391.6681, -391.1814, -391.649, -389.8702, -390.6613, 
    -388.4903, -389.0186, -388.7757, -388.5089, -389.3321, -390.2083, 
    -390.2276, -390.5083, -391.3071, -389.9391, -394.3147, -391.5576, 
    -387.6644, -388.4621, -388.5768, -388.2677, -390.3655, -389.6055, 
    -391.6609, -391.1081, -392.014, -391.5638, -391.4976, -390.9105, 
    -390.5503, -389.6402, -388.8996, -388.3126, -388.4492, -389.094, 
    -390.262, -391.3758, -391.1337, -391.9452, -389.7889, -390.6892, 
    -390.3411, -391.2578, -389.26, -390.9518, -388.8272, -389.0137, 
    -389.5904, -390.7498, -391.0161, -391.2898, -391.1211, -390.2917, 
    -390.1576, -389.5765, -389.4158, -388.9731, -388.6063, -388.9413, 
    -389.2929, -390.2923, -391.2012, -392.1823, -392.4226, -393.7236, 
    -392.7905, -394.329, -393.0198, -395.2861, -391.0597, -392.9826, 
    -389.6169, -389.962, -390.5855, -392.0252, -391.2535, -392.1563, 
    -390.1524, -389.1159, -388.8485, -388.3482, -388.8599, -388.8183, 
    -389.3079, -389.1506, -390.3255, -389.6945, -391.4958, -392.1494, 
    -394.1521, -395.283, -396.4345, -396.9423, -397.0969, -397.1614 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  47.78409, 47.8606, 47.84574, 47.90741, 47.87322, 47.91359, 47.79963, 
    47.86362, 47.82278, 47.79101, 48.02697, 47.91017, 48.14847, 48.07399, 
    48.26083, 48.13685, 48.28588, 48.2573, 48.34346, 48.31878, 48.41801, 
    48.35485, 48.47505, 48.40039, 48.41205, 48.3524, 47.93373, 48.01242, 
    47.92906, 47.94028, 47.93526, 47.87391, 47.84295, 47.77828, 47.79003, 
    47.83755, 47.94533, 47.90879, 48.00098, 47.99891, 48.10147, 48.05523, 
    48.22758, 48.17862, 48.31981, 48.28423, 48.31813, 48.30786, 48.31827, 
    48.26608, 48.28844, 48.24282, 48.06388, 48.11647, 47.95955, 47.86507, 
    47.80243, 47.75792, 47.76421, 47.7762, 47.83783, 47.89581, 47.93998, 
    47.96951, 47.9986, 48.08652, 48.13315, 48.23745, 48.21868, 48.25051, 
    48.28069, 48.33178, 48.32338, 48.34588, 48.24971, 48.31351, 48.20797, 
    48.23692, 48.00632, 47.91866, 47.88122, 47.84859, 47.76905, 47.82397, 
    47.80232, 47.85387, 47.8866, 47.87042, 47.97031, 47.93147, 48.13592, 
    48.04788, 48.27714, 48.22253, 48.2903, 48.25588, 48.31505, 48.26153, 
    48.35427, 48.36369, 48.36065, 48.40285, 48.25856, 48.31812, 47.86996, 
    47.87259, 47.8849, 47.83079, 47.82749, 47.77795, 47.82205, 47.84081, 
    47.88851, 47.91668, 47.94347, 48.00237, 48.0681, 48.16004, 48.22609, 
    48.27005, 48.24322, 48.26688, 48.24039, 48.22785, 48.35614, 48.28864, 
    48.39524, 48.38876, 48.34641, 48.38949, 47.87445, 47.85926, 47.80648, 
    47.84779, 47.77255, 47.81465, 47.83883, 47.93224, 47.95281, 47.97182, 
    48.0094, 48.05759, 48.14211, 48.21564, 48.28247, 48.27756, 48.27929, 
    48.29426, 48.25714, 48.30036, 48.30759, 48.28865, 48.38789, 48.35652, 
    48.38862, 48.3682, 47.8642, 47.88976, 47.87595, 47.90191, 47.88361, 
    47.96494, 47.98932, 48.1034, 48.05664, 48.13111, 48.06422, 48.07606, 
    48.13346, 48.06784, 48.21154, 48.11406, 48.29485, 48.19775, 48.30094, 
    48.28218, 48.31326, 48.34106, 48.36533, 48.42977, 48.41486, 48.46878, 
    47.92787, 47.96099, 47.95811, 47.99279, 48.01843, 48.07403, 48.16314, 
    48.12965, 48.19117, 48.2035, 48.11006, 48.1674, 47.98318, 48.01292, 
    47.99524, 47.93047, 48.13731, 48.03116, 48.22717, 48.16971, 48.3371, 
    48.25398, 48.40664, 48.47643, 48.54226, 48.61898, 47.9791, 47.9566, 
    47.99693, 48.05265, 48.10443, 48.17321, 48.18026, 48.19313, 48.22651, 
    48.25455, 48.19717, 48.26129, 48.01974, 48.14655, 47.94806, 48.0078, 
    48.04938, 48.03117, 48.12583, 48.14812, 48.23866, 48.19188, 48.45918, 
    48.34689, 48.67749, 48.58213, 47.94873, 47.97905, 48.08448, 48.03432, 
    48.17781, 48.2131, 48.24182, 48.27816, 48.28215, 48.30386, 48.26828, 
    48.30247, 48.17335, 48.2312, 48.07247, 48.1111, 48.09334, 48.07384, 
    48.13402, 48.19806, 48.19949, 48.22001, 48.27743, 48.1784, 48.47494, 
    48.29574, 48.0121, 48.0704, 48.07879, 48.0562, 48.20956, 48.154, 
    48.30334, 48.26292, 48.32915, 48.29624, 48.29139, 48.24942, 48.22308, 
    48.15654, 48.1024, 48.05948, 48.06947, 48.1166, 48.20199, 48.28248, 
    48.26478, 48.32412, 48.16741, 48.23323, 48.20778, 48.27386, 48.12875, 
    48.2524, 48.0971, 48.11074, 48.1529, 48.23766, 48.2562, 48.2762, 
    48.26387, 48.20417, 48.19436, 48.15189, 48.14013, 48.10777, 48.08096, 
    48.10544, 48.13115, 48.20422, 48.26972, 48.34145, 48.35902, 48.43182, 
    48.36376, 48.47599, 48.38046, 48.54587, 48.25936, 48.37776, 48.15483, 
    48.18007, 48.22564, 48.32996, 48.27355, 48.33954, 48.19398, 48.1182, 
    48.09866, 48.06208, 48.0995, 48.09646, 48.13225, 48.12075, 48.20664, 
    48.16051, 48.29126, 48.33904, 48.46311, 48.54566, 48.62976, 48.66684, 
    48.67813, 48.68285 ;

 FIRA_R =
  47.78409, 47.8606, 47.84574, 47.90741, 47.87322, 47.91359, 47.79963, 
    47.86362, 47.82278, 47.79101, 48.02697, 47.91017, 48.14847, 48.07399, 
    48.26083, 48.13685, 48.28588, 48.2573, 48.34346, 48.31878, 48.41801, 
    48.35485, 48.47505, 48.40039, 48.41205, 48.3524, 47.93373, 48.01242, 
    47.92906, 47.94028, 47.93526, 47.87391, 47.84295, 47.77828, 47.79003, 
    47.83755, 47.94533, 47.90879, 48.00098, 47.99891, 48.10147, 48.05523, 
    48.22758, 48.17862, 48.31981, 48.28423, 48.31813, 48.30786, 48.31827, 
    48.26608, 48.28844, 48.24282, 48.06388, 48.11647, 47.95955, 47.86507, 
    47.80243, 47.75792, 47.76421, 47.7762, 47.83783, 47.89581, 47.93998, 
    47.96951, 47.9986, 48.08652, 48.13315, 48.23745, 48.21868, 48.25051, 
    48.28069, 48.33178, 48.32338, 48.34588, 48.24971, 48.31351, 48.20797, 
    48.23692, 48.00632, 47.91866, 47.88122, 47.84859, 47.76905, 47.82397, 
    47.80232, 47.85387, 47.8866, 47.87042, 47.97031, 47.93147, 48.13592, 
    48.04788, 48.27714, 48.22253, 48.2903, 48.25588, 48.31505, 48.26153, 
    48.35427, 48.36369, 48.36065, 48.40285, 48.25856, 48.31812, 47.86996, 
    47.87259, 47.8849, 47.83079, 47.82749, 47.77795, 47.82205, 47.84081, 
    47.88851, 47.91668, 47.94347, 48.00237, 48.0681, 48.16004, 48.22609, 
    48.27005, 48.24322, 48.26688, 48.24039, 48.22785, 48.35614, 48.28864, 
    48.39524, 48.38876, 48.34641, 48.38949, 47.87445, 47.85926, 47.80648, 
    47.84779, 47.77255, 47.81465, 47.83883, 47.93224, 47.95281, 47.97182, 
    48.0094, 48.05759, 48.14211, 48.21564, 48.28247, 48.27756, 48.27929, 
    48.29426, 48.25714, 48.30036, 48.30759, 48.28865, 48.38789, 48.35652, 
    48.38862, 48.3682, 47.8642, 47.88976, 47.87595, 47.90191, 47.88361, 
    47.96494, 47.98932, 48.1034, 48.05664, 48.13111, 48.06422, 48.07606, 
    48.13346, 48.06784, 48.21154, 48.11406, 48.29485, 48.19775, 48.30094, 
    48.28218, 48.31326, 48.34106, 48.36533, 48.42977, 48.41486, 48.46878, 
    47.92787, 47.96099, 47.95811, 47.99279, 48.01843, 48.07403, 48.16314, 
    48.12965, 48.19117, 48.2035, 48.11006, 48.1674, 47.98318, 48.01292, 
    47.99524, 47.93047, 48.13731, 48.03116, 48.22717, 48.16971, 48.3371, 
    48.25398, 48.40664, 48.47643, 48.54226, 48.61898, 47.9791, 47.9566, 
    47.99693, 48.05265, 48.10443, 48.17321, 48.18026, 48.19313, 48.22651, 
    48.25455, 48.19717, 48.26129, 48.01974, 48.14655, 47.94806, 48.0078, 
    48.04938, 48.03117, 48.12583, 48.14812, 48.23866, 48.19188, 48.45918, 
    48.34689, 48.67749, 48.58213, 47.94873, 47.97905, 48.08448, 48.03432, 
    48.17781, 48.2131, 48.24182, 48.27816, 48.28215, 48.30386, 48.26828, 
    48.30247, 48.17335, 48.2312, 48.07247, 48.1111, 48.09334, 48.07384, 
    48.13402, 48.19806, 48.19949, 48.22001, 48.27743, 48.1784, 48.47494, 
    48.29574, 48.0121, 48.0704, 48.07879, 48.0562, 48.20956, 48.154, 
    48.30334, 48.26292, 48.32915, 48.29624, 48.29139, 48.24942, 48.22308, 
    48.15654, 48.1024, 48.05948, 48.06947, 48.1166, 48.20199, 48.28248, 
    48.26478, 48.32412, 48.16741, 48.23323, 48.20778, 48.27386, 48.12875, 
    48.2524, 48.0971, 48.11074, 48.1529, 48.23766, 48.2562, 48.2762, 
    48.26387, 48.20417, 48.19436, 48.15189, 48.14013, 48.10777, 48.08096, 
    48.10544, 48.13115, 48.20422, 48.26972, 48.34145, 48.35902, 48.43182, 
    48.36376, 48.47599, 48.38046, 48.54587, 48.25936, 48.37776, 48.15483, 
    48.18007, 48.22564, 48.32996, 48.27355, 48.33954, 48.19398, 48.1182, 
    48.09866, 48.06208, 48.0995, 48.09646, 48.13225, 48.12075, 48.20664, 
    48.16051, 48.29126, 48.33904, 48.46311, 48.54566, 48.62976, 48.66684, 
    48.67813, 48.68285 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  262.1302, 262.2068, 262.1919, 262.2535, 262.2194, 262.2597, 262.1458, 
    262.2097, 262.1689, 262.1371, 262.3731, 262.2563, 262.4946, 262.4201, 
    262.607, 262.483, 262.632, 262.6035, 262.6896, 262.6649, 262.7642, 
    262.701, 262.8212, 262.7466, 262.7582, 262.6985, 262.2799, 262.3586, 
    262.2752, 262.2864, 262.2814, 262.2201, 262.1891, 262.1244, 262.1362, 
    262.1837, 262.2915, 262.2549, 262.3471, 262.3451, 262.4476, 262.4014, 
    262.5737, 262.5247, 262.666, 262.6304, 262.6643, 262.654, 262.6644, 
    262.6122, 262.6346, 262.589, 262.41, 262.4626, 262.3057, 262.2112, 
    262.1486, 262.1041, 262.1104, 262.1223, 262.184, 262.2419, 262.2861, 
    262.3156, 262.3448, 262.4326, 262.4793, 262.5836, 262.5648, 262.5966, 
    262.6268, 262.6779, 262.6695, 262.692, 262.5959, 262.6597, 262.5541, 
    262.5831, 262.3525, 262.2648, 262.2274, 262.1947, 262.1152, 262.1701, 
    262.1485, 262.2, 262.2327, 262.2166, 262.3165, 262.2776, 262.4821, 
    262.394, 262.6233, 262.5687, 262.6364, 262.602, 262.6612, 262.6077, 
    262.7004, 262.7098, 262.7068, 262.749, 262.6047, 262.6642, 262.2161, 
    262.2188, 262.231, 262.1769, 262.1736, 262.1241, 262.1682, 262.187, 
    262.2346, 262.2628, 262.2896, 262.3485, 262.4142, 262.5062, 262.5722, 
    262.6162, 262.5894, 262.613, 262.5865, 262.574, 262.7023, 262.6348, 
    262.7414, 262.7349, 262.6925, 262.7356, 262.2206, 262.2054, 262.1526, 
    262.1939, 262.1187, 262.1608, 262.185, 262.2784, 262.299, 262.318, 
    262.3555, 262.4037, 262.4883, 262.5618, 262.6286, 262.6237, 262.6254, 
    262.6404, 262.6033, 262.6465, 262.6537, 262.6348, 262.734, 262.7027, 
    262.7348, 262.7144, 262.2104, 262.2359, 262.2221, 262.248, 262.2297, 
    262.3111, 262.3354, 262.4496, 262.4028, 262.4773, 262.4104, 262.4222, 
    262.4796, 262.414, 262.5577, 262.4602, 262.641, 262.5439, 262.6471, 
    262.6283, 262.6594, 262.6872, 262.7115, 262.7759, 262.761, 262.8149, 
    262.274, 262.3071, 262.3043, 262.3389, 262.3646, 262.4202, 262.5093, 
    262.4758, 262.5373, 262.5497, 262.4562, 262.5135, 262.3293, 262.3591, 
    262.3414, 262.2766, 262.4835, 262.3773, 262.5733, 262.5158, 262.6832, 
    262.6001, 262.7528, 262.8226, 262.8884, 262.9651, 262.3253, 262.3027, 
    262.3431, 262.3988, 262.4506, 262.5193, 262.5264, 262.5393, 262.5727, 
    262.6007, 262.5433, 262.6074, 262.3659, 262.4927, 262.2942, 262.3539, 
    262.3955, 262.3773, 262.472, 262.4943, 262.5848, 262.538, 262.8053, 
    262.693, 263.0236, 262.9283, 262.2949, 262.3252, 262.4306, 262.3805, 
    262.524, 262.5592, 262.588, 262.6243, 262.6283, 262.65, 262.6144, 
    262.6486, 262.5195, 262.5773, 262.4186, 262.4572, 262.4395, 262.42, 
    262.4802, 262.5442, 262.5456, 262.5662, 262.6236, 262.5245, 262.8211, 
    262.6419, 262.3582, 262.4165, 262.4249, 262.4023, 262.5557, 262.5002, 
    262.6495, 262.6091, 262.6753, 262.6424, 262.6375, 262.5956, 262.5692, 
    262.5027, 262.4485, 262.4056, 262.4156, 262.4627, 262.5481, 262.6286, 
    262.6109, 262.6703, 262.5135, 262.5794, 262.5539, 262.62, 262.4749, 
    262.5985, 262.4432, 262.4569, 262.4991, 262.5838, 262.6023, 262.6223, 
    262.61, 262.5503, 262.5405, 262.498, 262.4863, 262.4539, 262.4271, 
    262.4516, 262.4773, 262.5504, 262.6159, 262.6876, 262.7052, 262.778, 
    262.7099, 262.8221, 262.7266, 262.892, 262.6055, 262.7239, 262.501, 
    262.5262, 262.5718, 262.6761, 262.6197, 262.6857, 262.5401, 262.4644, 
    262.4448, 262.4082, 262.4456, 262.4426, 262.4784, 262.4669, 262.5528, 
    262.5067, 262.6374, 262.6852, 262.8093, 262.8918, 262.9759, 263.013, 
    263.0243, 263.029 ;

 FIRE_R =
  262.1302, 262.2068, 262.1919, 262.2535, 262.2194, 262.2597, 262.1458, 
    262.2097, 262.1689, 262.1371, 262.3731, 262.2563, 262.4946, 262.4201, 
    262.607, 262.483, 262.632, 262.6035, 262.6896, 262.6649, 262.7642, 
    262.701, 262.8212, 262.7466, 262.7582, 262.6985, 262.2799, 262.3586, 
    262.2752, 262.2864, 262.2814, 262.2201, 262.1891, 262.1244, 262.1362, 
    262.1837, 262.2915, 262.2549, 262.3471, 262.3451, 262.4476, 262.4014, 
    262.5737, 262.5247, 262.666, 262.6304, 262.6643, 262.654, 262.6644, 
    262.6122, 262.6346, 262.589, 262.41, 262.4626, 262.3057, 262.2112, 
    262.1486, 262.1041, 262.1104, 262.1223, 262.184, 262.2419, 262.2861, 
    262.3156, 262.3448, 262.4326, 262.4793, 262.5836, 262.5648, 262.5966, 
    262.6268, 262.6779, 262.6695, 262.692, 262.5959, 262.6597, 262.5541, 
    262.5831, 262.3525, 262.2648, 262.2274, 262.1947, 262.1152, 262.1701, 
    262.1485, 262.2, 262.2327, 262.2166, 262.3165, 262.2776, 262.4821, 
    262.394, 262.6233, 262.5687, 262.6364, 262.602, 262.6612, 262.6077, 
    262.7004, 262.7098, 262.7068, 262.749, 262.6047, 262.6642, 262.2161, 
    262.2188, 262.231, 262.1769, 262.1736, 262.1241, 262.1682, 262.187, 
    262.2346, 262.2628, 262.2896, 262.3485, 262.4142, 262.5062, 262.5722, 
    262.6162, 262.5894, 262.613, 262.5865, 262.574, 262.7023, 262.6348, 
    262.7414, 262.7349, 262.6925, 262.7356, 262.2206, 262.2054, 262.1526, 
    262.1939, 262.1187, 262.1608, 262.185, 262.2784, 262.299, 262.318, 
    262.3555, 262.4037, 262.4883, 262.5618, 262.6286, 262.6237, 262.6254, 
    262.6404, 262.6033, 262.6465, 262.6537, 262.6348, 262.734, 262.7027, 
    262.7348, 262.7144, 262.2104, 262.2359, 262.2221, 262.248, 262.2297, 
    262.3111, 262.3354, 262.4496, 262.4028, 262.4773, 262.4104, 262.4222, 
    262.4796, 262.414, 262.5577, 262.4602, 262.641, 262.5439, 262.6471, 
    262.6283, 262.6594, 262.6872, 262.7115, 262.7759, 262.761, 262.8149, 
    262.274, 262.3071, 262.3043, 262.3389, 262.3646, 262.4202, 262.5093, 
    262.4758, 262.5373, 262.5497, 262.4562, 262.5135, 262.3293, 262.3591, 
    262.3414, 262.2766, 262.4835, 262.3773, 262.5733, 262.5158, 262.6832, 
    262.6001, 262.7528, 262.8226, 262.8884, 262.9651, 262.3253, 262.3027, 
    262.3431, 262.3988, 262.4506, 262.5193, 262.5264, 262.5393, 262.5727, 
    262.6007, 262.5433, 262.6074, 262.3659, 262.4927, 262.2942, 262.3539, 
    262.3955, 262.3773, 262.472, 262.4943, 262.5848, 262.538, 262.8053, 
    262.693, 263.0236, 262.9283, 262.2949, 262.3252, 262.4306, 262.3805, 
    262.524, 262.5592, 262.588, 262.6243, 262.6283, 262.65, 262.6144, 
    262.6486, 262.5195, 262.5773, 262.4186, 262.4572, 262.4395, 262.42, 
    262.4802, 262.5442, 262.5456, 262.5662, 262.6236, 262.5245, 262.8211, 
    262.6419, 262.3582, 262.4165, 262.4249, 262.4023, 262.5557, 262.5002, 
    262.6495, 262.6091, 262.6753, 262.6424, 262.6375, 262.5956, 262.5692, 
    262.5027, 262.4485, 262.4056, 262.4156, 262.4627, 262.5481, 262.6286, 
    262.6109, 262.6703, 262.5135, 262.5794, 262.5539, 262.62, 262.4749, 
    262.5985, 262.4432, 262.4569, 262.4991, 262.5838, 262.6023, 262.6223, 
    262.61, 262.5503, 262.5405, 262.498, 262.4863, 262.4539, 262.4271, 
    262.4516, 262.4773, 262.5504, 262.6159, 262.6876, 262.7052, 262.778, 
    262.7099, 262.8221, 262.7266, 262.892, 262.6055, 262.7239, 262.501, 
    262.5262, 262.5718, 262.6761, 262.6197, 262.6857, 262.5401, 262.4644, 
    262.4448, 262.4082, 262.4456, 262.4426, 262.4784, 262.4669, 262.5528, 
    262.5067, 262.6374, 262.6852, 262.8093, 262.8918, 262.9759, 263.013, 
    263.0243, 263.029 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSAT =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FSA_R =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347 ;

 FSDSND =
  0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532 ;

 FSDSNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSDSNI =
  0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819 ;

 FSDSVD =
  0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128 ;

 FSDSVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSDSVI =
  0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223 ;

 FSDSVILN =
  0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376 ;

 FSH =
  336.8137, 337.7838, 337.5954, 338.3774, 337.9438, 338.4557, 337.0107, 
    337.8221, 337.3043, 336.9014, 339.8937, 338.4124, 341.4338, 340.4894, 
    342.8711, 341.2866, 343.1888, 342.8262, 343.9185, 343.6057, 345.1686, 
    344.0629, 345.893, 344.9447, 345.0929, 344.0319, 338.7111, 339.7091, 
    338.6518, 338.7942, 338.7304, 337.9526, 337.5602, 336.7399, 336.8889, 
    337.4916, 338.8582, 338.3947, 339.5637, 339.5373, 340.8377, 340.2515, 
    342.4366, 341.8159, 343.6188, 343.1677, 343.5975, 343.4672, 343.5992, 
    342.9376, 343.2211, 342.6299, 340.3612, 341.028, 339.0385, 337.8406, 
    337.0461, 336.4818, 336.5616, 336.7136, 337.4951, 338.2303, 338.7902, 
    339.1646, 339.5335, 340.6485, 341.2396, 342.5618, 342.3237, 342.7274, 
    343.1228, 343.7706, 343.6641, 343.9493, 342.7171, 343.539, 342.188, 
    342.555, 339.6319, 338.5199, 338.0454, 337.6316, 336.6229, 337.3194, 
    337.0448, 337.6984, 338.1134, 337.9082, 339.1748, 338.6824, 341.2746, 
    340.1584, 343.0778, 342.3726, 343.2447, 342.7953, 343.5585, 342.8799, 
    344.0556, 344.478, 344.1365, 344.9758, 342.8422, 343.5973, 337.9024, 
    337.9358, 338.0919, 337.4059, 337.364, 336.7357, 337.2949, 337.5329, 
    338.1376, 338.4948, 338.8346, 339.5814, 340.4149, 341.5804, 342.4177, 
    342.9879, 342.6349, 342.9476, 342.599, 342.44, 344.3819, 343.2236, 
    344.8791, 344.7968, 343.956, 344.806, 337.9594, 337.7668, 337.0976, 
    337.6213, 336.6673, 337.2011, 337.5079, 338.6923, 338.9529, 339.1939, 
    339.6704, 340.2815, 341.353, 342.2852, 343.1454, 343.0831, 343.105, 
    343.2949, 342.8242, 343.3721, 343.4639, 343.2237, 344.7857, 344.3867, 
    344.795, 344.5353, 337.8294, 338.1535, 337.9784, 338.3076, 338.0755, 
    339.1068, 339.4159, 340.8624, 340.2693, 341.2137, 340.3654, 340.5157, 
    341.2437, 340.4114, 342.2335, 340.9976, 343.3022, 342.0587, 343.3795, 
    343.1417, 343.5357, 343.8882, 344.4989, 345.3179, 345.1284, 345.8133, 
    338.6367, 339.0567, 339.0201, 339.4599, 339.785, 340.4899, 341.6196, 
    341.195, 341.9749, 342.1313, 340.9466, 341.6737, 339.3381, 339.7152, 
    339.4909, 338.6696, 341.2924, 339.9465, 342.4315, 341.7029, 343.8379, 
    342.7714, 345.024, 345.9106, 346.7463, 347.7204, 339.2863, 339.0009, 
    339.5123, 340.2189, 340.8754, 341.7473, 341.8366, 341.9998, 342.423, 
    342.7785, 342.0511, 342.8768, 339.802, 341.4093, 338.8927, 339.6503, 
    340.1774, 339.9465, 341.1465, 341.4291, 342.5771, 341.9839, 345.6915, 
    343.9622, 348.4629, 347.2527, 338.9011, 339.2855, 340.6224, 339.9865, 
    341.8056, 342.2531, 342.617, 343.0908, 343.1413, 343.4165, 342.9654, 
    343.3989, 341.7491, 342.4824, 340.4701, 340.9598, 340.7346, 340.4874, 
    341.2504, 342.0625, 342.0804, 342.3406, 343.082, 341.813, 345.892, 
    343.3141, 339.7046, 340.444, 340.5503, 340.2638, 342.2082, 341.5038, 
    343.4099, 342.8975, 343.7372, 343.3199, 343.2585, 342.7134, 342.3795, 
    341.5359, 340.8495, 340.3054, 340.432, 341.0297, 342.1123, 343.1456, 
    342.9212, 343.6734, 341.6738, 342.5083, 342.1856, 343.0362, 341.1836, 
    342.7517, 340.7824, 340.9552, 341.4898, 342.5645, 342.8122, 343.0659, 
    342.9095, 342.1399, 342.0155, 341.4769, 341.3279, 340.9176, 340.5776, 
    340.8881, 341.2141, 342.1404, 342.9838, 343.8932, 344.1159, 345.3441, 
    344.479, 345.9053, 344.6917, 346.7925, 342.8526, 344.6571, 341.5143, 
    341.8342, 342.4121, 343.7476, 343.0323, 343.869, 342.0107, 341.05, 
    340.8021, 340.3384, 340.8127, 340.7742, 341.228, 341.0822, 342.1712, 
    341.5863, 343.2568, 343.8626, 345.7413, 346.7896, 347.857, 348.3277, 
    348.471, 348.5309 ;

 FSH_G =
  343.5179, 344.4886, 344.3001, 345.0825, 344.6487, 345.1609, 343.715, 
    344.5269, 344.0088, 343.6057, 346.5996, 345.1175, 348.1406, 347.1957, 
    349.5787, 347.9933, 349.8965, 349.5338, 350.6267, 350.3137, 351.8773, 
    350.7711, 352.6022, 351.6533, 351.8016, 350.7401, 345.4164, 346.4149, 
    345.357, 345.4995, 345.4357, 344.6575, 344.2648, 343.4441, 343.5932, 
    344.1962, 345.5636, 345.0999, 346.2695, 346.2431, 347.5442, 346.9576, 
    349.1439, 348.5229, 350.3268, 349.8754, 350.3055, 350.1751, 350.3072, 
    349.6452, 349.9288, 349.3373, 347.0674, 347.7345, 345.7439, 344.5454, 
    343.7505, 343.1859, 343.2657, 343.4178, 344.1998, 344.9353, 345.4955, 
    345.8701, 346.2393, 347.3548, 347.9463, 349.2692, 349.031, 349.4349, 
    349.8306, 350.4787, 350.3721, 350.6574, 349.4246, 350.2469, 348.8952, 
    349.2624, 346.3377, 345.2251, 344.7504, 344.3362, 343.3271, 344.0239, 
    343.7492, 344.4031, 344.8183, 344.6131, 345.8804, 345.3877, 347.9813, 
    346.8645, 349.7855, 349.0799, 349.9524, 349.5028, 350.2664, 349.5875, 
    350.7638, 351.1864, 350.8448, 351.6845, 349.5498, 350.3053, 344.6072, 
    344.6407, 344.7968, 344.1104, 344.0685, 343.4399, 343.9995, 344.2375, 
    344.8426, 345.2, 345.5399, 346.2871, 347.1211, 348.2872, 349.125, 
    349.6956, 349.3423, 349.6552, 349.3064, 349.1473, 351.0902, 349.9314, 
    351.5877, 351.5053, 350.6642, 351.5146, 344.6642, 344.4716, 343.802, 
    344.326, 343.3715, 343.9056, 344.2125, 345.3976, 345.6583, 345.8995, 
    346.3762, 346.9876, 348.0597, 348.9925, 349.8531, 349.7908, 349.8127, 
    350.0027, 349.5318, 350.08, 350.1718, 349.9315, 351.4943, 351.095, 
    351.5035, 351.2437, 344.5342, 344.8585, 344.6833, 345.0127, 344.7805, 
    345.8123, 346.1216, 347.5689, 346.9755, 347.9203, 347.0717, 347.222, 
    347.9503, 347.1176, 348.9407, 347.7041, 350.0101, 348.7658, 350.0874, 
    349.8494, 350.2436, 350.5964, 351.2072, 352.0268, 351.8372, 352.5224, 
    345.3419, 345.7622, 345.7256, 346.1656, 346.4908, 347.1962, 348.3265, 
    347.9016, 348.682, 348.8385, 347.6531, 348.3806, 346.0437, 346.4211, 
    346.1967, 345.3749, 347.9991, 346.6525, 349.1388, 348.4098, 350.5461, 
    349.4789, 351.7327, 352.6198, 353.456, 354.4306, 345.9919, 345.7064, 
    346.218, 346.925, 347.5818, 348.4542, 348.5437, 348.7069, 349.1303, 
    349.486, 348.7582, 349.5844, 346.5078, 348.1161, 345.5981, 346.3561, 
    346.8835, 346.6525, 347.8531, 348.1359, 349.2845, 348.691, 352.4006, 
    350.6704, 355.1735, 353.9626, 345.6065, 345.9911, 347.3288, 346.6925, 
    348.5126, 348.9603, 349.3245, 349.7985, 349.849, 350.1244, 349.673, 
    350.1067, 348.4561, 349.1898, 347.1763, 347.6663, 347.4411, 347.1937, 
    347.9571, 348.7696, 348.7875, 349.0479, 349.7896, 348.52, 352.6012, 
    350.0219, 346.4104, 347.1502, 347.2566, 346.9699, 348.9154, 348.2106, 
    350.1178, 349.6051, 350.4453, 350.0277, 349.9663, 349.4209, 349.0869, 
    348.2428, 347.556, 347.0116, 347.1382, 347.7362, 348.8194, 349.8533, 
    349.6288, 350.3814, 348.3807, 349.2157, 348.8928, 349.7439, 347.8902, 
    349.4592, 347.4888, 347.6617, 348.1966, 349.2719, 349.5198, 349.7736, 
    349.6171, 348.847, 348.7226, 348.1837, 348.0346, 347.6241, 347.2839, 
    347.5946, 347.9207, 348.8476, 349.6914, 350.6013, 350.8242, 352.0529, 
    351.1874, 352.6145, 351.4001, 353.5021, 349.5602, 351.3656, 348.2211, 
    348.5412, 349.1195, 350.4556, 349.7399, 350.5772, 348.7178, 347.7566, 
    347.5086, 347.0446, 347.5192, 347.4806, 347.9346, 347.7888, 348.8784, 
    348.2932, 349.9646, 350.5707, 352.4504, 353.4993, 354.5673, 355.0383, 
    355.1816, 355.2415 ;

 FSH_NODYNLNDUSE =
  336.8137, 337.7838, 337.5954, 338.3774, 337.9438, 338.4557, 337.0107, 
    337.8221, 337.3043, 336.9014, 339.8937, 338.4124, 341.4338, 340.4894, 
    342.8711, 341.2866, 343.1888, 342.8262, 343.9185, 343.6057, 345.1686, 
    344.0629, 345.893, 344.9447, 345.0929, 344.0319, 338.7111, 339.7091, 
    338.6518, 338.7942, 338.7304, 337.9526, 337.5602, 336.7399, 336.8889, 
    337.4916, 338.8582, 338.3947, 339.5637, 339.5373, 340.8377, 340.2515, 
    342.4366, 341.8159, 343.6188, 343.1677, 343.5975, 343.4672, 343.5992, 
    342.9376, 343.2211, 342.6299, 340.3612, 341.028, 339.0385, 337.8406, 
    337.0461, 336.4818, 336.5616, 336.7136, 337.4951, 338.2303, 338.7902, 
    339.1646, 339.5335, 340.6485, 341.2396, 342.5618, 342.3237, 342.7274, 
    343.1228, 343.7706, 343.6641, 343.9493, 342.7171, 343.539, 342.188, 
    342.555, 339.6319, 338.5199, 338.0454, 337.6316, 336.6229, 337.3194, 
    337.0448, 337.6984, 338.1134, 337.9082, 339.1748, 338.6824, 341.2746, 
    340.1584, 343.0778, 342.3726, 343.2447, 342.7953, 343.5585, 342.8799, 
    344.0556, 344.478, 344.1365, 344.9758, 342.8422, 343.5973, 337.9024, 
    337.9358, 338.0919, 337.4059, 337.364, 336.7357, 337.2949, 337.5329, 
    338.1376, 338.4948, 338.8346, 339.5814, 340.4149, 341.5804, 342.4177, 
    342.9879, 342.6349, 342.9476, 342.599, 342.44, 344.3819, 343.2236, 
    344.8791, 344.7968, 343.956, 344.806, 337.9594, 337.7668, 337.0976, 
    337.6213, 336.6673, 337.2011, 337.5079, 338.6923, 338.9529, 339.1939, 
    339.6704, 340.2815, 341.353, 342.2852, 343.1454, 343.0831, 343.105, 
    343.2949, 342.8242, 343.3721, 343.4639, 343.2237, 344.7857, 344.3867, 
    344.795, 344.5353, 337.8294, 338.1535, 337.9784, 338.3076, 338.0755, 
    339.1068, 339.4159, 340.8624, 340.2693, 341.2137, 340.3654, 340.5157, 
    341.2437, 340.4114, 342.2335, 340.9976, 343.3022, 342.0587, 343.3795, 
    343.1417, 343.5357, 343.8882, 344.4989, 345.3179, 345.1284, 345.8133, 
    338.6367, 339.0567, 339.0201, 339.4599, 339.785, 340.4899, 341.6196, 
    341.195, 341.9749, 342.1313, 340.9466, 341.6737, 339.3381, 339.7152, 
    339.4909, 338.6696, 341.2924, 339.9465, 342.4315, 341.7029, 343.8379, 
    342.7714, 345.024, 345.9106, 346.7463, 347.7204, 339.2863, 339.0009, 
    339.5123, 340.2189, 340.8754, 341.7473, 341.8366, 341.9998, 342.423, 
    342.7785, 342.0511, 342.8768, 339.802, 341.4093, 338.8927, 339.6503, 
    340.1774, 339.9465, 341.1465, 341.4291, 342.5771, 341.9839, 345.6915, 
    343.9622, 348.4629, 347.2527, 338.9011, 339.2855, 340.6224, 339.9865, 
    341.8056, 342.2531, 342.617, 343.0908, 343.1413, 343.4165, 342.9654, 
    343.3989, 341.7491, 342.4824, 340.4701, 340.9598, 340.7346, 340.4874, 
    341.2504, 342.0625, 342.0804, 342.3406, 343.082, 341.813, 345.892, 
    343.3141, 339.7046, 340.444, 340.5503, 340.2638, 342.2082, 341.5038, 
    343.4099, 342.8975, 343.7372, 343.3199, 343.2585, 342.7134, 342.3795, 
    341.5359, 340.8495, 340.3054, 340.432, 341.0297, 342.1123, 343.1456, 
    342.9212, 343.6734, 341.6738, 342.5083, 342.1856, 343.0362, 341.1836, 
    342.7517, 340.7824, 340.9552, 341.4898, 342.5645, 342.8122, 343.0659, 
    342.9095, 342.1399, 342.0155, 341.4769, 341.3279, 340.9176, 340.5776, 
    340.8881, 341.2141, 342.1404, 342.9838, 343.8932, 344.1159, 345.3441, 
    344.479, 345.9053, 344.6917, 346.7925, 342.8526, 344.6571, 341.5143, 
    341.8342, 342.4121, 343.7476, 343.0323, 343.869, 342.0107, 341.05, 
    340.8021, 340.3384, 340.8127, 340.7742, 341.228, 341.0822, 342.1712, 
    341.5863, 343.2568, 343.8626, 345.7413, 346.7896, 347.857, 348.3277, 
    348.471, 348.5309 ;

 FSH_R =
  336.8137, 337.7838, 337.5954, 338.3774, 337.9438, 338.4557, 337.0107, 
    337.8221, 337.3043, 336.9014, 339.8937, 338.4124, 341.4338, 340.4894, 
    342.8711, 341.2866, 343.1888, 342.8262, 343.9185, 343.6057, 345.1686, 
    344.0629, 345.893, 344.9447, 345.0929, 344.0319, 338.7111, 339.7091, 
    338.6518, 338.7942, 338.7304, 337.9526, 337.5602, 336.7399, 336.8889, 
    337.4916, 338.8582, 338.3947, 339.5637, 339.5373, 340.8377, 340.2515, 
    342.4366, 341.8159, 343.6188, 343.1677, 343.5975, 343.4672, 343.5992, 
    342.9376, 343.2211, 342.6299, 340.3612, 341.028, 339.0385, 337.8406, 
    337.0461, 336.4818, 336.5616, 336.7136, 337.4951, 338.2303, 338.7902, 
    339.1646, 339.5335, 340.6485, 341.2396, 342.5618, 342.3237, 342.7274, 
    343.1228, 343.7706, 343.6641, 343.9493, 342.7171, 343.539, 342.188, 
    342.555, 339.6319, 338.5199, 338.0454, 337.6316, 336.6229, 337.3194, 
    337.0448, 337.6984, 338.1134, 337.9082, 339.1748, 338.6824, 341.2746, 
    340.1584, 343.0778, 342.3726, 343.2447, 342.7953, 343.5585, 342.8799, 
    344.0556, 344.478, 344.1365, 344.9758, 342.8422, 343.5973, 337.9024, 
    337.9358, 338.0919, 337.4059, 337.364, 336.7357, 337.2949, 337.5329, 
    338.1376, 338.4948, 338.8346, 339.5814, 340.4149, 341.5804, 342.4177, 
    342.9879, 342.6349, 342.9476, 342.599, 342.44, 344.3819, 343.2236, 
    344.8791, 344.7968, 343.956, 344.806, 337.9594, 337.7668, 337.0976, 
    337.6213, 336.6673, 337.2011, 337.5079, 338.6923, 338.9529, 339.1939, 
    339.6704, 340.2815, 341.353, 342.2852, 343.1454, 343.0831, 343.105, 
    343.2949, 342.8242, 343.3721, 343.4639, 343.2237, 344.7857, 344.3867, 
    344.795, 344.5353, 337.8294, 338.1535, 337.9784, 338.3076, 338.0755, 
    339.1068, 339.4159, 340.8624, 340.2693, 341.2137, 340.3654, 340.5157, 
    341.2437, 340.4114, 342.2335, 340.9976, 343.3022, 342.0587, 343.3795, 
    343.1417, 343.5357, 343.8882, 344.4989, 345.3179, 345.1284, 345.8133, 
    338.6367, 339.0567, 339.0201, 339.4599, 339.785, 340.4899, 341.6196, 
    341.195, 341.9749, 342.1313, 340.9466, 341.6737, 339.3381, 339.7152, 
    339.4909, 338.6696, 341.2924, 339.9465, 342.4315, 341.7029, 343.8379, 
    342.7714, 345.024, 345.9106, 346.7463, 347.7204, 339.2863, 339.0009, 
    339.5123, 340.2189, 340.8754, 341.7473, 341.8366, 341.9998, 342.423, 
    342.7785, 342.0511, 342.8768, 339.802, 341.4093, 338.8927, 339.6503, 
    340.1774, 339.9465, 341.1465, 341.4291, 342.5771, 341.9839, 345.6915, 
    343.9622, 348.4629, 347.2527, 338.9011, 339.2855, 340.6224, 339.9865, 
    341.8056, 342.2531, 342.617, 343.0908, 343.1413, 343.4165, 342.9654, 
    343.3989, 341.7491, 342.4824, 340.4701, 340.9598, 340.7346, 340.4874, 
    341.2504, 342.0625, 342.0804, 342.3406, 343.082, 341.813, 345.892, 
    343.3141, 339.7046, 340.444, 340.5503, 340.2638, 342.2082, 341.5038, 
    343.4099, 342.8975, 343.7372, 343.3199, 343.2585, 342.7134, 342.3795, 
    341.5359, 340.8495, 340.3054, 340.432, 341.0297, 342.1123, 343.1456, 
    342.9212, 343.6734, 341.6738, 342.5083, 342.1856, 343.0362, 341.1836, 
    342.7517, 340.7824, 340.9552, 341.4898, 342.5645, 342.8122, 343.0659, 
    342.9095, 342.1399, 342.0155, 341.4769, 341.3279, 340.9176, 340.5776, 
    340.8881, 341.2141, 342.1404, 342.9838, 343.8932, 344.1159, 345.3441, 
    344.479, 345.9053, 344.6917, 346.7925, 342.8526, 344.6571, 341.5143, 
    341.8342, 342.4121, 343.7476, 343.0323, 343.869, 342.0107, 341.05, 
    340.8021, 340.3384, 340.8127, 340.7742, 341.228, 341.0822, 342.1712, 
    341.5863, 343.2568, 343.8626, 345.7413, 346.7896, 347.857, 348.3277, 
    348.471, 348.5309 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -6.704242, -6.704774, -6.704673, -6.705097, -6.704865, -6.70514, -6.704355, 
    -6.704791, -6.704515, -6.704297, -6.705907, -6.705117, -6.706776, 
    -6.706263, -6.707569, -6.70669, -6.707748, -6.707554, -6.708166, 
    -6.707991, -6.708751, -6.708246, -6.709165, -6.708636, -6.708715, 
    -6.708228, -6.705286, -6.705805, -6.705253, -6.705328, -6.705297, 
    -6.704867, -6.704643, -6.704209, -6.70429, -6.704613, -6.705361, 
    -6.705114, -6.705758, -6.705744, -6.706456, -6.706134, -6.707342, 
    -6.707001, -6.707998, -6.707746, -6.707985, -6.707913, -6.707986, 
    -6.707616, -6.707774, -6.707451, -6.706192, -6.706558, -6.705463, 
    -6.704791, -6.704372, -6.704067, -6.70411, -6.70419, -6.704615, 
    -6.705024, -6.705333, -6.705538, -6.705742, -6.706332, -6.706668, 
    -6.707406, -6.707282, -6.7075, -6.707721, -6.70808, -6.708022, -6.708179, 
    -6.7075, -6.707948, -6.707209, -6.70741, -6.705761, -6.705183, -6.704906, 
    -6.704691, -6.704143, -6.704519, -6.70437, -6.704733, -6.704959, 
    -6.704849, -6.705544, -6.705272, -6.706688, -6.706078, -6.707695, 
    -6.707308, -6.707789, -6.707545, -6.70796, -6.707587, -6.70824, 
    -6.708377, -6.708282, -6.708661, -6.707566, -6.707981, -6.704844, 
    -6.704862, -6.704949, -6.704566, -6.704545, -6.704205, -6.70451, 
    -6.704638, -6.704975, -6.705168, -6.705354, -6.705764, -6.706217, 
    -6.706862, -6.707333, -6.707647, -6.707457, -6.707625, -6.707436, 
    -6.707349, -6.708323, -6.707773, -6.708606, -6.708561, -6.708181, 
    -6.708566, -6.704875, -6.704772, -6.704401, -6.704691, -6.704169, 
    -6.704456, -6.704619, -6.705269, -6.705421, -6.705551, -6.705815, 
    -6.706151, -6.706738, -6.707256, -6.707736, -6.707701, -6.707713, 
    -6.707816, -6.707555, -6.70786, -6.707907, -6.707777, -6.708555, 
    -6.708333, -6.70856, -6.708416, -6.704806, -6.704982, -6.704886, 
    -6.705064, -6.704936, -6.705495, -6.705663, -6.70646, -6.706142, 
    -6.706659, -6.706197, -6.706277, -6.706661, -6.706225, -6.70722, 
    -6.706531, -6.70782, -6.707115, -6.707863, -6.707733, -6.707952, 
    -6.708146, -6.708395, -6.708845, -6.708742, -6.709125, -6.705247, 
    -6.705472, -6.705459, -6.705699, -6.705876, -6.706267, -6.706889, 
    -6.706657, -6.70709, -6.707174, -6.706521, -6.706915, -6.705628, 
    -6.705828, -6.705714, -6.705261, -6.706701, -6.705956, -6.707339, 
    -6.706936, -6.708117, -6.707522, -6.708684, -6.709165, -6.709651, 
    -6.710182, -6.705602, -6.705449, -6.70573, -6.706107, -6.706478, 
    -6.70696, -6.707013, -6.707101, -6.707339, -6.707535, -6.707122, 
    -6.707586, -6.705861, -6.706769, -6.705384, -6.705791, -6.706088, 
    -6.705965, -6.706632, -6.706788, -6.707417, -6.707095, -6.70904, 
    -6.708177, -6.710611, -6.709923, -6.705393, -6.705605, -6.706334, 
    -6.705988, -6.706995, -6.707241, -6.707447, -6.7077, -6.707732, 
    -6.707882, -6.707635, -6.707875, -6.706961, -6.70737, -6.706258, 
    -6.706524, -6.706404, -6.706267, -6.706689, -6.707127, -6.707148, 
    -6.707286, -6.707659, -6.707, -6.709131, -6.707793, -6.705835, -6.706229, 
    -6.706299, -6.706144, -6.707216, -6.706826, -6.70788, -6.707597, 
    -6.708064, -6.707831, -6.707796, -6.7075, -6.707312, -6.706841, 
    -6.706462, -6.706168, -6.706237, -6.706561, -6.707157, -6.70773, 
    -6.707603, -6.708029, -6.706922, -6.707379, -6.707199, -6.707673, 
    -6.706648, -6.707486, -6.706431, -6.706525, -6.706818, -6.707403, 
    -6.70755, -6.707685, -6.707604, -6.707174, -6.707108, -6.706813, 
    -6.706727, -6.706506, -6.706317, -6.706487, -6.706662, -6.707179, 
    -6.707639, -6.708147, -6.708275, -6.708841, -6.708364, -6.709136, 
    -6.708457, -6.709646, -6.707551, -6.708459, -6.706835, -6.707012, 
    -6.707321, -6.708055, -6.70767, -6.708126, -6.707107, -6.706567, 
    -6.706441, -6.706183, -6.706447, -6.706426, -6.706677, -6.706597, 
    -6.707196, -6.706874, -6.707792, -6.708125, -6.709081, -6.709662, 
    -6.710274, -6.710539, -6.71062, -6.710654 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179 ;

 FSRND =
  0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234 ;

 FSRNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSRNI =
  0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666 ;

 FSRVD =
  0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223 ;

 FSRVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSRVI =
  0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_DENIT_vr =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_NIT =
  2.317337e-14, 2.33729e-14, 2.333404e-14, 2.349548e-14, 2.340585e-14, 
    2.351166e-14, 2.321374e-14, 2.338082e-14, 2.327409e-14, 2.319128e-14, 
    2.38104e-14, 2.350267e-14, 2.413232e-14, 2.393442e-14, 2.443319e-14, 
    2.410146e-14, 2.450036e-14, 2.442359e-14, 2.465506e-14, 2.458863e-14, 
    2.488593e-14, 2.468574e-14, 2.504078e-14, 2.483805e-14, 2.48697e-14, 
    2.467914e-14, 2.356446e-14, 2.377199e-14, 2.355219e-14, 2.358172e-14, 
    2.356846e-14, 2.340769e-14, 2.332688e-14, 2.315814e-14, 2.318872e-14, 
    2.331268e-14, 2.359498e-14, 2.349895e-14, 2.374136e-14, 2.373588e-14, 
    2.400724e-14, 2.388469e-14, 2.434323e-14, 2.421244e-14, 2.459139e-14, 
    2.449579e-14, 2.458689e-14, 2.455925e-14, 2.458724e-14, 2.444712e-14, 
    2.45071e-14, 2.438399e-14, 2.390765e-14, 2.404714e-14, 2.363234e-14, 
    2.338473e-14, 2.322104e-14, 2.310525e-14, 2.312159e-14, 2.315278e-14, 
    2.33134e-14, 2.346495e-14, 2.358079e-14, 2.365844e-14, 2.373508e-14, 
    2.396784e-14, 2.409154e-14, 2.436971e-14, 2.431939e-14, 2.440466e-14, 
    2.448629e-14, 2.462364e-14, 2.460101e-14, 2.466161e-14, 2.44024e-14, 
    2.457451e-14, 2.429073e-14, 2.436817e-14, 2.375593e-14, 2.352485e-14, 
    2.342696e-14, 2.334148e-14, 2.313417e-14, 2.327722e-14, 2.322077e-14, 
    2.335519e-14, 2.344081e-14, 2.339844e-14, 2.366056e-14, 2.355847e-14, 
    2.409888e-14, 2.386532e-14, 2.447677e-14, 2.432971e-14, 2.451207e-14, 
    2.441893e-14, 2.457863e-14, 2.443487e-14, 2.468419e-14, 2.473866e-14, 
    2.470142e-14, 2.48446e-14, 2.44269e-14, 2.458686e-14, 2.339727e-14, 
    2.340417e-14, 2.343636e-14, 2.329502e-14, 2.328638e-14, 2.315728e-14, 
    2.327214e-14, 2.332113e-14, 2.344577e-14, 2.351965e-14, 2.358999e-14, 
    2.374506e-14, 2.391886e-14, 2.416301e-14, 2.433922e-14, 2.445771e-14, 
    2.438502e-14, 2.444919e-14, 2.437745e-14, 2.434387e-14, 2.471824e-14, 
    2.450765e-14, 2.482397e-14, 2.480641e-14, 2.466303e-14, 2.480838e-14, 
    2.340902e-14, 2.336928e-14, 2.323159e-14, 2.33393e-14, 2.314324e-14, 
    2.325287e-14, 2.331603e-14, 2.356059e-14, 2.36145e-14, 2.366455e-14, 
    2.376356e-14, 2.389093e-14, 2.411524e-14, 2.431131e-14, 2.449103e-14, 
    2.447784e-14, 2.448248e-14, 2.452271e-14, 2.442311e-14, 2.453907e-14, 
    2.455856e-14, 2.450762e-14, 2.480405e-14, 2.471918e-14, 2.480603e-14, 
    2.475074e-14, 2.338219e-14, 2.344909e-14, 2.341292e-14, 2.348094e-14, 
    2.3433e-14, 2.364654e-14, 2.371076e-14, 2.401248e-14, 2.388842e-14, 
    2.408604e-14, 2.390845e-14, 2.393986e-14, 2.409247e-14, 2.391802e-14, 
    2.430046e-14, 2.404082e-14, 2.452427e-14, 2.426372e-14, 2.454064e-14, 
    2.449023e-14, 2.457371e-14, 2.46486e-14, 2.474301e-14, 2.491766e-14, 
    2.487716e-14, 2.502359e-14, 2.354901e-14, 2.363611e-14, 2.362844e-14, 
    2.371977e-14, 2.378743e-14, 2.393444e-14, 2.417121e-14, 2.408203e-14, 
    2.424588e-14, 2.427884e-14, 2.402996e-14, 2.41826e-14, 2.369448e-14, 
    2.377298e-14, 2.372623e-14, 2.355582e-14, 2.410253e-14, 2.382113e-14, 
    2.434211e-14, 2.418865e-14, 2.463791e-14, 2.441394e-14, 2.485487e-14, 
    2.504461e-14, 2.52239e-14, 2.543423e-14, 2.368373e-14, 2.362445e-14, 
    2.373064e-14, 2.387796e-14, 2.401509e-14, 2.419803e-14, 2.421679e-14, 
    2.425115e-14, 2.434029e-14, 2.441537e-14, 2.426201e-14, 2.44342e-14, 
    2.379119e-14, 2.412704e-14, 2.360202e-14, 2.375947e-14, 2.386923e-14, 
    2.382105e-14, 2.407181e-14, 2.413111e-14, 2.437286e-14, 2.424773e-14, 
    2.49977e-14, 2.466441e-14, 2.559502e-14, 2.533313e-14, 2.360376e-14, 
    2.368352e-14, 2.396221e-14, 2.382939e-14, 2.421026e-14, 2.43045e-14, 
    2.438125e-14, 2.447953e-14, 2.449016e-14, 2.45485e-14, 2.445292e-14, 
    2.454472e-14, 2.419839e-14, 2.435284e-14, 2.393024e-14, 2.403273e-14, 
    2.398555e-14, 2.393385e-14, 2.409359e-14, 2.426438e-14, 2.426805e-14, 
    2.432294e-14, 2.447798e-14, 2.421176e-14, 2.504085e-14, 2.452707e-14, 
    2.377065e-14, 2.392496e-14, 2.394706e-14, 2.388719e-14, 2.429503e-14, 
    2.414684e-14, 2.454708e-14, 2.443857e-14, 2.461649e-14, 2.452799e-14, 
    2.451497e-14, 2.440159e-14, 2.433112e-14, 2.41536e-14, 2.400965e-14, 
    2.389583e-14, 2.392227e-14, 2.404738e-14, 2.427485e-14, 2.449108e-14, 
    2.444362e-14, 2.460291e-14, 2.418248e-14, 2.435831e-14, 2.429026e-14, 
    2.446788e-14, 2.407965e-14, 2.441006e-14, 2.399556e-14, 2.403175e-14, 
    2.414389e-14, 2.437029e-14, 2.442054e-14, 2.447424e-14, 2.444109e-14, 
    2.428066e-14, 2.425443e-14, 2.414115e-14, 2.410991e-14, 2.402384e-14, 
    2.39527e-14, 2.401769e-14, 2.408603e-14, 2.428071e-14, 2.445684e-14, 
    2.464963e-14, 2.469694e-14, 2.492342e-14, 2.473897e-14, 2.504371e-14, 
    2.478447e-14, 2.523413e-14, 2.442929e-14, 2.477695e-14, 2.4149e-14, 
    2.421624e-14, 2.433811e-14, 2.461884e-14, 2.446708e-14, 2.464462e-14, 
    2.42534e-14, 2.40517e-14, 2.399967e-14, 2.390274e-14, 2.400188e-14, 
    2.399381e-14, 2.408887e-14, 2.40583e-14, 2.428718e-14, 2.416409e-14, 
    2.451461e-14, 2.464318e-14, 2.500819e-14, 2.523332e-14, 2.54636e-14, 
    2.556561e-14, 2.55967e-14, 2.56097e-14 ;

 F_NIT =
  3.862229e-11, 3.895483e-11, 3.889006e-11, 3.915913e-11, 3.900975e-11, 
    3.91861e-11, 3.868957e-11, 3.896803e-11, 3.879014e-11, 3.865213e-11, 
    3.9684e-11, 3.917112e-11, 4.022054e-11, 3.989069e-11, 4.072198e-11, 
    4.016909e-11, 4.083394e-11, 4.070598e-11, 4.109177e-11, 4.098104e-11, 
    4.147654e-11, 4.114291e-11, 4.173464e-11, 4.139675e-11, 4.14495e-11, 
    4.11319e-11, 3.92741e-11, 3.961999e-11, 3.925365e-11, 3.930286e-11, 
    3.928077e-11, 3.901281e-11, 3.887813e-11, 3.85969e-11, 3.864787e-11, 
    3.885446e-11, 3.932497e-11, 3.916492e-11, 3.956894e-11, 3.95598e-11, 
    4.001207e-11, 3.980781e-11, 4.057205e-11, 4.035406e-11, 4.098566e-11, 
    4.082632e-11, 4.097815e-11, 4.093208e-11, 4.097874e-11, 4.07452e-11, 
    4.084516e-11, 4.063998e-11, 3.984608e-11, 4.007857e-11, 3.938724e-11, 
    3.897455e-11, 3.870174e-11, 3.850875e-11, 3.853599e-11, 3.858797e-11, 
    3.885567e-11, 3.910825e-11, 3.930132e-11, 3.943073e-11, 3.955847e-11, 
    3.99464e-11, 4.015257e-11, 4.061618e-11, 4.053232e-11, 4.067444e-11, 
    4.081048e-11, 4.10394e-11, 4.100168e-11, 4.110269e-11, 4.067068e-11, 
    4.095752e-11, 4.048455e-11, 4.061362e-11, 3.959322e-11, 3.920809e-11, 
    3.904494e-11, 3.890246e-11, 3.855695e-11, 3.879537e-11, 3.870129e-11, 
    3.892531e-11, 3.906801e-11, 3.89974e-11, 3.943427e-11, 3.926411e-11, 
    4.01648e-11, 3.977553e-11, 4.079461e-11, 4.054952e-11, 4.085346e-11, 
    4.069822e-11, 4.096439e-11, 4.072479e-11, 4.114031e-11, 4.123111e-11, 
    4.116903e-11, 4.140766e-11, 4.071149e-11, 4.09781e-11, 3.899545e-11, 
    3.900696e-11, 3.906061e-11, 3.882503e-11, 3.881064e-11, 3.859547e-11, 
    3.878689e-11, 3.886856e-11, 3.907629e-11, 3.919942e-11, 3.931666e-11, 
    3.95751e-11, 3.986476e-11, 4.027168e-11, 4.056537e-11, 4.076285e-11, 
    4.06417e-11, 4.074864e-11, 4.062909e-11, 4.057311e-11, 4.119707e-11, 
    4.084608e-11, 4.137328e-11, 4.134403e-11, 4.110505e-11, 4.13473e-11, 
    3.901503e-11, 3.89488e-11, 3.871931e-11, 3.889884e-11, 3.857207e-11, 
    3.875479e-11, 3.886005e-11, 3.926764e-11, 3.93575e-11, 3.944091e-11, 
    3.960593e-11, 3.981822e-11, 4.019208e-11, 4.051885e-11, 4.081839e-11, 
    4.07964e-11, 4.080413e-11, 4.087118e-11, 4.070518e-11, 4.089846e-11, 
    4.093093e-11, 4.084603e-11, 4.134009e-11, 4.119863e-11, 4.134338e-11, 
    4.125124e-11, 3.897032e-11, 3.908181e-11, 3.902153e-11, 3.913491e-11, 
    3.9055e-11, 3.94109e-11, 3.951793e-11, 4.002081e-11, 3.981403e-11, 
    4.014339e-11, 3.984742e-11, 3.989977e-11, 4.015412e-11, 3.986337e-11, 
    4.050077e-11, 4.006803e-11, 4.087378e-11, 4.043953e-11, 4.090106e-11, 
    4.081705e-11, 4.095619e-11, 4.108101e-11, 4.123835e-11, 4.152944e-11, 
    4.146193e-11, 4.170599e-11, 3.924834e-11, 3.939352e-11, 3.938073e-11, 
    3.953295e-11, 3.964572e-11, 3.989074e-11, 4.028535e-11, 4.013671e-11, 
    4.04098e-11, 4.046474e-11, 4.004993e-11, 4.030433e-11, 3.949081e-11, 
    3.962163e-11, 3.954371e-11, 3.925971e-11, 4.017088e-11, 3.970188e-11, 
    4.057018e-11, 4.031442e-11, 4.106318e-11, 4.06899e-11, 4.142479e-11, 
    4.174102e-11, 4.203983e-11, 4.239039e-11, 3.947288e-11, 3.937409e-11, 
    3.955107e-11, 3.97966e-11, 4.002515e-11, 4.033005e-11, 4.036131e-11, 
    4.041858e-11, 4.056714e-11, 4.069228e-11, 4.043668e-11, 4.072366e-11, 
    3.965198e-11, 4.021173e-11, 3.93367e-11, 3.959912e-11, 3.978204e-11, 
    3.970175e-11, 4.011969e-11, 4.021851e-11, 4.062144e-11, 4.041289e-11, 
    4.166283e-11, 4.110735e-11, 4.265837e-11, 4.222189e-11, 3.93396e-11, 
    3.947253e-11, 3.993702e-11, 3.971566e-11, 4.035044e-11, 4.05075e-11, 
    4.063541e-11, 4.079922e-11, 4.081693e-11, 4.091417e-11, 4.075487e-11, 
    4.090787e-11, 4.033065e-11, 4.058806e-11, 3.988374e-11, 4.005456e-11, 
    3.997593e-11, 3.988975e-11, 4.015599e-11, 4.044064e-11, 4.044674e-11, 
    4.053824e-11, 4.079663e-11, 4.035294e-11, 4.173475e-11, 4.087846e-11, 
    3.961775e-11, 3.987494e-11, 3.991176e-11, 3.981198e-11, 4.049172e-11, 
    4.024472e-11, 4.09118e-11, 4.073094e-11, 4.102748e-11, 4.087998e-11, 
    4.085829e-11, 4.066932e-11, 4.055187e-11, 4.025599e-11, 4.001608e-11, 
    3.982639e-11, 3.987045e-11, 4.007897e-11, 4.045808e-11, 4.081846e-11, 
    4.073937e-11, 4.100485e-11, 4.030414e-11, 4.059717e-11, 4.048377e-11, 
    4.07798e-11, 4.013274e-11, 4.068344e-11, 3.99926e-11, 4.005292e-11, 
    4.023982e-11, 4.061715e-11, 4.07009e-11, 4.07904e-11, 4.073515e-11, 
    4.046776e-11, 4.042404e-11, 4.023524e-11, 4.018318e-11, 4.003974e-11, 
    3.992117e-11, 4.002948e-11, 4.014339e-11, 4.046784e-11, 4.07614e-11, 
    4.108272e-11, 4.116157e-11, 4.153903e-11, 4.123162e-11, 4.173952e-11, 
    4.130746e-11, 4.205689e-11, 4.071549e-11, 4.129491e-11, 4.024834e-11, 
    4.036041e-11, 4.056351e-11, 4.10314e-11, 4.077846e-11, 4.107436e-11, 
    4.042233e-11, 4.008617e-11, 3.999945e-11, 3.98379e-11, 4.000314e-11, 
    3.998969e-11, 4.014812e-11, 4.009716e-11, 4.047863e-11, 4.027349e-11, 
    4.085768e-11, 4.107197e-11, 4.168032e-11, 4.205554e-11, 4.243934e-11, 
    4.260935e-11, 4.266116e-11, 4.268283e-11 ;

 F_NIT_vr =
  2.478151e-10, 2.489173e-10, 2.487025e-10, 2.49592e-10, 2.490983e-10, 
    2.496803e-10, 2.480373e-10, 2.489591e-10, 2.483703e-10, 2.479122e-10, 
    2.513175e-10, 2.496296e-10, 2.530751e-10, 2.519958e-10, 2.547082e-10, 
    2.529062e-10, 2.550716e-10, 2.546558e-10, 2.559074e-10, 2.555482e-10, 
    2.571496e-10, 2.560722e-10, 2.579806e-10, 2.56892e-10, 2.570617e-10, 
    2.560353e-10, 2.499713e-10, 2.511091e-10, 2.499034e-10, 2.500656e-10, 
    2.499926e-10, 2.491072e-10, 2.486612e-10, 2.477287e-10, 2.478976e-10, 
    2.485824e-10, 2.501366e-10, 2.496085e-10, 2.509393e-10, 2.509093e-10, 
    2.523924e-10, 2.517233e-10, 2.542199e-10, 2.535093e-10, 2.555629e-10, 
    2.550456e-10, 2.55538e-10, 2.553883e-10, 2.555392e-10, 2.547813e-10, 
    2.551054e-10, 2.544388e-10, 2.518517e-10, 2.526126e-10, 2.503432e-10, 
    2.4898e-10, 2.480765e-10, 2.474358e-10, 2.475258e-10, 2.476984e-10, 
    2.485858e-10, 2.494211e-10, 2.500582e-10, 2.504842e-10, 2.509042e-10, 
    2.521766e-10, 2.528512e-10, 2.543627e-10, 2.540899e-10, 2.545517e-10, 
    2.549939e-10, 2.557359e-10, 2.556136e-10, 2.559403e-10, 2.545384e-10, 
    2.554696e-10, 2.539322e-10, 2.543523e-10, 2.510198e-10, 2.497521e-10, 
    2.492126e-10, 2.487413e-10, 2.475952e-10, 2.483863e-10, 2.48074e-10, 
    2.488161e-10, 2.492879e-10, 2.490541e-10, 2.504956e-10, 2.499344e-10, 
    2.528907e-10, 2.516163e-10, 2.549427e-10, 2.541453e-10, 2.55133e-10, 
    2.546288e-10, 2.554922e-10, 2.547147e-10, 2.560616e-10, 2.563553e-10, 
    2.56154e-10, 2.569253e-10, 2.546699e-10, 2.555352e-10, 2.490491e-10, 
    2.490872e-10, 2.492643e-10, 2.484841e-10, 2.484364e-10, 2.477223e-10, 
    2.483571e-10, 2.486276e-10, 2.493146e-10, 2.497208e-10, 2.501071e-10, 
    2.50958e-10, 2.519084e-10, 2.532392e-10, 2.541966e-10, 2.548385e-10, 
    2.544446e-10, 2.547918e-10, 2.54403e-10, 2.542205e-10, 2.562445e-10, 
    2.551072e-10, 2.568136e-10, 2.567192e-10, 2.559459e-10, 2.567291e-10, 
    2.491134e-10, 2.48894e-10, 2.481335e-10, 2.487281e-10, 2.476442e-10, 
    2.482504e-10, 2.485987e-10, 2.499455e-10, 2.502416e-10, 2.505163e-10, 
    2.510589e-10, 2.517554e-10, 2.529789e-10, 2.540445e-10, 2.550186e-10, 
    2.549468e-10, 2.549718e-10, 2.55189e-10, 2.546497e-10, 2.552769e-10, 
    2.553818e-10, 2.551065e-10, 2.567058e-10, 2.562486e-10, 2.567161e-10, 
    2.56418e-10, 2.489649e-10, 2.493331e-10, 2.491335e-10, 2.495081e-10, 
    2.492435e-10, 2.504176e-10, 2.507694e-10, 2.524191e-10, 2.517416e-10, 
    2.5282e-10, 2.518507e-10, 2.520222e-10, 2.528537e-10, 2.519024e-10, 
    2.539846e-10, 2.525714e-10, 2.551971e-10, 2.537839e-10, 2.552851e-10, 
    2.550122e-10, 2.554632e-10, 2.558676e-10, 2.563763e-10, 2.573158e-10, 
    2.570977e-10, 2.57884e-10, 2.498826e-10, 2.503606e-10, 2.503186e-10, 
    2.508192e-10, 2.511895e-10, 2.519936e-10, 2.532838e-10, 2.52798e-10, 
    2.536892e-10, 2.538682e-10, 2.525133e-10, 2.533445e-10, 2.506783e-10, 
    2.511078e-10, 2.508519e-10, 2.49916e-10, 2.529072e-10, 2.513704e-10, 
    2.542092e-10, 2.533753e-10, 2.558091e-10, 2.545977e-10, 2.569777e-10, 
    2.57996e-10, 2.589561e-10, 2.600774e-10, 2.506217e-10, 2.502961e-10, 
    2.508783e-10, 2.516844e-10, 2.524329e-10, 2.534293e-10, 2.535311e-10, 
    2.537174e-10, 2.54201e-10, 2.546081e-10, 2.537755e-10, 2.547094e-10, 
    2.512067e-10, 2.530407e-10, 2.501694e-10, 2.510328e-10, 2.516332e-10, 
    2.513698e-10, 2.527391e-10, 2.530616e-10, 2.543744e-10, 2.536956e-10, 
    2.577436e-10, 2.559506e-10, 2.609326e-10, 2.595381e-10, 2.501822e-10, 
    2.506196e-10, 2.521441e-10, 2.514184e-10, 2.534952e-10, 2.540071e-10, 
    2.54423e-10, 2.549553e-10, 2.550123e-10, 2.553279e-10, 2.548103e-10, 
    2.55307e-10, 2.534285e-10, 2.542674e-10, 2.51967e-10, 2.525258e-10, 
    2.522685e-10, 2.519858e-10, 2.528568e-10, 2.537855e-10, 2.538054e-10, 
    2.541028e-10, 2.549417e-10, 2.534986e-10, 2.579733e-10, 2.552066e-10, 
    2.510969e-10, 2.519401e-10, 2.520608e-10, 2.517339e-10, 2.53955e-10, 
    2.531495e-10, 2.553202e-10, 2.547327e-10, 2.556946e-10, 2.552163e-10, 
    2.551454e-10, 2.545316e-10, 2.541489e-10, 2.531842e-10, 2.523994e-10, 
    2.517781e-10, 2.51922e-10, 2.526046e-10, 2.538416e-10, 2.55014e-10, 
    2.547567e-10, 2.55618e-10, 2.533389e-10, 2.542937e-10, 2.539239e-10, 
    2.548871e-10, 2.527838e-10, 2.545782e-10, 2.523252e-10, 2.525222e-10, 
    2.531327e-10, 2.543623e-10, 2.546346e-10, 2.549252e-10, 2.547454e-10, 
    2.538751e-10, 2.537325e-10, 2.531162e-10, 2.529456e-10, 2.524768e-10, 
    2.52088e-10, 2.524427e-10, 2.528145e-10, 2.538735e-10, 2.548282e-10, 
    2.558699e-10, 2.561251e-10, 2.573429e-10, 2.563506e-10, 2.579873e-10, 
    2.565943e-10, 2.590065e-10, 2.546821e-10, 2.565598e-10, 2.531607e-10, 
    2.53526e-10, 2.541873e-10, 2.557062e-10, 2.548859e-10, 2.558452e-10, 
    2.537267e-10, 2.526284e-10, 2.523447e-10, 2.518154e-10, 2.523563e-10, 
    2.523123e-10, 2.528303e-10, 2.526633e-10, 2.539079e-10, 2.532391e-10, 
    2.551399e-10, 2.558345e-10, 2.577983e-10, 2.590032e-10, 2.602318e-10, 
    2.60774e-10, 2.609391e-10, 2.610078e-10,
  1.2614e-10, 1.27101e-10, 1.26914e-10, 1.276906e-10, 1.272597e-10, 
    1.277685e-10, 1.263347e-10, 1.271392e-10, 1.266254e-10, 1.262265e-10, 
    1.292027e-10, 1.277254e-10, 1.30745e-10, 1.297976e-10, 1.321827e-10, 
    1.305973e-10, 1.325032e-10, 1.32137e-10, 1.332409e-10, 1.329243e-10, 
    1.343395e-10, 1.333871e-10, 1.350756e-10, 1.34112e-10, 1.342625e-10, 
    1.333557e-10, 1.280223e-10, 1.290184e-10, 1.279634e-10, 1.281052e-10, 
    1.280416e-10, 1.272685e-10, 1.268795e-10, 1.260668e-10, 1.262142e-10, 
    1.268113e-10, 1.28169e-10, 1.277076e-10, 1.288721e-10, 1.288457e-10, 
    1.301466e-10, 1.295594e-10, 1.317534e-10, 1.311285e-10, 1.329375e-10, 
    1.324817e-10, 1.329161e-10, 1.327843e-10, 1.329178e-10, 1.322494e-10, 
    1.325356e-10, 1.319482e-10, 1.296693e-10, 1.303374e-10, 1.283485e-10, 
    1.271579e-10, 1.263699e-10, 1.258118e-10, 1.258906e-10, 1.260409e-10, 
    1.268148e-10, 1.275441e-10, 1.28101e-10, 1.28474e-10, 1.288419e-10, 
    1.299576e-10, 1.3055e-10, 1.318798e-10, 1.316396e-10, 1.320467e-10, 
    1.324364e-10, 1.330912e-10, 1.329834e-10, 1.332721e-10, 1.320361e-10, 
    1.32857e-10, 1.315028e-10, 1.318727e-10, 1.289413e-10, 1.278321e-10, 
    1.273611e-10, 1.269499e-10, 1.259512e-10, 1.266406e-10, 1.263686e-10, 
    1.270161e-10, 1.27428e-10, 1.272242e-10, 1.284842e-10, 1.279938e-10, 
    1.305851e-10, 1.294665e-10, 1.323909e-10, 1.316889e-10, 1.325594e-10, 
    1.321149e-10, 1.328767e-10, 1.321911e-10, 1.333797e-10, 1.336391e-10, 
    1.334618e-10, 1.341434e-10, 1.321531e-10, 1.32916e-10, 1.272185e-10, 
    1.272517e-10, 1.274066e-10, 1.267263e-10, 1.266847e-10, 1.260627e-10, 
    1.266162e-10, 1.268521e-10, 1.27452e-10, 1.278072e-10, 1.281453e-10, 
    1.288898e-10, 1.297231e-10, 1.30892e-10, 1.317343e-10, 1.323001e-10, 
    1.319531e-10, 1.322594e-10, 1.31917e-10, 1.317567e-10, 1.335419e-10, 
    1.325383e-10, 1.340453e-10, 1.339618e-10, 1.33279e-10, 1.339712e-10, 
    1.272751e-10, 1.270839e-10, 1.264208e-10, 1.269396e-10, 1.259951e-10, 
    1.265234e-10, 1.268275e-10, 1.280039e-10, 1.282631e-10, 1.285033e-10, 
    1.289786e-10, 1.295895e-10, 1.306636e-10, 1.31601e-10, 1.324591e-10, 
    1.323961e-10, 1.324183e-10, 1.326101e-10, 1.32135e-10, 1.326882e-10, 
    1.327811e-10, 1.325382e-10, 1.339506e-10, 1.335466e-10, 1.3396e-10, 
    1.336969e-10, 1.27146e-10, 1.274679e-10, 1.272939e-10, 1.276211e-10, 
    1.273905e-10, 1.284168e-10, 1.287251e-10, 1.301716e-10, 1.295774e-10, 
    1.305238e-10, 1.296735e-10, 1.298239e-10, 1.305544e-10, 1.297194e-10, 
    1.315491e-10, 1.303073e-10, 1.326176e-10, 1.313735e-10, 1.326957e-10, 
    1.324553e-10, 1.328535e-10, 1.332103e-10, 1.3366e-10, 1.344908e-10, 
    1.342983e-10, 1.349943e-10, 1.279483e-10, 1.283667e-10, 1.2833e-10, 
    1.287685e-10, 1.290931e-10, 1.29798e-10, 1.309313e-10, 1.305047e-10, 
    1.312884e-10, 1.314459e-10, 1.302555e-10, 1.309858e-10, 1.286472e-10, 
    1.290238e-10, 1.287996e-10, 1.279812e-10, 1.306028e-10, 1.292548e-10, 
    1.317483e-10, 1.310149e-10, 1.331594e-10, 1.320912e-10, 1.341923e-10, 
    1.350939e-10, 1.35945e-10, 1.369414e-10, 1.285955e-10, 1.283109e-10, 
    1.288207e-10, 1.295271e-10, 1.301843e-10, 1.310596e-10, 1.311494e-10, 
    1.313136e-10, 1.317395e-10, 1.32098e-10, 1.313654e-10, 1.32188e-10, 
    1.291109e-10, 1.307201e-10, 1.282032e-10, 1.28959e-10, 1.294855e-10, 
    1.292546e-10, 1.30456e-10, 1.307398e-10, 1.318951e-10, 1.312975e-10, 
    1.34871e-10, 1.332855e-10, 1.377022e-10, 1.364626e-10, 1.282115e-10, 
    1.285945e-10, 1.299309e-10, 1.292945e-10, 1.311182e-10, 1.315685e-10, 
    1.319351e-10, 1.324042e-10, 1.324549e-10, 1.327332e-10, 1.322773e-10, 
    1.327152e-10, 1.310615e-10, 1.317995e-10, 1.297781e-10, 1.302689e-10, 
    1.300431e-10, 1.297954e-10, 1.305603e-10, 1.313769e-10, 1.313946e-10, 
    1.316568e-10, 1.323964e-10, 1.311256e-10, 1.350757e-10, 1.326307e-10, 
    1.290127e-10, 1.297524e-10, 1.298585e-10, 1.295716e-10, 1.315233e-10, 
    1.308149e-10, 1.327264e-10, 1.322088e-10, 1.330573e-10, 1.326354e-10, 
    1.325734e-10, 1.320323e-10, 1.316959e-10, 1.308473e-10, 1.301584e-10, 
    1.296132e-10, 1.297399e-10, 1.303391e-10, 1.31427e-10, 1.324594e-10, 
    1.32233e-10, 1.329928e-10, 1.309856e-10, 1.318258e-10, 1.315007e-10, 
    1.323489e-10, 1.304934e-10, 1.320722e-10, 1.300909e-10, 1.302642e-10, 
    1.308008e-10, 1.318827e-10, 1.321228e-10, 1.32379e-10, 1.322209e-10, 
    1.314547e-10, 1.313294e-10, 1.307878e-10, 1.306383e-10, 1.302265e-10, 
    1.298858e-10, 1.30197e-10, 1.305241e-10, 1.314551e-10, 1.322961e-10, 
    1.332154e-10, 1.334408e-10, 1.345181e-10, 1.336407e-10, 1.350894e-10, 
    1.338569e-10, 1.359932e-10, 1.321642e-10, 1.338212e-10, 1.308253e-10, 
    1.311469e-10, 1.31729e-10, 1.330683e-10, 1.323449e-10, 1.331912e-10, 
    1.313245e-10, 1.303597e-10, 1.301107e-10, 1.296463e-10, 1.301213e-10, 
    1.300827e-10, 1.305378e-10, 1.303915e-10, 1.31486e-10, 1.308977e-10, 
    1.325717e-10, 1.331846e-10, 1.349212e-10, 1.359897e-10, 1.370808e-10, 
    1.375634e-10, 1.377104e-10, 1.377718e-10,
  1.185433e-10, 1.195951e-10, 1.193904e-10, 1.20241e-10, 1.197688e-10, 
    1.203263e-10, 1.187562e-10, 1.196369e-10, 1.190744e-10, 1.186379e-10, 
    1.21899e-10, 1.20279e-10, 1.235922e-10, 1.225517e-10, 1.251728e-10, 
    1.2343e-10, 1.255255e-10, 1.251225e-10, 1.263374e-10, 1.259889e-10, 
    1.27548e-10, 1.264984e-10, 1.283596e-10, 1.272971e-10, 1.27463e-10, 
    1.264638e-10, 1.206044e-10, 1.216968e-10, 1.205398e-10, 1.206953e-10, 
    1.206255e-10, 1.197785e-10, 1.193526e-10, 1.184631e-10, 1.186244e-10, 
    1.192779e-10, 1.207652e-10, 1.202595e-10, 1.21536e-10, 1.215071e-10, 
    1.229348e-10, 1.222902e-10, 1.247005e-10, 1.240134e-10, 1.260034e-10, 
    1.255017e-10, 1.259798e-10, 1.258347e-10, 1.259817e-10, 1.252462e-10, 
    1.255611e-10, 1.249147e-10, 1.224108e-10, 1.231444e-10, 1.209619e-10, 
    1.196575e-10, 1.187948e-10, 1.181841e-10, 1.182704e-10, 1.184348e-10, 
    1.192817e-10, 1.200804e-10, 1.206906e-10, 1.210995e-10, 1.215029e-10, 
    1.227274e-10, 1.233779e-10, 1.248396e-10, 1.245754e-10, 1.250232e-10, 
    1.254518e-10, 1.261726e-10, 1.260539e-10, 1.263719e-10, 1.250114e-10, 
    1.259149e-10, 1.244249e-10, 1.248317e-10, 1.216123e-10, 1.203959e-10, 
    1.198801e-10, 1.194297e-10, 1.183367e-10, 1.19091e-10, 1.187934e-10, 
    1.19502e-10, 1.199532e-10, 1.1973e-10, 1.211107e-10, 1.205731e-10, 
    1.234165e-10, 1.221883e-10, 1.254018e-10, 1.246296e-10, 1.255872e-10, 
    1.250982e-10, 1.259365e-10, 1.251819e-10, 1.264903e-10, 1.267761e-10, 
    1.265807e-10, 1.273316e-10, 1.251401e-10, 1.259797e-10, 1.197237e-10, 
    1.197601e-10, 1.199298e-10, 1.191848e-10, 1.191393e-10, 1.184587e-10, 
    1.190643e-10, 1.193226e-10, 1.199794e-10, 1.203686e-10, 1.207391e-10, 
    1.215555e-10, 1.2247e-10, 1.237537e-10, 1.246796e-10, 1.253018e-10, 
    1.249201e-10, 1.252571e-10, 1.248804e-10, 1.247041e-10, 1.26669e-10, 
    1.25564e-10, 1.272235e-10, 1.271315e-10, 1.263794e-10, 1.271418e-10, 
    1.197857e-10, 1.195763e-10, 1.188505e-10, 1.194183e-10, 1.183846e-10, 
    1.189627e-10, 1.192956e-10, 1.205842e-10, 1.208682e-10, 1.211317e-10, 
    1.216529e-10, 1.223231e-10, 1.235027e-10, 1.24533e-10, 1.254768e-10, 
    1.254075e-10, 1.254319e-10, 1.256431e-10, 1.251202e-10, 1.25729e-10, 
    1.258313e-10, 1.255639e-10, 1.271191e-10, 1.26674e-10, 1.271295e-10, 
    1.268396e-10, 1.196444e-10, 1.199969e-10, 1.198063e-10, 1.201647e-10, 
    1.199121e-10, 1.210368e-10, 1.213749e-10, 1.229624e-10, 1.223099e-10, 
    1.233491e-10, 1.224153e-10, 1.225805e-10, 1.233829e-10, 1.224657e-10, 
    1.24476e-10, 1.231114e-10, 1.256513e-10, 1.242829e-10, 1.257372e-10, 
    1.254727e-10, 1.259109e-10, 1.263038e-10, 1.267991e-10, 1.277147e-10, 
    1.275024e-10, 1.282698e-10, 1.205232e-10, 1.209819e-10, 1.209416e-10, 
    1.214224e-10, 1.217785e-10, 1.22552e-10, 1.237968e-10, 1.233281e-10, 
    1.241893e-10, 1.243624e-10, 1.230544e-10, 1.238567e-10, 1.212894e-10, 
    1.217026e-10, 1.214565e-10, 1.205594e-10, 1.23436e-10, 1.21956e-10, 
    1.246949e-10, 1.238887e-10, 1.262477e-10, 1.250721e-10, 1.273856e-10, 
    1.283798e-10, 1.293189e-10, 1.304194e-10, 1.212327e-10, 1.209206e-10, 
    1.214797e-10, 1.222548e-10, 1.229762e-10, 1.239378e-10, 1.240364e-10, 
    1.24217e-10, 1.246853e-10, 1.250795e-10, 1.24274e-10, 1.251785e-10, 
    1.217983e-10, 1.235648e-10, 1.208027e-10, 1.216315e-10, 1.222091e-10, 
    1.219557e-10, 1.232746e-10, 1.235863e-10, 1.248565e-10, 1.241992e-10, 
    1.281341e-10, 1.263867e-10, 1.312603e-10, 1.298906e-10, 1.208117e-10, 
    1.212316e-10, 1.22698e-10, 1.219994e-10, 1.240022e-10, 1.244972e-10, 
    1.249004e-10, 1.254164e-10, 1.254722e-10, 1.257785e-10, 1.252768e-10, 
    1.257587e-10, 1.239399e-10, 1.247513e-10, 1.225302e-10, 1.230691e-10, 
    1.228211e-10, 1.225492e-10, 1.233892e-10, 1.242867e-10, 1.24306e-10, 
    1.245943e-10, 1.254082e-10, 1.240103e-10, 1.283601e-10, 1.25666e-10, 
    1.216903e-10, 1.225021e-10, 1.226184e-10, 1.223035e-10, 1.244476e-10, 
    1.236689e-10, 1.25771e-10, 1.252014e-10, 1.261353e-10, 1.256709e-10, 
    1.256026e-10, 1.250073e-10, 1.246373e-10, 1.237045e-10, 1.229478e-10, 
    1.223492e-10, 1.224883e-10, 1.231462e-10, 1.243417e-10, 1.254772e-10, 
    1.252281e-10, 1.260642e-10, 1.238565e-10, 1.247801e-10, 1.244227e-10, 
    1.253556e-10, 1.233156e-10, 1.250515e-10, 1.228736e-10, 1.230639e-10, 
    1.236534e-10, 1.248428e-10, 1.251068e-10, 1.253887e-10, 1.252147e-10, 
    1.243721e-10, 1.242343e-10, 1.236391e-10, 1.234749e-10, 1.230225e-10, 
    1.226484e-10, 1.229901e-10, 1.233494e-10, 1.243725e-10, 1.252975e-10, 
    1.263094e-10, 1.265576e-10, 1.277449e-10, 1.267779e-10, 1.283751e-10, 
    1.270164e-10, 1.293724e-10, 1.251526e-10, 1.269768e-10, 1.236803e-10, 
    1.240337e-10, 1.246738e-10, 1.261476e-10, 1.253512e-10, 1.262828e-10, 
    1.24229e-10, 1.231689e-10, 1.228954e-10, 1.223855e-10, 1.22907e-10, 
    1.228646e-10, 1.233644e-10, 1.232037e-10, 1.244065e-10, 1.237598e-10, 
    1.256008e-10, 1.262755e-10, 1.281893e-10, 1.293683e-10, 1.305733e-10, 
    1.311067e-10, 1.312692e-10, 1.313372e-10,
  1.213295e-10, 1.224836e-10, 1.222589e-10, 1.231927e-10, 1.226743e-10, 
    1.232864e-10, 1.215631e-10, 1.225295e-10, 1.219121e-10, 1.214332e-10, 
    1.250149e-10, 1.232345e-10, 1.268775e-10, 1.257324e-10, 1.286186e-10, 
    1.26699e-10, 1.290074e-10, 1.285631e-10, 1.299027e-10, 1.295182e-10, 
    1.312389e-10, 1.300803e-10, 1.321352e-10, 1.309618e-10, 1.31145e-10, 
    1.300422e-10, 1.235918e-10, 1.247925e-10, 1.235209e-10, 1.236917e-10, 
    1.23615e-10, 1.22685e-10, 1.222175e-10, 1.212415e-10, 1.214184e-10, 
    1.221355e-10, 1.237686e-10, 1.23213e-10, 1.246155e-10, 1.245837e-10, 
    1.261539e-10, 1.254448e-10, 1.280981e-10, 1.273412e-10, 1.295343e-10, 
    1.28981e-10, 1.295083e-10, 1.293483e-10, 1.295103e-10, 1.286994e-10, 
    1.290466e-10, 1.283341e-10, 1.255774e-10, 1.263845e-10, 1.239846e-10, 
    1.225522e-10, 1.216054e-10, 1.209356e-10, 1.210302e-10, 1.212106e-10, 
    1.221397e-10, 1.230163e-10, 1.236865e-10, 1.241357e-10, 1.245792e-10, 
    1.259259e-10, 1.266417e-10, 1.282514e-10, 1.279602e-10, 1.284537e-10, 
    1.289261e-10, 1.29721e-10, 1.2959e-10, 1.299408e-10, 1.284407e-10, 
    1.294367e-10, 1.277945e-10, 1.282426e-10, 1.246997e-10, 1.233628e-10, 
    1.227965e-10, 1.22302e-10, 1.211029e-10, 1.219304e-10, 1.216039e-10, 
    1.223814e-10, 1.228767e-10, 1.226316e-10, 1.24148e-10, 1.235574e-10, 
    1.266842e-10, 1.253327e-10, 1.288709e-10, 1.280199e-10, 1.290753e-10, 
    1.285363e-10, 1.294605e-10, 1.286286e-10, 1.300714e-10, 1.303867e-10, 
    1.301712e-10, 1.309998e-10, 1.285825e-10, 1.295082e-10, 1.226248e-10, 
    1.226647e-10, 1.228509e-10, 1.220333e-10, 1.219834e-10, 1.212367e-10, 
    1.21901e-10, 1.221845e-10, 1.229054e-10, 1.233329e-10, 1.237398e-10, 
    1.246369e-10, 1.256425e-10, 1.270553e-10, 1.28075e-10, 1.287607e-10, 
    1.283401e-10, 1.287114e-10, 1.282963e-10, 1.28102e-10, 1.302686e-10, 
    1.290498e-10, 1.308805e-10, 1.307789e-10, 1.299491e-10, 1.307904e-10, 
    1.226928e-10, 1.224629e-10, 1.216665e-10, 1.222895e-10, 1.211555e-10, 
    1.217896e-10, 1.22155e-10, 1.235697e-10, 1.238816e-10, 1.241712e-10, 
    1.24744e-10, 1.25481e-10, 1.267789e-10, 1.279135e-10, 1.289536e-10, 
    1.288772e-10, 1.289041e-10, 1.29137e-10, 1.285606e-10, 1.292317e-10, 
    1.293445e-10, 1.290497e-10, 1.307653e-10, 1.302741e-10, 1.307767e-10, 
    1.304568e-10, 1.225376e-10, 1.229246e-10, 1.227154e-10, 1.231089e-10, 
    1.228316e-10, 1.24067e-10, 1.244385e-10, 1.261843e-10, 1.254665e-10, 
    1.266099e-10, 1.255824e-10, 1.257641e-10, 1.266472e-10, 1.256378e-10, 
    1.278508e-10, 1.263484e-10, 1.29146e-10, 1.276382e-10, 1.292408e-10, 
    1.289491e-10, 1.294322e-10, 1.298656e-10, 1.30412e-10, 1.314229e-10, 
    1.311885e-10, 1.32036e-10, 1.235027e-10, 1.240066e-10, 1.239622e-10, 
    1.244907e-10, 1.248821e-10, 1.257327e-10, 1.271028e-10, 1.265867e-10, 
    1.275349e-10, 1.277256e-10, 1.262855e-10, 1.271687e-10, 1.243445e-10, 
    1.247987e-10, 1.245282e-10, 1.235424e-10, 1.267055e-10, 1.250773e-10, 
    1.280919e-10, 1.272039e-10, 1.298038e-10, 1.285076e-10, 1.310595e-10, 
    1.321577e-10, 1.331954e-10, 1.344129e-10, 1.242821e-10, 1.239392e-10, 
    1.245536e-10, 1.254059e-10, 1.261994e-10, 1.27258e-10, 1.273665e-10, 
    1.275654e-10, 1.280813e-10, 1.285157e-10, 1.276283e-10, 1.286248e-10, 
    1.249041e-10, 1.268473e-10, 1.238097e-10, 1.247206e-10, 1.253556e-10, 
    1.250769e-10, 1.265278e-10, 1.26871e-10, 1.2827e-10, 1.275459e-10, 
    1.318862e-10, 1.299573e-10, 1.353436e-10, 1.338277e-10, 1.238195e-10, 
    1.24281e-10, 1.258934e-10, 1.25125e-10, 1.273288e-10, 1.278741e-10, 
    1.283183e-10, 1.288871e-10, 1.289486e-10, 1.292863e-10, 1.287331e-10, 
    1.292644e-10, 1.272602e-10, 1.28154e-10, 1.257087e-10, 1.263017e-10, 
    1.260287e-10, 1.257296e-10, 1.266539e-10, 1.276422e-10, 1.276634e-10, 
    1.279811e-10, 1.288784e-10, 1.273378e-10, 1.321361e-10, 1.291626e-10, 
    1.247851e-10, 1.25678e-10, 1.258058e-10, 1.254594e-10, 1.278194e-10, 
    1.269618e-10, 1.29278e-10, 1.286501e-10, 1.296798e-10, 1.291676e-10, 
    1.290923e-10, 1.284361e-10, 1.280284e-10, 1.270011e-10, 1.261682e-10, 
    1.255096e-10, 1.256626e-10, 1.263865e-10, 1.277028e-10, 1.289541e-10, 
    1.286795e-10, 1.296014e-10, 1.271684e-10, 1.281859e-10, 1.277921e-10, 
    1.2882e-10, 1.26573e-10, 1.284851e-10, 1.260865e-10, 1.262959e-10, 
    1.269448e-10, 1.28255e-10, 1.285458e-10, 1.288565e-10, 1.286647e-10, 
    1.277363e-10, 1.275846e-10, 1.269291e-10, 1.267483e-10, 1.262503e-10, 
    1.258387e-10, 1.262147e-10, 1.266102e-10, 1.277367e-10, 1.28756e-10, 
    1.298718e-10, 1.301456e-10, 1.314564e-10, 1.303889e-10, 1.321527e-10, 
    1.306523e-10, 1.332549e-10, 1.285964e-10, 1.306084e-10, 1.269744e-10, 
    1.273635e-10, 1.280688e-10, 1.296934e-10, 1.288152e-10, 1.298426e-10, 
    1.275786e-10, 1.264115e-10, 1.261105e-10, 1.255496e-10, 1.261233e-10, 
    1.260766e-10, 1.266267e-10, 1.264498e-10, 1.277742e-10, 1.27062e-10, 
    1.290904e-10, 1.298345e-10, 1.319471e-10, 1.332501e-10, 1.34583e-10, 
    1.351735e-10, 1.353534e-10, 1.354287e-10,
  1.320191e-10, 1.33252e-10, 1.330118e-10, 1.3401e-10, 1.334558e-10, 
    1.341102e-10, 1.322685e-10, 1.333011e-10, 1.326414e-10, 1.321298e-10, 
    1.359596e-10, 1.340547e-10, 1.379546e-10, 1.367277e-10, 1.398219e-10, 
    1.377633e-10, 1.402392e-10, 1.397623e-10, 1.412004e-10, 1.407875e-10, 
    1.426366e-10, 1.413913e-10, 1.436005e-10, 1.423386e-10, 1.425356e-10, 
    1.413503e-10, 1.344368e-10, 1.357216e-10, 1.343608e-10, 1.345436e-10, 
    1.344616e-10, 1.334672e-10, 1.329677e-10, 1.319251e-10, 1.32114e-10, 
    1.3288e-10, 1.346258e-10, 1.340317e-10, 1.355318e-10, 1.354978e-10, 
    1.371791e-10, 1.364196e-10, 1.392633e-10, 1.384516e-10, 1.408048e-10, 
    1.402108e-10, 1.407768e-10, 1.406051e-10, 1.407791e-10, 1.399086e-10, 
    1.402812e-10, 1.395166e-10, 1.365616e-10, 1.374263e-10, 1.348569e-10, 
    1.333254e-10, 1.323137e-10, 1.315985e-10, 1.316995e-10, 1.318921e-10, 
    1.328845e-10, 1.338214e-10, 1.345379e-10, 1.350185e-10, 1.35493e-10, 
    1.369351e-10, 1.377019e-10, 1.394278e-10, 1.391154e-10, 1.396449e-10, 
    1.401518e-10, 1.410053e-10, 1.408646e-10, 1.412414e-10, 1.396309e-10, 
    1.407e-10, 1.389376e-10, 1.394184e-10, 1.356222e-10, 1.341918e-10, 
    1.335866e-10, 1.33058e-10, 1.317772e-10, 1.326609e-10, 1.323121e-10, 
    1.331427e-10, 1.336721e-10, 1.334101e-10, 1.350316e-10, 1.343999e-10, 
    1.377474e-10, 1.362997e-10, 1.400926e-10, 1.391795e-10, 1.40312e-10, 
    1.397334e-10, 1.407256e-10, 1.398325e-10, 1.413818e-10, 1.417205e-10, 
    1.414889e-10, 1.423794e-10, 1.397831e-10, 1.407769e-10, 1.334028e-10, 
    1.334455e-10, 1.336446e-10, 1.327709e-10, 1.327175e-10, 1.319199e-10, 
    1.326295e-10, 1.329323e-10, 1.337028e-10, 1.341598e-10, 1.34595e-10, 
    1.355548e-10, 1.366314e-10, 1.381451e-10, 1.392386e-10, 1.399743e-10, 
    1.395229e-10, 1.399214e-10, 1.39476e-10, 1.392675e-10, 1.415935e-10, 
    1.402846e-10, 1.422511e-10, 1.421419e-10, 1.412504e-10, 1.421542e-10, 
    1.334755e-10, 1.332298e-10, 1.323789e-10, 1.330446e-10, 1.318333e-10, 
    1.325105e-10, 1.329009e-10, 1.344131e-10, 1.347467e-10, 1.350564e-10, 
    1.356694e-10, 1.364584e-10, 1.378489e-10, 1.390654e-10, 1.401813e-10, 
    1.400994e-10, 1.401282e-10, 1.403782e-10, 1.397595e-10, 1.404799e-10, 
    1.40601e-10, 1.402845e-10, 1.421273e-10, 1.415994e-10, 1.421396e-10, 
    1.417957e-10, 1.333097e-10, 1.337233e-10, 1.334997e-10, 1.339204e-10, 
    1.336239e-10, 1.34945e-10, 1.353426e-10, 1.372118e-10, 1.364428e-10, 
    1.376678e-10, 1.36567e-10, 1.367616e-10, 1.377079e-10, 1.366263e-10, 
    1.389982e-10, 1.373876e-10, 1.403879e-10, 1.387703e-10, 1.404896e-10, 
    1.401765e-10, 1.406952e-10, 1.411607e-10, 1.417476e-10, 1.428343e-10, 
    1.425822e-10, 1.434938e-10, 1.343414e-10, 1.348804e-10, 1.348329e-10, 
    1.353982e-10, 1.358173e-10, 1.367279e-10, 1.38196e-10, 1.376429e-10, 
    1.386593e-10, 1.388638e-10, 1.3732e-10, 1.382667e-10, 1.352419e-10, 
    1.35728e-10, 1.354384e-10, 1.343839e-10, 1.377702e-10, 1.360263e-10, 
    1.392567e-10, 1.383044e-10, 1.410943e-10, 1.397028e-10, 1.424436e-10, 
    1.436248e-10, 1.447416e-10, 1.460533e-10, 1.351751e-10, 1.348083e-10, 
    1.354656e-10, 1.363781e-10, 1.372279e-10, 1.383624e-10, 1.384788e-10, 
    1.38692e-10, 1.392453e-10, 1.397114e-10, 1.387595e-10, 1.398284e-10, 
    1.358409e-10, 1.379222e-10, 1.346697e-10, 1.356444e-10, 1.363242e-10, 
    1.360257e-10, 1.375797e-10, 1.379475e-10, 1.394478e-10, 1.38671e-10, 
    1.433327e-10, 1.412592e-10, 1.470566e-10, 1.454227e-10, 1.346802e-10, 
    1.351739e-10, 1.369002e-10, 1.360772e-10, 1.384383e-10, 1.390231e-10, 
    1.394995e-10, 1.4011e-10, 1.40176e-10, 1.405385e-10, 1.399447e-10, 
    1.40515e-10, 1.383648e-10, 1.393233e-10, 1.367022e-10, 1.373375e-10, 
    1.37045e-10, 1.367246e-10, 1.377149e-10, 1.387745e-10, 1.387971e-10, 
    1.391379e-10, 1.40101e-10, 1.384479e-10, 1.436017e-10, 1.40406e-10, 
    1.357134e-10, 1.366694e-10, 1.368063e-10, 1.364352e-10, 1.389644e-10, 
    1.380449e-10, 1.405296e-10, 1.398556e-10, 1.40961e-10, 1.404111e-10, 
    1.403303e-10, 1.39626e-10, 1.391886e-10, 1.38087e-10, 1.371944e-10, 
    1.36489e-10, 1.366528e-10, 1.374284e-10, 1.388394e-10, 1.40182e-10, 
    1.398872e-10, 1.408768e-10, 1.382663e-10, 1.393575e-10, 1.389352e-10, 
    1.400379e-10, 1.376282e-10, 1.396788e-10, 1.371069e-10, 1.373312e-10, 
    1.380267e-10, 1.394317e-10, 1.397436e-10, 1.400772e-10, 1.398713e-10, 
    1.388753e-10, 1.387125e-10, 1.380097e-10, 1.378161e-10, 1.372824e-10, 
    1.368414e-10, 1.372443e-10, 1.376681e-10, 1.388757e-10, 1.399693e-10, 
    1.411673e-10, 1.414614e-10, 1.428705e-10, 1.417229e-10, 1.436197e-10, 
    1.420063e-10, 1.448059e-10, 1.397981e-10, 1.419588e-10, 1.380584e-10, 
    1.384755e-10, 1.392319e-10, 1.409758e-10, 1.400327e-10, 1.41136e-10, 
    1.387062e-10, 1.374552e-10, 1.371326e-10, 1.365319e-10, 1.371463e-10, 
    1.370963e-10, 1.376856e-10, 1.374961e-10, 1.389159e-10, 1.381522e-10, 
    1.403282e-10, 1.411273e-10, 1.433981e-10, 1.448006e-10, 1.462365e-10, 
    1.468731e-10, 1.470672e-10, 1.471484e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24572.8, 24593.05, 24589.08, 24605.65, 24596.42, 24607.33, 24576.87, 
    24593.86, 24582.98, 24574.6, 24638.56, 24606.4, 24672.95, 24651.7, 
    24705.54, 24669.61, 24712.92, 24704.49, 24730.11, 24722.7, 24756.31, 
    24733.55, 24774.2, 24750.83, 24754.45, 24732.81, 24612.8, 24634.51, 
    24611.52, 24614.59, 24613.21, 24596.61, 24588.35, 24571.27, 24574.35, 
    24586.91, 24615.98, 24606.01, 24631.29, 24630.71, 24659.47, 24646.41, 
    24695.72, 24681.6, 24723, 24712.42, 24722.51, 24719.44, 24722.54, 
    24707.07, 24713.67, 24700.16, 24648.85, 24663.75, 24619.88, 24594.27, 
    24577.61, 24565.96, 24567.6, 24570.73, 24586.98, 24602.5, 24614.5, 
    24622.61, 24630.63, 24655.27, 24668.54, 24698.61, 24693.14, 24702.42, 
    24711.37, 24726.6, 24724.08, 24730.85, 24702.17, 24721.13, 24690.04, 
    24698.44, 24632.82, 24608.69, 24598.6, 24589.84, 24568.86, 24583.3, 
    24577.58, 24591.24, 24600.02, 24595.67, 24622.83, 24612.18, 24669.34, 
    24644.36, 24710.32, 24694.26, 24714.21, 24703.98, 24721.59, 24705.72, 
    24733.38, 24739.55, 24735.32, 24751.58, 24704.85, 24722.51, 24595.54, 
    24596.25, 24599.56, 24585.11, 24584.23, 24571.18, 24582.79, 24587.77, 
    24600.53, 24608.15, 24615.46, 24631.68, 24650.04, 24676.28, 24695.29, 
    24708.23, 24700.27, 24707.29, 24699.45, 24695.8, 24737.25, 24713.73, 
    24749.23, 24747.23, 24731.01, 24747.46, 24596.75, 24592.68, 24578.68, 
    24589.62, 24569.77, 24580.83, 24587.25, 24612.4, 24618.01, 24623.25, 
    24633.62, 24647.08, 24671.1, 24692.27, 24711.89, 24710.44, 24710.96, 
    24715.39, 24704.44, 24717.2, 24719.36, 24713.73, 24746.96, 24737.36, 
    24747.19, 24740.92, 24594, 24600.87, 24597.15, 24604.15, 24599.22, 
    24621.37, 24628.09, 24660.04, 24646.81, 24667.95, 24648.94, 24652.28, 
    24668.65, 24649.96, 24691.1, 24663.08, 24715.57, 24687.13, 24717.38, 
    24711.81, 24721.04, 24729.39, 24740.05, 24759.96, 24755.31, 24772.21, 
    24611.2, 24620.27, 24619.47, 24629.03, 24636.13, 24651.7, 24677.17, 
    24667.51, 24685.2, 24688.75, 24661.91, 24678.41, 24626.39, 24634.62, 
    24629.71, 24611.91, 24669.73, 24639.69, 24695.61, 24679.06, 24728.2, 
    24703.44, 24752.76, 24774.66, 24795.74, 24820.79, 24625.26, 24619.05, 
    24630.17, 24645.7, 24660.32, 24680.06, 24682.07, 24685.77, 24695.41, 
    24703.59, 24686.94, 24705.65, 24636.54, 24672.38, 24616.72, 24633.2, 
    24644.78, 24639.68, 24666.42, 24672.82, 24698.96, 24685.4, 24769.21, 
    24731.17, 24840.08, 24808.77, 24616.89, 24625.24, 24654.66, 24640.56, 
    24681.37, 24691.53, 24699.86, 24710.63, 24711.8, 24718.25, 24707.71, 
    24717.83, 24680.1, 24696.77, 24651.26, 24662.21, 24657.16, 24651.64, 
    24668.77, 24687.2, 24687.59, 24693.53, 24710.48, 24681.54, 24774.23, 
    24715.89, 24634.37, 24650.7, 24653.05, 24646.68, 24690.5, 24674.53, 
    24718.09, 24706.13, 24725.8, 24715.98, 24714.54, 24702.09, 24694.42, 
    24675.26, 24659.74, 24647.6, 24650.41, 24663.79, 24688.33, 24711.91, 
    24706.69, 24724.29, 24678.4, 24697.38, 24690, 24709.36, 24667.26, 
    24703.02, 24658.22, 24662.11, 24674.21, 24698.68, 24704.16, 24710.05, 
    24706.41, 24688.96, 24686.12, 24673.91, 24670.53, 24661.26, 24653.65, 
    24660.6, 24667.95, 24688.96, 24708.14, 24729.51, 24734.82, 24760.63, 
    24739.6, 24774.57, 24744.76, 24796.97, 24705.12, 24743.89, 24674.76, 
    24682.02, 24695.18, 24726.07, 24709.26, 24728.95, 24686.01, 24664.26, 
    24658.67, 24648.34, 24658.91, 24658.04, 24668.26, 24664.96, 24689.66, 
    24676.41, 24714.51, 24728.79, 24770.42, 24796.86, 24824.3, 24836.53, 
    24840.28, 24841.86 ;

 GC_ICE1 =
  17680.35, 17712.78, 17706.42, 17732.96, 17718.19, 17735.64, 17686.87, 
    17714.08, 17696.66, 17683.24, 17785.63, 17734.16, 17840.63, 17806.65, 
    17892.65, 17835.3, 17904.42, 17890.96, 17931.83, 17920.01, 17973.63, 
    17937.32, 18002.16, 17964.89, 17970.66, 17936.14, 17744.41, 17779.16, 
    17742.37, 17747.28, 17745.07, 17718.49, 17705.26, 17677.9, 17682.83, 
    17702.95, 17749.5, 17733.54, 17774, 17773.08, 17819.08, 17798.19, 
    17876.99, 17854.46, 17920.5, 17903.62, 17919.71, 17914.81, 17919.77, 
    17895.08, 17905.61, 17884.07, 17802.09, 17825.93, 17755.73, 17714.73, 
    17688.06, 17669.4, 17672.02, 17677.04, 17703.06, 17727.92, 17747.13, 
    17760.11, 17772.95, 17812.36, 17833.59, 17881.58, 17872.86, 17887.67, 
    17901.95, 17926.24, 17922.21, 17933.01, 17887.27, 17917.52, 17867.91, 
    17881.32, 17776.46, 17737.83, 17721.67, 17707.64, 17674.04, 17697.17, 
    17688.02, 17709.89, 17723.94, 17716.97, 17760.46, 17743.42, 17834.85, 
    17794.91, 17900.28, 17874.65, 17906.48, 17890.15, 17918.25, 17892.94, 
    17937.05, 17946.91, 17940.14, 17966.09, 17891.55, 17919.71, 17716.78, 
    17717.91, 17723.21, 17700.07, 17698.66, 17677.77, 17696.35, 17704.33, 
    17724.76, 17736.97, 17748.67, 17774.62, 17804.01, 17845.96, 17876.29, 
    17896.94, 17884.24, 17895.44, 17882.93, 17877.1, 17943.24, 17905.71, 
    17962.34, 17959.15, 17933.27, 17959.51, 17718.71, 17712.19, 17689.77, 
    17707.29, 17675.51, 17693.22, 17703.5, 17743.77, 17752.76, 17761.14, 
    17777.73, 17799.26, 17837.68, 17871.47, 17902.78, 17900.46, 17901.28, 
    17908.36, 17890.89, 17911.25, 17914.7, 17905.7, 17958.72, 17943.4, 
    17959.08, 17949.09, 17714.31, 17725.3, 17719.35, 17730.56, 17722.66, 
    17758.12, 17768.88, 17819.99, 17798.83, 17832.64, 17802.24, 17807.58, 
    17833.76, 17803.86, 17869.6, 17824.86, 17908.64, 17863.27, 17911.53, 
    17902.64, 17917.38, 17930.69, 17947.7, 17979.44, 17972.03, 17998.97, 
    17741.84, 17756.37, 17755.09, 17770.38, 17781.75, 17806.65, 17847.39, 
    17831.94, 17860.19, 17865.87, 17822.98, 17849.36, 17766.16, 17779.32, 
    17771.47, 17742.98, 17835.49, 17787.44, 17876.8, 17850.4, 17928.79, 
    17889.29, 17967.96, 18002.89, 18036.49, 18076.38, 17764.36, 17754.42, 
    17772.21, 17797.06, 17820.43, 17852, 17855.21, 17861.1, 17876.48, 
    17889.53, 17862.97, 17892.82, 17782.4, 17839.73, 17750.68, 17777.06, 
    17795.58, 17787.43, 17830.19, 17840.43, 17882.14, 17860.52, 17994.19, 
    17933.53, 18107.03, 18057.26, 17750.96, 17764.32, 17811.39, 17788.83, 
    17854.09, 17870.29, 17883.59, 17900.77, 17902.63, 17912.91, 17896.1, 
    17912.25, 17852.06, 17878.66, 17805.94, 17823.46, 17815.38, 17806.56, 
    17833.94, 17863.39, 17864.01, 17873.49, 17900.52, 17854.35, 18002.21, 
    17909.16, 17778.92, 17805.05, 17808.8, 17798.62, 17868.66, 17843.15, 
    17912.66, 17893.59, 17924.97, 17909.29, 17907, 17887.13, 17874.9, 
    17844.33, 17819.51, 17800.1, 17804.59, 17825.98, 17865.19, 17902.8, 
    17894.48, 17922.56, 17849.35, 17879.62, 17867.85, 17898.73, 17831.53, 
    17888.63, 17817.09, 17823.29, 17842.65, 17881.7, 17890.44, 17899.84, 
    17894.03, 17866.19, 17861.67, 17842.17, 17836.77, 17821.94, 17809.77, 
    17820.88, 17832.64, 17866.2, 17896.8, 17930.88, 17939.35, 17980.52, 
    17946.98, 18002.74, 17955.21, 18038.45, 17891.98, 17953.83, 17843.53, 
    17855.12, 17876.11, 17925.4, 17898.58, 17929.99, 17861.49, 17826.73, 
    17817.8, 17801.27, 17818.18, 17816.79, 17833.13, 17827.86, 17867.31, 
    17846.16, 17906.95, 17929.74, 17996.13, 18038.29, 18081.95, 18101.39, 
    18107.35, 18109.85 ;

 GC_LIQ1 =
  5232.711, 5234.74, 5234.342, 5236.003, 5235.078, 5236.171, 5233.119, 
    5234.821, 5233.731, 5232.892, 5239.312, 5236.078, 5242.792, 5240.64, 
    5246.142, 5242.454, 5246.903, 5246.033, 5248.677, 5247.912, 5251.378, 
    5249.032, 5253.228, 5250.812, 5251.186, 5248.956, 5236.72, 5238.904, 
    5236.592, 5236.9, 5236.762, 5235.097, 5234.27, 5232.558, 5232.866, 
    5234.125, 5237.039, 5236.04, 5238.579, 5238.521, 5241.427, 5240.105, 
    5245.129, 5243.674, 5247.943, 5246.851, 5247.892, 5247.575, 5247.896, 
    5246.299, 5246.98, 5245.587, 5240.352, 5241.86, 5237.43, 5234.862, 
    5233.193, 5232.026, 5232.19, 5232.504, 5234.132, 5235.688, 5236.891, 
    5237.704, 5238.512, 5241.001, 5242.345, 5245.427, 5244.863, 5245.82, 
    5246.743, 5248.314, 5248.054, 5248.753, 5245.794, 5247.75, 5244.543, 
    5245.41, 5238.733, 5236.308, 5235.296, 5234.418, 5232.316, 5233.763, 
    5233.19, 5234.559, 5235.438, 5235.002, 5237.726, 5236.658, 5242.426, 
    5239.898, 5246.635, 5244.979, 5247.037, 5245.98, 5247.797, 5246.161, 
    5249.014, 5249.647, 5249.214, 5250.89, 5246.071, 5247.892, 5234.99, 
    5235.061, 5235.393, 5233.944, 5233.856, 5232.549, 5233.711, 5234.211, 
    5235.49, 5236.254, 5236.987, 5238.618, 5240.473, 5243.129, 5245.085, 
    5246.419, 5245.599, 5246.323, 5245.514, 5245.137, 5249.41, 5246.986, 
    5250.646, 5250.44, 5248.77, 5250.463, 5235.111, 5234.703, 5233.3, 
    5234.396, 5232.408, 5233.516, 5234.159, 5236.681, 5237.243, 5237.769, 
    5238.814, 5240.173, 5242.605, 5244.773, 5246.797, 5246.647, 5246.7, 
    5247.158, 5246.028, 5247.345, 5247.568, 5246.986, 5250.413, 5249.421, 
    5250.436, 5249.789, 5234.835, 5235.524, 5235.151, 5235.854, 5235.358, 
    5237.58, 5238.255, 5241.484, 5240.146, 5242.285, 5240.361, 5240.699, 
    5242.356, 5240.464, 5244.652, 5241.793, 5247.176, 5244.244, 5247.363, 
    5246.789, 5247.741, 5248.603, 5249.698, 5251.755, 5251.274, 5253.021, 
    5236.56, 5237.47, 5237.389, 5238.35, 5239.067, 5240.641, 5243.219, 
    5242.241, 5244.045, 5244.411, 5241.674, 5243.345, 5238.084, 5238.915, 
    5238.419, 5236.631, 5242.466, 5239.427, 5245.118, 5243.412, 5248.479, 
    5245.925, 5251.011, 5253.274, 5255.456, 5258.074, 5237.97, 5237.348, 
    5238.465, 5240.034, 5241.513, 5243.515, 5243.723, 5244.104, 5245.097, 
    5245.94, 5244.224, 5246.153, 5239.108, 5242.734, 5237.113, 5238.771, 
    5239.94, 5239.426, 5242.13, 5242.779, 5245.463, 5244.066, 5252.711, 
    5248.786, 5260.12, 5256.808, 5237.131, 5237.968, 5240.94, 5239.514, 
    5243.65, 5244.697, 5245.557, 5246.667, 5246.788, 5247.453, 5246.365, 
    5247.409, 5243.52, 5245.238, 5240.596, 5241.705, 5241.193, 5240.635, 
    5242.368, 5244.251, 5244.292, 5244.904, 5246.651, 5243.667, 5253.23, 
    5247.209, 5238.889, 5240.539, 5240.777, 5240.133, 5244.591, 5242.952, 
    5247.437, 5246.203, 5248.232, 5247.218, 5247.07, 5245.786, 5244.995, 
    5243.026, 5241.454, 5240.226, 5240.51, 5241.864, 5244.367, 5246.798, 
    5246.261, 5248.077, 5243.344, 5245.3, 5244.539, 5246.535, 5242.215, 
    5245.882, 5241.301, 5241.694, 5242.919, 5245.434, 5245.999, 5246.607, 
    5246.231, 5244.432, 5244.14, 5242.889, 5242.547, 5241.608, 5240.838, 
    5241.542, 5242.286, 5244.433, 5246.41, 5248.615, 5249.163, 5251.824, 
    5249.652, 5253.265, 5250.185, 5255.583, 5246.099, 5250.096, 5242.975, 
    5243.717, 5245.073, 5248.26, 5246.526, 5248.557, 5244.128, 5241.911, 
    5241.346, 5240.3, 5241.37, 5241.282, 5242.316, 5241.983, 5244.504, 
    5243.142, 5247.066, 5248.541, 5252.836, 5255.573, 5258.445, 5259.743, 
    5260.141, 5260.309 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.756585e-09, 8.795193e-09, 8.787688e-09, 8.818827e-09, 8.801554e-09, 
    8.821944e-09, 8.764413e-09, 8.796724e-09, 8.776098e-09, 8.760061e-09, 
    8.87926e-09, 8.820217e-09, 8.940603e-09, 8.902943e-09, 8.997554e-09, 
    8.934742e-09, 9.01022e-09, 8.995744e-09, 9.03932e-09, 9.026836e-09, 
    9.082572e-09, 9.045082e-09, 9.111468e-09, 9.073621e-09, 9.079541e-09, 
    9.043845e-09, 8.8321e-09, 8.871908e-09, 8.829741e-09, 8.835419e-09, 
    8.832871e-09, 8.80191e-09, 8.786307e-09, 8.753635e-09, 8.759567e-09, 
    8.783564e-09, 8.83797e-09, 8.819503e-09, 8.866051e-09, 8.865e-09, 
    8.916823e-09, 8.893457e-09, 8.980567e-09, 8.955808e-09, 9.027357e-09, 
    9.009362e-09, 9.026511e-09, 9.021312e-09, 9.026579e-09, 9.000188e-09, 
    9.011495e-09, 8.988273e-09, 8.897833e-09, 8.924411e-09, 8.845142e-09, 
    8.797481e-09, 8.76583e-09, 8.743369e-09, 8.746544e-09, 8.752597e-09, 
    8.783704e-09, 8.812955e-09, 8.835245e-09, 8.850156e-09, 8.864848e-09, 
    8.909318e-09, 8.93286e-09, 8.985571e-09, 8.976061e-09, 8.992175e-09, 
    9.007572e-09, 9.033421e-09, 9.029167e-09, 9.040555e-09, 8.991751e-09, 
    9.024185e-09, 8.970643e-09, 8.985286e-09, 8.868836e-09, 8.824486e-09, 
    8.805629e-09, 8.78913e-09, 8.748986e-09, 8.776707e-09, 8.765779e-09, 
    8.791781e-09, 8.808303e-09, 8.800131e-09, 8.850564e-09, 8.830956e-09, 
    8.934255e-09, 8.889759e-09, 9.005777e-09, 8.978013e-09, 9.012431e-09, 
    8.994869e-09, 9.024961e-09, 8.997878e-09, 9.044794e-09, 9.055013e-09, 
    9.048028e-09, 9.07485e-09, 8.996377e-09, 9.02651e-09, 8.799902e-09, 
    8.801234e-09, 8.807444e-09, 8.780151e-09, 8.778481e-09, 8.753473e-09, 
    8.775726e-09, 8.785202e-09, 8.80926e-09, 8.82349e-09, 8.837017e-09, 
    8.866762e-09, 8.89998e-09, 8.946435e-09, 8.979812e-09, 9.002187e-09, 
    8.988468e-09, 9.00058e-09, 8.98704e-09, 8.980694e-09, 9.051184e-09, 
    9.0116e-09, 9.070993e-09, 9.067707e-09, 9.040826e-09, 9.068077e-09, 
    8.802171e-09, 8.794502e-09, 8.767875e-09, 8.788713e-09, 8.750749e-09, 
    8.771998e-09, 8.784216e-09, 8.831365e-09, 8.841726e-09, 8.851331e-09, 
    8.870304e-09, 8.894652e-09, 8.937367e-09, 8.974536e-09, 9.008469e-09, 
    9.005982e-09, 9.006857e-09, 9.014437e-09, 8.995661e-09, 9.01752e-09, 
    9.021188e-09, 9.011596e-09, 9.067266e-09, 9.051363e-09, 9.067636e-09, 
    9.057282e-09, 8.796994e-09, 8.809899e-09, 8.802925e-09, 8.816038e-09, 
    8.8068e-09, 8.847875e-09, 8.860192e-09, 8.917825e-09, 8.894173e-09, 
    8.931816e-09, 8.897997e-09, 8.90399e-09, 8.933042e-09, 8.899825e-09, 
    8.972485e-09, 8.92322e-09, 9.014731e-09, 8.965531e-09, 9.017815e-09, 
    9.008321e-09, 9.02404e-09, 9.038118e-09, 9.055833e-09, 9.088511e-09, 
    9.080944e-09, 9.108275e-09, 8.829137e-09, 8.845873e-09, 8.844402e-09, 
    8.861918e-09, 8.874872e-09, 8.902953e-09, 8.947992e-09, 8.931056e-09, 
    8.962149e-09, 8.968391e-09, 8.921153e-09, 8.950155e-09, 8.857076e-09, 
    8.872113e-09, 8.863161e-09, 8.830456e-09, 8.934957e-09, 8.881324e-09, 
    8.980364e-09, 8.951308e-09, 9.03611e-09, 8.993934e-09, 9.076778e-09, 
    9.11219e-09, 9.145526e-09, 9.184478e-09, 8.85501e-09, 8.843637e-09, 
    8.864002e-09, 8.892176e-09, 8.918321e-09, 8.95308e-09, 8.956637e-09, 
    8.963148e-09, 8.980017e-09, 8.994199e-09, 8.965206e-09, 8.997755e-09, 
    8.875597e-09, 8.939613e-09, 8.839336e-09, 8.869528e-09, 8.890516e-09, 
    8.881311e-09, 8.929121e-09, 8.940389e-09, 8.98618e-09, 8.962509e-09, 
    9.103449e-09, 9.04109e-09, 9.214142e-09, 9.165777e-09, 8.839663e-09, 
    8.854971e-09, 8.908249e-09, 8.8829e-09, 8.955401e-09, 8.973248e-09, 
    8.987757e-09, 9.006302e-09, 9.008306e-09, 9.019295e-09, 9.001288e-09, 
    9.018583e-09, 8.953154e-09, 8.982393e-09, 8.902161e-09, 8.921687e-09, 
    8.912704e-09, 8.902851e-09, 8.933263e-09, 8.965662e-09, 8.966357e-09, 
    8.976746e-09, 9.006017e-09, 8.955695e-09, 9.111494e-09, 9.015269e-09, 
    8.871664e-09, 8.901148e-09, 8.905363e-09, 8.893941e-09, 8.971458e-09, 
    8.94337e-09, 9.019026e-09, 8.99858e-09, 9.032083e-09, 9.015434e-09, 
    9.012984e-09, 8.991602e-09, 8.978289e-09, 8.944657e-09, 8.917294e-09, 
    8.895597e-09, 8.900643e-09, 8.924476e-09, 8.967644e-09, 9.008486e-09, 
    8.99954e-09, 9.029536e-09, 8.950144e-09, 8.983433e-09, 8.970566e-09, 
    9.004117e-09, 8.930606e-09, 8.993198e-09, 8.914606e-09, 8.921496e-09, 
    8.942813e-09, 8.98569e-09, 8.995179e-09, 9.005308e-09, 8.999058e-09, 
    8.968741e-09, 8.963775e-09, 8.942295e-09, 8.936363e-09, 8.919996e-09, 
    8.906446e-09, 8.918827e-09, 8.931828e-09, 8.968755e-09, 9.002033e-09, 
    9.038318e-09, 9.047199e-09, 9.089592e-09, 9.055081e-09, 9.112029e-09, 
    9.063609e-09, 9.147431e-09, 8.996828e-09, 9.062188e-09, 8.943783e-09, 
    8.956539e-09, 8.979608e-09, 9.032526e-09, 9.003959e-09, 9.037369e-09, 
    8.963581e-09, 8.925298e-09, 8.915395e-09, 8.896916e-09, 8.915817e-09, 
    8.91428e-09, 8.932367e-09, 8.926555e-09, 8.96998e-09, 8.946654e-09, 
    9.012923e-09, 9.037106e-09, 9.10541e-09, 9.147281e-09, 9.189909e-09, 
    9.208728e-09, 9.214456e-09, 9.216851e-09 ;

 H2OCAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  6.177402, 6.205632, 6.200137, 6.222954, 6.210289, 6.22524, 6.183118, 
    6.206756, 6.191658, 6.179939, 6.267385, 6.223972, 6.31266, 6.284832, 
    6.354875, 6.308327, 6.364285, 6.353526, 6.385933, 6.376639, 6.423027, 
    6.390226, 6.444653, 6.416328, 6.420756, 6.389305, 6.23269, 6.261971, 
    6.230959, 6.235128, 6.233256, 6.210552, 6.199131, 6.175246, 6.179577, 
    6.197122, 6.237004, 6.223445, 6.257643, 6.25687, 6.295077, 6.277833, 
    6.34226, 6.323907, 6.377027, 6.363643, 6.376398, 6.372529, 6.376449, 
    6.356827, 6.36523, 6.347979, 6.281061, 6.300684, 6.242271, 6.207314, 
    6.184154, 6.167755, 6.170072, 6.17449, 6.197224, 6.218643, 6.234998, 
    6.245953, 6.256759, 6.289546, 6.306933, 6.345977, 6.338917, 6.350878, 
    6.362312, 6.381542, 6.378374, 6.386856, 6.35056, 6.37467, 6.334898, 
    6.345762, 6.259711, 6.227101, 6.213283, 6.201193, 6.171854, 6.192107, 
    6.184118, 6.203131, 6.215233, 6.209245, 6.246253, 6.23185, 6.307964, 
    6.27511, 6.360978, 6.340366, 6.365924, 6.352874, 6.375246, 6.355109, 
    6.390013, 6.402422, 6.392425, 6.417244, 6.353994, 6.3764, 6.209078, 
    6.210055, 6.214603, 6.194624, 6.193403, 6.175128, 6.191386, 6.198319, 
    6.215934, 6.22637, 6.2363, 6.258168, 6.282648, 6.316973, 6.341701, 
    6.35831, 6.348121, 6.357116, 6.347062, 6.342352, 6.399561, 6.365309, 
    6.414361, 6.411904, 6.387058, 6.412181, 6.21074, 6.205123, 6.185648, 
    6.200885, 6.17314, 6.188663, 6.1976, 6.232153, 6.239758, 6.246819, 
    6.260775, 6.278715, 6.310263, 6.337789, 6.362978, 6.36113, 6.36178, 
    6.367416, 6.353463, 6.369709, 6.372439, 6.365304, 6.411575, 6.399692, 
    6.411852, 6.404115, 6.206948, 6.216403, 6.211293, 6.220905, 6.214133, 
    6.244282, 6.253339, 6.295821, 6.278362, 6.306159, 6.281181, 6.285604, 
    6.307073, 6.282529, 6.336272, 6.29981, 6.367635, 6.331121, 6.369928, 
    6.362869, 6.374558, 6.38504, 6.403032, 6.427464, 6.421803, 6.442258, 
    6.230514, 6.242809, 6.241724, 6.254603, 6.26414, 6.284837, 6.318123, 
    6.305593, 6.328605, 6.333231, 6.298274, 6.319726, 6.251044, 6.262112, 
    6.255519, 6.231484, 6.308482, 6.268896, 6.34211, 6.320577, 6.383545, 
    6.352185, 6.418687, 6.445199, 6.470194, 6.499485, 6.249523, 6.241162, 
    6.256135, 6.276893, 6.296184, 6.321889, 6.324522, 6.329346, 6.341851, 
    6.352377, 6.330874, 6.355017, 6.264685, 6.311924, 6.238004, 6.26021, 
    6.275667, 6.268881, 6.304161, 6.312494, 6.346427, 6.328871, 6.438652, 
    6.387259, 6.521831, 6.485416, 6.238243, 6.249493, 6.288749, 6.270051, 
    6.323606, 6.336832, 6.347594, 6.361371, 6.362857, 6.371029, 6.357642, 
    6.370499, 6.321944, 6.343615, 6.284251, 6.29867, 6.292034, 6.28476, 
    6.307224, 6.331213, 6.331723, 6.339427, 6.361177, 6.323823, 6.444688, 
    6.368052, 6.261775, 6.283512, 6.286616, 6.278188, 6.335505, 6.314702, 
    6.37083, 6.35563, 6.380545, 6.368157, 6.366336, 6.350449, 6.340571, 
    6.315655, 6.295425, 6.27941, 6.283131, 6.300732, 6.332682, 6.362994, 
    6.356347, 6.378649, 6.319714, 6.344388, 6.334846, 6.359745, 6.305261, 
    6.351651, 6.293437, 6.298527, 6.314289, 6.346067, 6.353105, 6.360631, 
    6.355986, 6.333493, 6.329811, 6.313904, 6.309519, 6.297419, 6.287414, 
    6.296556, 6.306166, 6.333501, 6.358199, 6.38519, 6.391804, 6.428282, 
    6.402479, 6.44509, 6.408862, 6.47164, 6.35434, 6.407791, 6.315005, 
    6.324448, 6.341553, 6.380882, 6.359628, 6.384487, 6.329667, 6.301341, 
    6.294021, 6.280383, 6.294333, 6.293197, 6.306561, 6.302265, 6.33441, 
    6.317131, 6.366292, 6.384289, 6.440114, 6.471518, 6.503567, 6.517746, 
    6.522065, 6.523871,
  3.94925, 3.968676, 3.964894, 3.980599, 3.971881, 3.982172, 3.953182, 
    3.96945, 3.959059, 3.950994, 4.011191, 3.9813, 4.041689, 4.023084, 
    4.069917, 4.038793, 4.07621, 4.069013, 4.090688, 4.084471, 4.112349, 
    4.093559, 4.126805, 4.10787, 4.11083, 4.092943, 3.987301, 4.007463, 
    3.986109, 3.988979, 3.98769, 3.972062, 3.964204, 3.947765, 3.950745, 
    3.962819, 3.990271, 3.980936, 4.004479, 4.003946, 4.029933, 4.018382, 
    4.061479, 4.049207, 4.08473, 4.075779, 4.08431, 4.081721, 4.084344, 
    4.07122, 4.07684, 4.065303, 4.020564, 4.033681, 3.993896, 3.969836, 
    3.953895, 3.94261, 3.944204, 3.947245, 3.96289, 3.977631, 3.988889, 
    3.996431, 4.00387, 4.026238, 4.03786, 4.063966, 4.059243, 4.067243, 
    4.074889, 4.087751, 4.085632, 4.091306, 4.067029, 4.083155, 4.056555, 
    4.06382, 4.005908, 3.983453, 3.973943, 3.965621, 3.945431, 3.959368, 
    3.95387, 3.966954, 3.975284, 3.971162, 3.996637, 3.986722, 4.038549, 
    4.016507, 4.073997, 4.060212, 4.077304, 4.068576, 4.08354, 4.070071, 
    4.093418, 4.098579, 4.095031, 4.10848, 4.069325, 4.084311, 3.971047, 
    3.97172, 3.97485, 3.961101, 3.96026, 3.947684, 3.958872, 3.963643, 
    3.975766, 3.98295, 3.989786, 4.004841, 4.021625, 4.044571, 4.061104, 
    4.072211, 4.065398, 4.071413, 4.064689, 4.06154, 4.09667, 4.076893, 
    4.106554, 4.104912, 4.091441, 4.105097, 3.972191, 3.968325, 3.954923, 
    3.965409, 3.946315, 3.956997, 3.963149, 3.986932, 3.992165, 3.997027, 
    4.006635, 4.018989, 4.040085, 4.058489, 4.075333, 4.074097, 4.074533, 
    4.078302, 4.06897, 4.079835, 4.081662, 4.07689, 4.104692, 4.096756, 
    4.104877, 4.099708, 3.969581, 3.976089, 3.972572, 3.979188, 3.974527, 
    3.995282, 4.001517, 4.030432, 4.018746, 4.037342, 4.020644, 4.0236, 
    4.037955, 4.021544, 4.057476, 4.033099, 4.078449, 4.054033, 4.079982, 
    4.07526, 4.083079, 4.090091, 4.098985, 4.115313, 4.111528, 4.125203, 
    3.985802, 3.994267, 3.993519, 4.002386, 4.008953, 4.023087, 4.045339, 
    4.036962, 4.052347, 4.055441, 4.032069, 4.046412, 3.999936, 4.007557, 
    4.003017, 3.986471, 4.038895, 4.012228, 4.061378, 4.04698, 4.089091, 
    4.068117, 4.109446, 4.127172, 4.143886, 4.163485, 3.998888, 3.993132, 
    4.003441, 4.017735, 4.030672, 4.047858, 4.049617, 4.052843, 4.061204, 
    4.068244, 4.053866, 4.070009, 4.009332, 4.041196, 3.990959, 4.006248, 
    4.016891, 4.012218, 4.036004, 4.041575, 4.064266, 4.052525, 4.122796, 
    4.091577, 4.178435, 4.15407, 3.991122, 3.998868, 4.025703, 4.013023, 
    4.049005, 4.057849, 4.065045, 4.074259, 4.075253, 4.080719, 4.071764, 
    4.080364, 4.047894, 4.062384, 4.022695, 4.032334, 4.027897, 4.023036, 
    4.038052, 4.054093, 4.054432, 4.059585, 4.074136, 4.04915, 4.126836, 
    4.078733, 4.007324, 4.022204, 4.024276, 4.018626, 4.056962, 4.043052, 
    4.080585, 4.070419, 4.087083, 4.078798, 4.07758, 4.066954, 4.060349, 
    4.04369, 4.030166, 4.019459, 4.021946, 4.033713, 4.055075, 4.075345, 
    4.0709, 4.085815, 4.046402, 4.062902, 4.056522, 4.073172, 4.03674, 
    4.067764, 4.028836, 4.032238, 4.042776, 4.064026, 4.06873, 4.073765, 
    4.070657, 4.055617, 4.053154, 4.042519, 4.039587, 4.031497, 4.024809, 
    4.030921, 4.037346, 4.055622, 4.072138, 4.090191, 4.094615, 4.115863, 
    4.09862, 4.127105, 4.10289, 4.144858, 4.06956, 4.10217, 4.043254, 
    4.049568, 4.061007, 4.087312, 4.073093, 4.089723, 4.053058, 4.034122, 
    4.029225, 4.02011, 4.029434, 4.028675, 4.037609, 4.034736, 4.056229, 
    4.044675, 4.07755, 4.08959, 4.12377, 4.144773, 4.166212, 4.175701, 
    4.178591, 4.1798,
  3.268149, 3.285393, 3.282035, 3.295979, 3.288238, 3.297376, 3.271639, 
    3.28608, 3.276855, 3.269697, 3.323152, 3.296601, 3.350864, 3.333825, 
    3.376728, 3.348211, 3.382497, 3.3759, 3.395771, 3.390071, 3.415585, 
    3.398404, 3.428849, 3.411477, 3.414192, 3.397839, 3.30193, 3.31984, 
    3.300872, 3.303421, 3.302276, 3.288399, 3.281422, 3.266832, 3.269477, 
    3.280193, 3.304568, 3.296278, 3.317189, 3.316716, 3.340097, 3.329542, 
    3.368996, 3.357751, 3.390308, 3.382102, 3.389923, 3.38755, 3.389954, 
    3.377924, 3.383075, 3.3725, 3.331517, 3.34353, 3.307788, 3.286422, 
    3.272272, 3.262258, 3.263672, 3.266371, 3.280256, 3.293343, 3.303341, 
    3.310039, 3.316648, 3.336712, 3.347356, 3.371274, 3.366947, 3.374278, 
    3.381286, 3.393078, 3.391135, 3.396337, 3.374082, 3.388864, 3.364484, 
    3.371141, 3.318457, 3.298513, 3.290069, 3.282681, 3.26476, 3.27713, 
    3.27225, 3.283864, 3.291259, 3.2876, 3.310223, 3.301416, 3.347988, 
    3.327876, 3.380468, 3.367835, 3.383501, 3.3755, 3.389217, 3.37687, 
    3.398274, 3.402956, 3.399753, 3.412038, 3.376187, 3.389924, 3.287498, 
    3.288095, 3.290874, 3.278668, 3.277921, 3.26676, 3.276689, 3.280924, 
    3.291687, 3.298067, 3.304137, 3.31751, 3.332489, 3.353504, 3.368653, 
    3.378832, 3.372587, 3.3781, 3.371938, 3.369052, 3.401205, 3.383124, 
    3.41027, 3.408765, 3.396461, 3.408934, 3.288513, 3.285081, 3.273185, 
    3.282492, 3.265545, 3.275026, 3.280486, 3.301602, 3.306251, 3.310569, 
    3.319105, 3.330081, 3.349395, 3.366256, 3.381694, 3.380561, 3.38096, 
    3.384415, 3.375861, 3.385821, 3.387496, 3.38312, 3.408563, 3.401284, 
    3.408733, 3.403991, 3.286196, 3.291974, 3.288851, 3.294726, 3.290587, 
    3.309019, 3.314558, 3.340553, 3.329866, 3.346882, 3.331591, 3.334298, 
    3.347443, 3.332415, 3.365327, 3.342995, 3.38455, 3.362172, 3.385956, 
    3.381627, 3.388794, 3.395223, 3.403329, 3.418305, 3.414833, 3.427379, 
    3.300599, 3.308117, 3.307453, 3.31533, 3.321164, 3.333828, 3.354208, 
    3.346534, 3.360628, 3.363463, 3.342053, 3.35519, 3.313153, 3.319924, 
    3.31589, 3.301193, 3.348305, 3.324074, 3.368904, 3.355711, 3.394306, 
    3.375079, 3.412923, 3.429185, 3.444526, 3.46252, 3.312223, 3.307109, 
    3.316267, 3.328968, 3.340774, 3.356515, 3.358127, 3.361083, 3.368744, 
    3.375196, 3.36202, 3.376814, 3.3215, 3.350412, 3.305179, 3.318761, 
    3.328217, 3.324064, 3.345657, 3.35076, 3.37155, 3.360791, 3.425169, 
    3.396585, 3.476254, 3.453875, 3.305324, 3.312204, 3.336223, 3.32478, 
    3.357566, 3.365669, 3.372264, 3.380709, 3.38162, 3.386631, 3.378423, 
    3.386306, 3.356549, 3.369825, 3.333469, 3.342296, 3.338233, 3.333781, 
    3.347533, 3.362228, 3.362539, 3.36726, 3.380594, 3.3577, 3.428875, 
    3.384809, 3.319717, 3.333019, 3.334917, 3.329759, 3.364856, 3.352113, 
    3.386508, 3.377189, 3.392466, 3.38487, 3.383753, 3.374014, 3.36796, 
    3.352697, 3.34031, 3.330506, 3.332784, 3.343559, 3.363127, 3.381704, 
    3.37763, 3.391303, 3.355182, 3.3703, 3.364453, 3.379712, 3.346331, 
    3.374754, 3.339092, 3.342208, 3.35186, 3.37133, 3.375642, 3.380256, 
    3.377408, 3.363624, 3.361368, 3.351624, 3.348939, 3.34153, 3.335405, 
    3.341001, 3.346886, 3.363628, 3.378765, 3.395315, 3.399372, 3.418809, 
    3.402993, 3.429122, 3.406907, 3.445417, 3.376401, 3.406248, 3.352298, 
    3.358082, 3.368563, 3.392674, 3.37964, 3.394885, 3.361279, 3.343932, 
    3.339449, 3.331102, 3.33964, 3.338945, 3.347127, 3.344496, 3.364185, 
    3.3536, 3.383726, 3.394764, 3.426064, 3.44534, 3.465026, 3.473742, 
    3.476397, 3.477508,
  2.990303, 3.006691, 3.003499, 3.016756, 3.009396, 3.018085, 2.993618, 
    3.007343, 2.998576, 2.991774, 3.042611, 3.017348, 3.069009, 3.052777, 
    3.093672, 3.06648, 3.099176, 3.092882, 3.111847, 3.106405, 3.130761, 
    3.114361, 3.143439, 3.126837, 3.129431, 3.113822, 3.022417, 3.039459, 
    3.02141, 3.023835, 3.022747, 3.009548, 3.002915, 2.989051, 2.991564, 
    3.001748, 3.024926, 3.017042, 3.036937, 3.036487, 3.05875, 3.048697, 
    3.086297, 3.075575, 3.106632, 3.0988, 3.106264, 3.103999, 3.106294, 
    3.094813, 3.099728, 3.089639, 3.050579, 3.062021, 3.02799, 3.007668, 
    2.99422, 2.984706, 2.98605, 2.988613, 3.001807, 3.01425, 3.023759, 
    3.030133, 3.036422, 3.055525, 3.065667, 3.08847, 3.084343, 3.091335, 
    3.098022, 3.109276, 3.107421, 3.112387, 3.091148, 3.105253, 3.081995, 
    3.088343, 3.038142, 3.019167, 3.011136, 3.004112, 2.987083, 2.998836, 
    2.994199, 3.005238, 3.012269, 3.008789, 3.030307, 3.021928, 3.066269, 
    3.047111, 3.097241, 3.085189, 3.100135, 3.092501, 3.10559, 3.093808, 
    3.114236, 3.118699, 3.115649, 3.127373, 3.093156, 3.106265, 3.008692, 
    3.009259, 3.011902, 3.000298, 2.999588, 2.988983, 2.998418, 3.002443, 
    3.012676, 3.018742, 3.024517, 3.037243, 3.051504, 3.071526, 3.08597, 
    3.09568, 3.089723, 3.094982, 3.089103, 3.08635, 3.117027, 3.099775, 
    3.125685, 3.124247, 3.112506, 3.124409, 3.009658, 3.006394, 2.995087, 
    3.003933, 2.987829, 2.996837, 3.002026, 3.022105, 3.026528, 3.030636, 
    3.03876, 3.049211, 3.06761, 3.083684, 3.098411, 3.09733, 3.09771, 
    3.101008, 3.092846, 3.102349, 3.103947, 3.099771, 3.124054, 3.117102, 
    3.124216, 3.119688, 3.007455, 3.012948, 3.009979, 3.015565, 3.011629, 
    3.029161, 3.034432, 3.059185, 3.049006, 3.065215, 3.050649, 3.053226, 
    3.065749, 3.051434, 3.082798, 3.061511, 3.101136, 3.079789, 3.102477, 
    3.098347, 3.105187, 3.111324, 3.119055, 3.133361, 3.130044, 3.142034, 
    3.021151, 3.028303, 3.027672, 3.035167, 3.04072, 3.052779, 3.072197, 
    3.064884, 3.078318, 3.081021, 3.060614, 3.073133, 3.033096, 3.03954, 
    3.0357, 3.021716, 3.066571, 3.04349, 3.086209, 3.07363, 3.110449, 
    3.092099, 3.128219, 3.14376, 3.158431, 3.175649, 3.03221, 3.027345, 
    3.036059, 3.04815, 3.059396, 3.074396, 3.075933, 3.078751, 3.086057, 
    3.092211, 3.079644, 3.093755, 3.041039, 3.068579, 3.025508, 3.038432, 
    3.047436, 3.043482, 3.064049, 3.068912, 3.088732, 3.078473, 3.13992, 
    3.112623, 3.188801, 3.167376, 3.025646, 3.032193, 3.05506, 3.044164, 
    3.075399, 3.083125, 3.089414, 3.097471, 3.09834, 3.103122, 3.095289, 
    3.102812, 3.074429, 3.087088, 3.052438, 3.060846, 3.056975, 3.052735, 
    3.065836, 3.079842, 3.080139, 3.084641, 3.097359, 3.075526, 3.143462, 
    3.101381, 3.039343, 3.052007, 3.053816, 3.048904, 3.08235, 3.0702, 
    3.103005, 3.094113, 3.108692, 3.101441, 3.100375, 3.091083, 3.085309, 
    3.070757, 3.058953, 3.049616, 3.051785, 3.062048, 3.0807, 3.09842, 
    3.094532, 3.107582, 3.073126, 3.087541, 3.081964, 3.09652, 3.064691, 
    3.091788, 3.057794, 3.060762, 3.069959, 3.088522, 3.092636, 3.097038, 
    3.094321, 3.081174, 3.079023, 3.069735, 3.067175, 3.060116, 3.054281, 
    3.059612, 3.065219, 3.081178, 3.095615, 3.111412, 3.115285, 3.133842, 
    3.118733, 3.143698, 3.122469, 3.159281, 3.093359, 3.121841, 3.070377, 
    3.075891, 3.085884, 3.10889, 3.096451, 3.111001, 3.078938, 3.062404, 
    3.058134, 3.050184, 3.058316, 3.057654, 3.065449, 3.062942, 3.081709, 
    3.071618, 3.100349, 3.110885, 3.140777, 3.159209, 3.178049, 3.186395, 
    3.188938, 3.190002,
  2.975095, 2.991747, 2.988503, 3.001985, 2.994498, 3.003337, 2.978463, 
    2.992411, 2.983499, 2.976589, 3.028315, 3.002587, 3.05465, 3.038612, 
    3.079055, 3.05215, 3.084508, 3.078274, 3.09707, 3.091673, 3.115842, 
    3.099563, 3.128441, 3.111946, 3.114521, 3.099028, 3.007746, 3.025101, 
    3.006721, 3.009189, 3.008081, 2.994653, 2.987909, 2.973825, 2.976377, 
    2.986722, 3.0103, 3.002275, 3.022534, 3.022075, 3.044513, 3.034522, 
    3.071753, 3.061143, 3.091898, 3.084136, 3.091534, 3.089288, 3.091563, 
    3.080186, 3.085055, 3.075062, 3.036441, 3.047744, 3.01342, 2.99274, 
    2.979074, 2.969413, 2.970777, 2.973379, 2.986783, 2.999436, 3.009112, 
    3.015602, 3.022009, 3.041326, 3.051346, 3.073904, 3.069819, 3.07674, 
    3.083364, 3.09452, 3.09268, 3.097605, 3.076556, 3.09053, 3.067495, 
    3.073779, 3.02376, 3.004438, 2.996267, 2.989126, 2.971826, 2.983763, 
    2.979053, 2.99027, 2.99742, 2.993881, 3.015779, 3.007248, 3.051941, 
    3.032904, 3.082591, 3.070657, 3.085458, 3.077896, 3.090865, 3.079191, 
    3.09944, 3.103867, 3.100841, 3.112478, 3.078545, 3.091534, 2.993783, 
    2.994359, 2.997047, 2.985249, 2.984528, 2.973755, 2.983339, 2.987429, 
    2.997834, 3.004006, 3.009884, 3.022845, 3.037355, 3.057139, 3.071429, 
    3.081045, 3.075145, 3.080353, 3.074531, 3.071806, 3.102207, 3.085101, 
    3.110802, 3.109374, 3.097723, 3.109535, 2.994765, 2.991446, 2.979955, 
    2.988944, 2.972584, 2.981732, 2.987005, 3.007428, 3.011931, 3.016115, 
    3.024391, 3.035046, 3.053267, 3.069166, 3.08375, 3.082679, 3.083056, 
    3.086323, 3.078237, 3.087653, 3.089236, 3.085098, 3.109183, 3.102283, 
    3.109344, 3.104849, 2.992524, 2.998111, 2.995091, 3.000773, 2.99677, 
    3.014611, 3.01998, 3.044941, 3.034836, 3.0509, 3.036512, 3.039057, 
    3.051427, 3.037287, 3.068289, 3.04724, 3.08645, 3.065311, 3.08778, 
    3.083687, 3.090466, 3.09655, 3.104221, 3.118425, 3.11513, 3.127044, 
    3.006458, 3.013739, 3.013096, 3.02073, 3.026389, 3.038615, 3.057803, 
    3.050573, 3.063857, 3.066531, 3.046354, 3.058728, 3.01862, 3.025185, 
    3.021273, 3.007032, 3.05224, 3.029212, 3.071666, 3.05922, 3.095682, 
    3.077497, 3.113317, 3.12876, 3.143356, 3.160506, 3.017718, 3.012763, 
    3.021639, 3.033963, 3.04515, 3.059978, 3.061498, 3.064286, 3.071516, 
    3.077608, 3.065169, 3.079138, 3.026712, 3.054225, 3.010893, 3.024056, 
    3.033235, 3.029204, 3.049748, 3.054554, 3.074164, 3.064011, 3.124943, 
    3.097839, 3.173622, 3.152262, 3.011034, 3.0177, 3.040867, 3.029899, 
    3.060969, 3.068613, 3.074839, 3.082819, 3.08368, 3.088419, 3.080658, 
    3.088111, 3.060009, 3.072536, 3.038278, 3.046583, 3.042759, 3.038572, 
    3.051514, 3.065364, 3.065659, 3.070114, 3.082706, 3.061095, 3.128462, 
    3.086691, 3.024985, 3.037853, 3.039639, 3.034733, 3.067846, 3.055828, 
    3.088303, 3.079492, 3.09394, 3.086753, 3.085697, 3.076492, 3.070775, 
    3.056379, 3.044713, 3.035459, 3.037634, 3.047771, 3.066213, 3.083759, 
    3.079908, 3.09284, 3.058722, 3.072984, 3.067465, 3.081876, 3.050382, 
    3.077188, 3.043568, 3.0465, 3.05559, 3.073955, 3.07803, 3.08239, 
    3.079698, 3.066682, 3.064554, 3.055368, 3.052838, 3.045861, 3.040099, 
    3.045364, 3.050904, 3.066687, 3.08098, 3.096638, 3.10048, 3.118901, 
    3.1039, 3.128696, 3.107607, 3.144201, 3.078745, 3.106985, 3.056004, 
    3.061456, 3.071344, 3.094136, 3.081808, 3.09623, 3.064471, 3.048122, 
    3.043904, 3.036038, 3.044083, 3.043429, 3.051132, 3.048655, 3.067212, 
    3.05723, 3.085671, 3.096115, 3.125794, 3.14413, 3.162899, 3.171222, 
    3.17376, 3.174821,
  2.975602, 2.994002, 2.990413, 3.005335, 2.997046, 3.006833, 2.979321, 
    2.994736, 2.984883, 2.977252, 3.034556, 3.006002, 3.064565, 3.046093, 
    3.092759, 3.061682, 3.099072, 3.091855, 3.113637, 3.107377, 3.135455, 
    3.116532, 3.150133, 3.130921, 3.133918, 3.115911, 3.01172, 3.030984, 
    3.010584, 3.01332, 3.012092, 2.997217, 2.989757, 2.9742, 2.977017, 
    2.988446, 3.014552, 3.005657, 3.028132, 3.027622, 3.052884, 3.041461, 
    3.084312, 3.072057, 3.107638, 3.098642, 3.107215, 3.104612, 3.107249, 
    3.094068, 3.099707, 3.088139, 3.043597, 3.056605, 3.018013, 2.9951, 
    2.979995, 2.96933, 2.970838, 2.973709, 2.988513, 3.002512, 3.013235, 
    3.020434, 3.027549, 3.049215, 3.060756, 3.086799, 3.082077, 3.09008, 
    3.097748, 3.110678, 3.108545, 3.114259, 3.089868, 3.106052, 3.079391, 
    3.086655, 3.029493, 3.008053, 2.999003, 2.991103, 2.971995, 2.985175, 
    2.979971, 2.992368, 3.00028, 2.996363, 3.020632, 3.011168, 3.061442, 
    3.03966, 3.096853, 3.083045, 3.100173, 3.091418, 3.10644, 3.092916, 
    3.116388, 3.12153, 3.118015, 3.131541, 3.092169, 3.107216, 2.996254, 
    2.996892, 2.999867, 2.986817, 2.98602, 2.974123, 2.984706, 2.989227, 
    3.000738, 3.007575, 3.01409, 3.028477, 3.044647, 3.067436, 3.083938, 
    3.095062, 3.088234, 3.094262, 3.087525, 3.084374, 3.119603, 3.09976, 
    3.129591, 3.127931, 3.114395, 3.128118, 2.997341, 2.993669, 2.980968, 
    2.990902, 2.972831, 2.982931, 2.988757, 3.011367, 3.016361, 3.021003, 
    3.030196, 3.042045, 3.06297, 3.081322, 3.098195, 3.096955, 3.097391, 
    3.101176, 3.091813, 3.102716, 3.104552, 3.099757, 3.127708, 3.11969, 
    3.127896, 3.122671, 2.994862, 3.001045, 2.997702, 3.003993, 2.99956, 
    3.019335, 3.025295, 3.053377, 3.041811, 3.060242, 3.043677, 3.046604, 
    3.060848, 3.044569, 3.080308, 3.056024, 3.101323, 3.076868, 3.102864, 
    3.098122, 3.105977, 3.113035, 3.121941, 3.138462, 3.134626, 3.148505, 
    3.010292, 3.018366, 3.017653, 3.026128, 3.032416, 3.046097, 3.068202, 
    3.059865, 3.07519, 3.078278, 3.055004, 3.069269, 3.023784, 3.031077, 
    3.026731, 3.010928, 3.061786, 3.035555, 3.084212, 3.069836, 3.112028, 
    3.090956, 3.132518, 3.150504, 3.167412, 3.186846, 3.022783, 3.017284, 
    3.027138, 3.040839, 3.053617, 3.070711, 3.072466, 3.075684, 3.084038, 
    3.091085, 3.076704, 3.092855, 3.032774, 3.064075, 3.015209, 3.029823, 
    3.040029, 3.035546, 3.058914, 3.064455, 3.0871, 3.075367, 3.146054, 
    3.11453, 3.201745, 3.177498, 3.015366, 3.022763, 3.048687, 3.036318, 
    3.071856, 3.080683, 3.087881, 3.097116, 3.098114, 3.103604, 3.094614, 
    3.103248, 3.070748, 3.085218, 3.045709, 3.055268, 3.050865, 3.046046, 
    3.06095, 3.07693, 3.077271, 3.082418, 3.096984, 3.072001, 3.150156, 
    3.101601, 3.030856, 3.045219, 3.047275, 3.041697, 3.079797, 3.065924, 
    3.10347, 3.093265, 3.110007, 3.101674, 3.10045, 3.089793, 3.083182, 
    3.066558, 3.053114, 3.042505, 3.044967, 3.056636, 3.07791, 3.098206, 
    3.093746, 3.10873, 3.069262, 3.085736, 3.079356, 3.096025, 3.059645, 
    3.090597, 3.051796, 3.055173, 3.065649, 3.086859, 3.091573, 3.09662, 
    3.093504, 3.078453, 3.075994, 3.065393, 3.062475, 3.054437, 3.047803, 
    3.053864, 3.060246, 3.078458, 3.094988, 3.113136, 3.117597, 3.139016, 
    3.121569, 3.15043, 3.125876, 3.168368, 3.0924, 3.125153, 3.066126, 
    3.072417, 3.083839, 3.110233, 3.095947, 3.112662, 3.075898, 3.057041, 
    3.052183, 3.043149, 3.05239, 3.051637, 3.060509, 3.057654, 3.079065, 
    3.067541, 3.10042, 3.112529, 3.147048, 3.168288, 3.189563, 3.199017, 
    3.201901, 3.203108,
  3.25515, 3.278626, 3.274039, 3.293146, 3.282522, 3.295069, 3.259885, 
    3.279566, 3.266977, 3.25725, 3.330328, 3.294003, 3.368102, 3.344811, 
    3.403897, 3.364459, 3.411954, 3.402744, 3.4306, 3.422575, 3.458685, 
    3.434315, 3.477687, 3.452834, 3.456701, 3.433517, 3.301347, 3.325852, 
    3.299887, 3.303405, 3.301825, 3.282741, 3.2732, 3.253366, 3.256951, 
    3.271524, 3.304989, 3.29356, 3.322283, 3.321645, 3.353359, 3.338991, 
    3.393142, 3.377584, 3.42291, 3.411404, 3.422368, 3.419036, 3.422411, 
    3.405566, 3.412764, 3.398011, 3.341673, 3.35805, 3.309445, 3.280032, 
    3.260744, 3.247179, 3.249091, 3.252741, 3.27161, 3.289525, 3.303295, 
    3.312564, 3.321554, 3.348738, 3.363289, 3.396305, 3.3903, 3.400483, 
    3.410263, 3.426805, 3.424072, 3.431397, 3.400212, 3.420879, 3.386889, 
    3.396122, 3.323986, 3.296636, 3.285028, 3.27492, 3.250562, 3.267349, 
    3.260714, 3.276538, 3.286664, 3.281648, 3.312818, 3.300638, 3.364155, 
    3.33673, 3.40912, 3.391531, 3.413361, 3.402188, 3.421375, 3.404098, 
    3.434131, 3.440738, 3.43622, 3.453634, 3.403145, 3.422369, 3.281508, 
    3.282326, 3.286136, 3.269445, 3.268428, 3.253268, 3.266751, 3.272522, 
    3.287252, 3.296021, 3.304396, 3.322716, 3.342993, 3.371733, 3.392666, 
    3.406835, 3.398133, 3.405813, 3.39723, 3.39322, 3.43826, 3.412832, 
    3.451119, 3.448978, 3.431572, 3.449219, 3.282899, 3.278201, 3.261984, 
    3.274663, 3.251625, 3.264487, 3.271923, 3.300894, 3.307318, 3.313298, 
    3.324866, 3.339723, 3.366086, 3.389341, 3.410833, 3.40925, 3.409807, 
    3.414642, 3.402691, 3.416611, 3.418959, 3.412828, 3.448692, 3.438373, 
    3.448933, 3.442206, 3.279727, 3.287645, 3.283362, 3.291425, 3.285742, 
    3.311147, 3.318736, 3.35398, 3.33943, 3.36264, 3.341774, 3.345454, 
    3.363405, 3.342894, 3.388053, 3.357317, 3.41483, 3.383685, 3.4168, 
    3.41074, 3.420783, 3.429827, 3.441267, 3.462571, 3.457615, 3.475575, 
    3.299512, 3.3099, 3.308981, 3.319778, 3.327646, 3.344816, 3.372702, 
    3.362164, 3.381556, 3.385475, 3.356032, 3.374054, 3.316848, 3.32597, 
    3.320532, 3.30033, 3.36459, 3.331579, 3.393014, 3.374772, 3.428535, 
    3.401599, 3.454893, 3.478169, 3.500344, 3.526617, 3.315592, 3.308506, 
    3.32104, 3.33821, 3.354283, 3.37588, 3.378103, 3.382183, 3.392793, 
    3.401764, 3.383477, 3.404019, 3.328095, 3.367483, 3.305835, 3.3244, 
    3.337192, 3.331568, 3.360964, 3.367963, 3.396688, 3.381781, 3.472398, 
    3.431745, 3.546502, 3.513958, 3.306037, 3.315567, 3.348075, 3.332537, 
    3.37733, 3.388529, 3.397683, 3.409456, 3.41073, 3.417746, 3.406263, 
    3.417291, 3.375926, 3.394294, 3.344328, 3.356364, 3.350816, 3.344752, 
    3.363534, 3.383764, 3.384196, 3.390733, 3.409287, 3.377513, 3.477717, 
    3.415185, 3.325692, 3.343712, 3.346297, 3.339286, 3.387403, 3.36982, 
    3.417575, 3.404543, 3.425944, 3.415278, 3.413714, 3.400118, 3.391705, 
    3.370623, 3.353649, 3.340301, 3.343396, 3.358089, 3.385008, 3.410847, 
    3.405155, 3.424309, 3.374044, 3.394952, 3.386843, 3.408063, 3.361886, 
    3.401142, 3.351989, 3.356244, 3.369473, 3.396381, 3.402385, 3.408822, 
    3.404847, 3.385696, 3.382577, 3.36915, 3.365461, 3.355317, 3.346962, 
    3.354594, 3.362645, 3.385703, 3.406739, 3.429956, 3.435683, 3.463288, 
    3.440788, 3.478072, 3.446331, 3.501632, 3.403439, 3.4454, 3.370076, 
    3.378041, 3.39254, 3.426234, 3.407963, 3.429348, 3.382455, 3.3586, 
    3.352476, 3.34111, 3.352736, 3.351788, 3.362978, 3.359374, 3.386474, 
    3.371866, 3.413676, 3.429178, 3.473686, 3.501524, 3.530303, 3.542899, 
    3.546709, 3.548304,
  3.812404, 3.852934, 3.844962, 3.878334, 3.859723, 3.881718, 3.820525, 
    3.854569, 3.832741, 3.816003, 3.945438, 3.879841, 4.016917, 3.9726, 
    4.0849, 4.009933, 4.100402, 4.082691, 4.136672, 4.120995, 4.192385, 
    4.143967, 4.230845, 4.180668, 4.188404, 4.142398, 3.892797, 3.937106, 
    3.890215, 3.896438, 3.893641, 3.860107, 3.843507, 3.809351, 3.81549, 
    3.840604, 3.899245, 3.879062, 3.93048, 3.929298, 3.988771, 3.961649, 
    4.064365, 4.034974, 4.121645, 4.09934, 4.12059, 4.114112, 4.120675, 
    4.088104, 4.101967, 4.07364, 3.96669, 3.997692, 3.907157, 3.855382, 
    3.822002, 3.79879, 3.802048, 3.808282, 3.840752, 3.871976, 3.896244, 
    3.912713, 3.929128, 3.980017, 4.007693, 4.070387, 4.058969, 4.078363, 
    4.09714, 4.129245, 4.123909, 4.138236, 4.077845, 4.117692, 4.052507, 
    4.070038, 3.93364, 3.884478, 3.864101, 3.846492, 3.804559, 3.833384, 
    3.82195, 3.849302, 3.866963, 3.8582, 3.913166, 3.891543, 4.009351, 
    3.957408, 4.094937, 4.061305, 4.103119, 4.081625, 4.118658, 4.085285, 
    4.143604, 4.156631, 4.147716, 4.182265, 4.083458, 4.120592, 3.857955, 
    3.859381, 3.866039, 3.837005, 3.835247, 3.809183, 3.83235, 3.842333, 
    3.867992, 3.883395, 3.898193, 3.931282, 3.969173, 4.023899, 4.06346, 
    4.090541, 4.073873, 4.088578, 4.07215, 4.064515, 4.151737, 4.102098, 
    4.177244, 4.172979, 4.138579, 4.173459, 3.860382, 3.852194, 3.824134, 
    3.846046, 3.806374, 3.828444, 3.841294, 3.891994, 3.903378, 3.914021, 
    3.935273, 3.963025, 4.013051, 4.057151, 4.098239, 4.095187, 4.096261, 
    4.105595, 4.082589, 4.109408, 4.113962, 4.10209, 4.172409, 4.151959, 
    4.172888, 4.159535, 3.85485, 3.868681, 3.861191, 3.875309, 3.865349, 
    3.910188, 3.923913, 3.989951, 3.962474, 4.006452, 3.966879, 3.973812, 
    4.007916, 3.968988, 4.05471, 3.996296, 4.105959, 4.046456, 4.109774, 
    4.098059, 4.117507, 4.135157, 4.157677, 4.200199, 4.190238, 4.226539, 
    3.889552, 3.907967, 3.906333, 3.92584, 3.940441, 3.972609, 4.025766, 
    4.005544, 4.042442, 4.049835, 3.99385, 4.028354, 3.920425, 3.937324, 
    3.927236, 3.890998, 4.010183, 3.947774, 4.064123, 4.029699, 4.132627, 
    4.080498, 4.184784, 4.231829, 4.277548, 4.332257, 3.918117, 3.905488, 
    3.928177, 3.960183, 3.990527, 4.031775, 4.035948, 4.043624, 4.063704, 
    4.080813, 4.046063, 4.085135, 3.941278, 4.015729, 3.900746, 3.934407, 
    3.958275, 3.947752, 4.00325, 4.01665, 4.071117, 4.042866, 4.220076, 
    4.138918, 4.374617, 4.306068, 3.901103, 3.918072, 3.978762, 3.949562, 
    4.034495, 4.055613, 4.073015, 4.095584, 4.098041, 4.111609, 4.089443, 
    4.110726, 4.031862, 4.066556, 3.971689, 3.994482, 3.98395, 3.972489, 
    4.008162, 4.046605, 4.04742, 4.059791, 4.095261, 4.034841, 4.230907, 
    4.106647, 3.936809, 3.970528, 3.975404, 3.962203, 4.053481, 4.020219, 
    4.111277, 4.086139, 4.127563, 4.106827, 4.103802, 4.077664, 4.061635, 
    4.021763, 3.989323, 3.96411, 3.969933, 3.997767, 4.048954, 4.098266, 
    4.087315, 4.124372, 4.028336, 4.06781, 4.052423, 4.092904, 4.005011, 
    4.079623, 3.986172, 3.994255, 4.019551, 4.070532, 4.082003, 4.094365, 
    4.086722, 4.050253, 4.044366, 4.01893, 4.011852, 3.992491, 3.97666, 
    3.991118, 4.006463, 4.050266, 4.090358, 4.135411, 4.146657, 4.201642, 
    4.156729, 4.231632, 4.167714, 4.280232, 4.084022, 4.165865, 4.020711, 
    4.035831, 4.063221, 4.12813, 4.09271, 4.13422, 4.044136, 3.99874, 
    3.987096, 3.965631, 3.98759, 3.985791, 4.007098, 4.000216, 4.051723, 
    4.024156, 4.103727, 4.133886, 4.222693, 4.280006, 4.339907, 4.366785, 
    4.375067, 4.378545,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24855.36, 24876.16, 24872.09, 24889.11, 24879.63, 24890.83, 24859.54, 
    24877, 24865.82, 24857.22, 24922.92, 24889.88, 24958.25, 24936.42, 
    24991.74, 24954.83, 24999.33, 24990.66, 25016.99, 25009.37, 25043.91, 
    25020.53, 25062.3, 25038.28, 25042, 25019.77, 24896.45, 24918.76, 
    24895.14, 24898.3, 24896.88, 24879.83, 24871.34, 24853.79, 24856.95, 
    24869.85, 24899.72, 24889.48, 24915.45, 24914.86, 24944.41, 24930.99, 
    24981.65, 24967.14, 25009.69, 24998.81, 25009.18, 25006.02, 25009.22, 
    24993.31, 25000.09, 24986.22, 24933.49, 24948.8, 24903.72, 24877.41, 
    24860.3, 24848.33, 24850.02, 24853.24, 24869.93, 24885.88, 24898.2, 
    24906.53, 24914.77, 24940.08, 24953.72, 24984.62, 24979, 24988.54, 
    24997.73, 25013.38, 25010.79, 25017.75, 24988.28, 25007.76, 24975.81, 
    24984.45, 24917.03, 24892.23, 24881.87, 24872.87, 24851.32, 24866.15, 
    24860.28, 24874.31, 24883.32, 24878.85, 24906.76, 24895.82, 24954.54, 
    24928.88, 24996.66, 24980.15, 25000.66, 24990.14, 25008.23, 24991.93, 
    25020.35, 25026.7, 25022.34, 25039.05, 24991.04, 25009.18, 24878.73, 
    24879.46, 24882.85, 24868.01, 24867.11, 24853.7, 24865.62, 24870.74, 
    24883.85, 24891.68, 24899.19, 24915.85, 24934.72, 24961.68, 24981.21, 
    24994.51, 24986.33, 24993.54, 24985.48, 24981.73, 25024.33, 25000.16, 
    25036.64, 25034.58, 25017.91, 25034.81, 24879.97, 24875.79, 24861.4, 
    24872.64, 24852.25, 24863.62, 24870.21, 24896.05, 24901.81, 24907.19, 
    24917.84, 24931.67, 24956.36, 24978.1, 24998.27, 24996.78, 24997.3, 
    25001.87, 24990.61, 25003.73, 25005.95, 25000.15, 25034.31, 25024.44, 
    25034.54, 25028.1, 24877.14, 24884.2, 24880.38, 24887.57, 24882.5, 
    24905.25, 24912.16, 24944.99, 24931.4, 24953.12, 24933.58, 24937.02, 
    24953.83, 24934.63, 24976.9, 24948.12, 25002.04, 24972.82, 25003.9, 
    24998.18, 25007.67, 25016.25, 25027.2, 25047.66, 25042.88, 25060.25, 
    24894.81, 24904.13, 24903.31, 24913.13, 24920.42, 24936.42, 24962.59, 
    24952.67, 24970.84, 24974.49, 24946.91, 24963.86, 24910.41, 24918.87, 
    24913.82, 24895.54, 24954.95, 24924.08, 24981.54, 24964.53, 25015.03, 
    24989.58, 25040.26, 25062.77, 25084.43, 25110.18, 24909.26, 24902.88, 
    24914.29, 24930.26, 24945.27, 24965.56, 24967.62, 24971.42, 24981.33, 
    24989.74, 24972.63, 24991.86, 24920.84, 24957.67, 24900.48, 24917.41, 
    24929.31, 24924.07, 24951.54, 24958.12, 24984.98, 24971.05, 25057.16, 
    25018.08, 25130, 25097.82, 24900.66, 24909.23, 24939.46, 24924.97, 
    24966.91, 24977.34, 24985.91, 24996.97, 24998.18, 25004.8, 24993.97, 
    25004.37, 24965.6, 24982.73, 24935.96, 24947.22, 24942.03, 24936.36, 
    24953.96, 24972.9, 24973.3, 24979.4, 24996.82, 24967.08, 25062.33, 
    25002.38, 24918.61, 24935.39, 24937.8, 24931.26, 24976.29, 24959.87, 
    25004.64, 24992.35, 25012.57, 25002.47, 25000.99, 24988.19, 24980.31, 
    24960.63, 24944.68, 24932.21, 24935.1, 24948.84, 24974.06, 24998.29, 
    24992.93, 25011.01, 24963.85, 24983.35, 24975.77, 24995.66, 24952.41, 
    24989.15, 24943.12, 24947.11, 24959.55, 24984.69, 24990.32, 24996.38, 
    24992.63, 24974.7, 24971.79, 24959.24, 24955.77, 24946.24, 24938.42, 
    24945.56, 24953.12, 24974.71, 24994.42, 25016.38, 25021.83, 25048.35, 
    25026.74, 25062.67, 25032.04, 25085.69, 24991.31, 25031.15, 24960.12, 
    24967.57, 24981.09, 25012.84, 24995.57, 25015.8, 24971.68, 24949.32, 
    24943.58, 24932.96, 24943.82, 24942.94, 24953.43, 24950.05, 24975.42, 
    24961.8, 25000.95, 25015.64, 25058.41, 25085.59, 25113.78, 25126.36, 
    25130.21, 25131.83 ;

 HCSOI =
  24855.36, 24876.16, 24872.09, 24889.11, 24879.63, 24890.83, 24859.54, 
    24877, 24865.82, 24857.22, 24922.92, 24889.88, 24958.25, 24936.42, 
    24991.74, 24954.83, 24999.33, 24990.66, 25016.99, 25009.37, 25043.91, 
    25020.53, 25062.3, 25038.28, 25042, 25019.77, 24896.45, 24918.76, 
    24895.14, 24898.3, 24896.88, 24879.83, 24871.34, 24853.79, 24856.95, 
    24869.85, 24899.72, 24889.48, 24915.45, 24914.86, 24944.41, 24930.99, 
    24981.65, 24967.14, 25009.69, 24998.81, 25009.18, 25006.02, 25009.22, 
    24993.31, 25000.09, 24986.22, 24933.49, 24948.8, 24903.72, 24877.41, 
    24860.3, 24848.33, 24850.02, 24853.24, 24869.93, 24885.88, 24898.2, 
    24906.53, 24914.77, 24940.08, 24953.72, 24984.62, 24979, 24988.54, 
    24997.73, 25013.38, 25010.79, 25017.75, 24988.28, 25007.76, 24975.81, 
    24984.45, 24917.03, 24892.23, 24881.87, 24872.87, 24851.32, 24866.15, 
    24860.28, 24874.31, 24883.32, 24878.85, 24906.76, 24895.82, 24954.54, 
    24928.88, 24996.66, 24980.15, 25000.66, 24990.14, 25008.23, 24991.93, 
    25020.35, 25026.7, 25022.34, 25039.05, 24991.04, 25009.18, 24878.73, 
    24879.46, 24882.85, 24868.01, 24867.11, 24853.7, 24865.62, 24870.74, 
    24883.85, 24891.68, 24899.19, 24915.85, 24934.72, 24961.68, 24981.21, 
    24994.51, 24986.33, 24993.54, 24985.48, 24981.73, 25024.33, 25000.16, 
    25036.64, 25034.58, 25017.91, 25034.81, 24879.97, 24875.79, 24861.4, 
    24872.64, 24852.25, 24863.62, 24870.21, 24896.05, 24901.81, 24907.19, 
    24917.84, 24931.67, 24956.36, 24978.1, 24998.27, 24996.78, 24997.3, 
    25001.87, 24990.61, 25003.73, 25005.95, 25000.15, 25034.31, 25024.44, 
    25034.54, 25028.1, 24877.14, 24884.2, 24880.38, 24887.57, 24882.5, 
    24905.25, 24912.16, 24944.99, 24931.4, 24953.12, 24933.58, 24937.02, 
    24953.83, 24934.63, 24976.9, 24948.12, 25002.04, 24972.82, 25003.9, 
    24998.18, 25007.67, 25016.25, 25027.2, 25047.66, 25042.88, 25060.25, 
    24894.81, 24904.13, 24903.31, 24913.13, 24920.42, 24936.42, 24962.59, 
    24952.67, 24970.84, 24974.49, 24946.91, 24963.86, 24910.41, 24918.87, 
    24913.82, 24895.54, 24954.95, 24924.08, 24981.54, 24964.53, 25015.03, 
    24989.58, 25040.26, 25062.77, 25084.43, 25110.18, 24909.26, 24902.88, 
    24914.29, 24930.26, 24945.27, 24965.56, 24967.62, 24971.42, 24981.33, 
    24989.74, 24972.63, 24991.86, 24920.84, 24957.67, 24900.48, 24917.41, 
    24929.31, 24924.07, 24951.54, 24958.12, 24984.98, 24971.05, 25057.16, 
    25018.08, 25130, 25097.82, 24900.66, 24909.23, 24939.46, 24924.97, 
    24966.91, 24977.34, 24985.91, 24996.97, 24998.18, 25004.8, 24993.97, 
    25004.37, 24965.6, 24982.73, 24935.96, 24947.22, 24942.03, 24936.36, 
    24953.96, 24972.9, 24973.3, 24979.4, 24996.82, 24967.08, 25062.33, 
    25002.38, 24918.61, 24935.39, 24937.8, 24931.26, 24976.29, 24959.87, 
    25004.64, 24992.35, 25012.57, 25002.47, 25000.99, 24988.19, 24980.31, 
    24960.63, 24944.68, 24932.21, 24935.1, 24948.84, 24974.06, 24998.29, 
    24992.93, 25011.01, 24963.85, 24983.35, 24975.77, 24995.66, 24952.41, 
    24989.15, 24943.12, 24947.11, 24959.55, 24984.69, 24990.32, 24996.38, 
    24992.63, 24974.7, 24971.79, 24959.24, 24955.77, 24946.24, 24938.42, 
    24945.56, 24953.12, 24974.71, 24994.42, 25016.38, 25021.83, 25048.35, 
    25026.74, 25062.67, 25032.04, 25085.69, 24991.31, 25031.15, 24960.12, 
    24967.57, 24981.09, 25012.84, 24995.57, 25015.8, 24971.68, 24949.32, 
    24943.58, 24932.96, 24943.82, 24942.94, 24953.43, 24950.05, 24975.42, 
    24961.8, 25000.95, 25015.64, 25058.41, 25085.59, 25113.78, 25126.36, 
    25130.21, 25131.83 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.215762e-08, 6.243169e-08, 6.237841e-08, 6.259947e-08, 6.247685e-08, 
    6.26216e-08, 6.221319e-08, 6.244257e-08, 6.229614e-08, 6.21823e-08, 
    6.302847e-08, 6.260934e-08, 6.346394e-08, 6.319659e-08, 6.386823e-08, 
    6.342233e-08, 6.395815e-08, 6.385538e-08, 6.416472e-08, 6.40761e-08, 
    6.447177e-08, 6.420563e-08, 6.46769e-08, 6.440823e-08, 6.445025e-08, 
    6.419685e-08, 6.269369e-08, 6.297628e-08, 6.267695e-08, 6.271725e-08, 
    6.269916e-08, 6.247938e-08, 6.236861e-08, 6.213668e-08, 6.217878e-08, 
    6.234914e-08, 6.273537e-08, 6.260426e-08, 6.29347e-08, 6.292724e-08, 
    6.329513e-08, 6.312926e-08, 6.374764e-08, 6.357188e-08, 6.40798e-08, 
    6.395206e-08, 6.40738e-08, 6.403688e-08, 6.407428e-08, 6.388693e-08, 
    6.39672e-08, 6.380235e-08, 6.316031e-08, 6.334899e-08, 6.278628e-08, 
    6.244793e-08, 6.222324e-08, 6.20638e-08, 6.208634e-08, 6.212931e-08, 
    6.235014e-08, 6.255778e-08, 6.271602e-08, 6.282187e-08, 6.292617e-08, 
    6.324185e-08, 6.340898e-08, 6.378317e-08, 6.371565e-08, 6.383004e-08, 
    6.393935e-08, 6.412285e-08, 6.409265e-08, 6.417349e-08, 6.382704e-08, 
    6.405729e-08, 6.367719e-08, 6.378114e-08, 6.295448e-08, 6.263964e-08, 
    6.250578e-08, 6.238865e-08, 6.210367e-08, 6.230047e-08, 6.222289e-08, 
    6.240747e-08, 6.252476e-08, 6.246675e-08, 6.282476e-08, 6.268557e-08, 
    6.341888e-08, 6.310301e-08, 6.39266e-08, 6.372951e-08, 6.397384e-08, 
    6.384917e-08, 6.406279e-08, 6.387053e-08, 6.420358e-08, 6.427612e-08, 
    6.422655e-08, 6.441695e-08, 6.385987e-08, 6.40738e-08, 6.246512e-08, 
    6.247458e-08, 6.251866e-08, 6.232491e-08, 6.231306e-08, 6.213552e-08, 
    6.229349e-08, 6.236077e-08, 6.253156e-08, 6.263257e-08, 6.27286e-08, 
    6.293975e-08, 6.317556e-08, 6.350534e-08, 6.374228e-08, 6.390112e-08, 
    6.380372e-08, 6.388971e-08, 6.379359e-08, 6.374854e-08, 6.424895e-08, 
    6.396795e-08, 6.438957e-08, 6.436624e-08, 6.417542e-08, 6.436887e-08, 
    6.248122e-08, 6.242679e-08, 6.223777e-08, 6.238569e-08, 6.211619e-08, 
    6.226703e-08, 6.235377e-08, 6.268847e-08, 6.276202e-08, 6.283021e-08, 
    6.296489e-08, 6.313774e-08, 6.344097e-08, 6.370482e-08, 6.394571e-08, 
    6.392806e-08, 6.393427e-08, 6.398808e-08, 6.385479e-08, 6.400997e-08, 
    6.403601e-08, 6.396792e-08, 6.436311e-08, 6.425022e-08, 6.436574e-08, 
    6.429224e-08, 6.244449e-08, 6.253608e-08, 6.248658e-08, 6.257967e-08, 
    6.251409e-08, 6.280568e-08, 6.289311e-08, 6.330224e-08, 6.313434e-08, 
    6.340156e-08, 6.316149e-08, 6.320403e-08, 6.341026e-08, 6.317446e-08, 
    6.369027e-08, 6.334054e-08, 6.399017e-08, 6.36409e-08, 6.401206e-08, 
    6.394467e-08, 6.405626e-08, 6.415619e-08, 6.428195e-08, 6.451393e-08, 
    6.446022e-08, 6.465423e-08, 6.267265e-08, 6.279146e-08, 6.278102e-08, 
    6.290536e-08, 6.299733e-08, 6.319667e-08, 6.35164e-08, 6.339616e-08, 
    6.361689e-08, 6.366121e-08, 6.332587e-08, 6.353175e-08, 6.2871e-08, 
    6.297773e-08, 6.291419e-08, 6.268202e-08, 6.342385e-08, 6.304312e-08, 
    6.37462e-08, 6.353994e-08, 6.414194e-08, 6.384253e-08, 6.443064e-08, 
    6.468203e-08, 6.491868e-08, 6.51952e-08, 6.285632e-08, 6.277559e-08, 
    6.292016e-08, 6.312016e-08, 6.330577e-08, 6.355251e-08, 6.357777e-08, 
    6.362399e-08, 6.374373e-08, 6.384442e-08, 6.363859e-08, 6.386966e-08, 
    6.300247e-08, 6.345691e-08, 6.274506e-08, 6.295939e-08, 6.310837e-08, 
    6.304303e-08, 6.338242e-08, 6.346242e-08, 6.378748e-08, 6.361945e-08, 
    6.461998e-08, 6.417729e-08, 6.540579e-08, 6.506244e-08, 6.274738e-08, 
    6.285605e-08, 6.323427e-08, 6.305431e-08, 6.356899e-08, 6.369568e-08, 
    6.379868e-08, 6.393034e-08, 6.394456e-08, 6.402257e-08, 6.389474e-08, 
    6.401752e-08, 6.355304e-08, 6.37606e-08, 6.319105e-08, 6.332966e-08, 
    6.326589e-08, 6.319594e-08, 6.341183e-08, 6.364183e-08, 6.364677e-08, 
    6.372051e-08, 6.392831e-08, 6.357108e-08, 6.467708e-08, 6.399399e-08, 
    6.297455e-08, 6.318386e-08, 6.321378e-08, 6.313269e-08, 6.368298e-08, 
    6.348358e-08, 6.402067e-08, 6.387551e-08, 6.411335e-08, 6.399516e-08, 
    6.397777e-08, 6.382598e-08, 6.373148e-08, 6.349272e-08, 6.329847e-08, 
    6.314445e-08, 6.318027e-08, 6.334945e-08, 6.365591e-08, 6.394584e-08, 
    6.388233e-08, 6.409527e-08, 6.353167e-08, 6.376798e-08, 6.367664e-08, 
    6.391483e-08, 6.339297e-08, 6.383731e-08, 6.327939e-08, 6.332831e-08, 
    6.347963e-08, 6.378401e-08, 6.385137e-08, 6.392327e-08, 6.387891e-08, 
    6.366369e-08, 6.362843e-08, 6.347595e-08, 6.343384e-08, 6.331766e-08, 
    6.322146e-08, 6.330935e-08, 6.340164e-08, 6.366378e-08, 6.390003e-08, 
    6.415761e-08, 6.422066e-08, 6.452161e-08, 6.427662e-08, 6.468089e-08, 
    6.433715e-08, 6.493221e-08, 6.386308e-08, 6.432707e-08, 6.348652e-08, 
    6.357706e-08, 6.374083e-08, 6.41165e-08, 6.39137e-08, 6.415087e-08, 
    6.362706e-08, 6.335529e-08, 6.328499e-08, 6.315381e-08, 6.328799e-08, 
    6.327708e-08, 6.340547e-08, 6.336422e-08, 6.367249e-08, 6.35069e-08, 
    6.397733e-08, 6.414901e-08, 6.463389e-08, 6.493114e-08, 6.523376e-08, 
    6.536735e-08, 6.540802e-08, 6.542501e-08 ;

 HR_vr =
  2.70791e-07, 2.715254e-07, 2.713828e-07, 2.719745e-07, 2.716464e-07, 
    2.720337e-07, 2.709401e-07, 2.715544e-07, 2.711623e-07, 2.708573e-07, 
    2.731212e-07, 2.720009e-07, 2.74284e-07, 2.735708e-07, 2.753612e-07, 
    2.741729e-07, 2.756007e-07, 2.753273e-07, 2.761504e-07, 2.759147e-07, 
    2.76966e-07, 2.762592e-07, 2.775106e-07, 2.767974e-07, 2.769089e-07, 
    2.762358e-07, 2.722268e-07, 2.729817e-07, 2.721819e-07, 2.722897e-07, 
    2.722414e-07, 2.716531e-07, 2.713563e-07, 2.70735e-07, 2.708479e-07, 
    2.713043e-07, 2.723381e-07, 2.719875e-07, 2.728713e-07, 2.728514e-07, 
    2.738338e-07, 2.73391e-07, 2.750403e-07, 2.74572e-07, 2.759245e-07, 
    2.755846e-07, 2.759085e-07, 2.758104e-07, 2.759098e-07, 2.754112e-07, 
    2.756249e-07, 2.751861e-07, 2.734739e-07, 2.739775e-07, 2.724744e-07, 
    2.715686e-07, 2.70967e-07, 2.705395e-07, 2.706e-07, 2.707151e-07, 
    2.713069e-07, 2.718631e-07, 2.722866e-07, 2.725697e-07, 2.728485e-07, 
    2.736912e-07, 2.741373e-07, 2.751348e-07, 2.749551e-07, 2.752597e-07, 
    2.755508e-07, 2.76039e-07, 2.759587e-07, 2.761736e-07, 2.752518e-07, 
    2.758645e-07, 2.748527e-07, 2.751296e-07, 2.729234e-07, 2.720822e-07, 
    2.717235e-07, 2.714101e-07, 2.706464e-07, 2.711739e-07, 2.70966e-07, 
    2.714607e-07, 2.717747e-07, 2.716194e-07, 2.725774e-07, 2.722051e-07, 
    2.741638e-07, 2.733208e-07, 2.755169e-07, 2.749921e-07, 2.756426e-07, 
    2.753108e-07, 2.758792e-07, 2.753677e-07, 2.762537e-07, 2.764465e-07, 
    2.763147e-07, 2.768207e-07, 2.753393e-07, 2.759085e-07, 2.71615e-07, 
    2.716403e-07, 2.717584e-07, 2.712393e-07, 2.712076e-07, 2.707318e-07, 
    2.711553e-07, 2.713354e-07, 2.717929e-07, 2.720632e-07, 2.723202e-07, 
    2.728847e-07, 2.735145e-07, 2.743945e-07, 2.750261e-07, 2.754491e-07, 
    2.751898e-07, 2.754187e-07, 2.751628e-07, 2.750428e-07, 2.763743e-07, 
    2.756268e-07, 2.76748e-07, 2.766861e-07, 2.761787e-07, 2.76693e-07, 
    2.716581e-07, 2.715124e-07, 2.710059e-07, 2.714023e-07, 2.7068e-07, 
    2.710843e-07, 2.713166e-07, 2.722127e-07, 2.724096e-07, 2.725919e-07, 
    2.72952e-07, 2.734137e-07, 2.742228e-07, 2.749262e-07, 2.755678e-07, 
    2.755208e-07, 2.755373e-07, 2.756805e-07, 2.753257e-07, 2.757387e-07, 
    2.758079e-07, 2.756268e-07, 2.766778e-07, 2.763778e-07, 2.766847e-07, 
    2.764895e-07, 2.715598e-07, 2.71805e-07, 2.716725e-07, 2.719216e-07, 
    2.717461e-07, 2.725261e-07, 2.727598e-07, 2.738526e-07, 2.734045e-07, 
    2.741177e-07, 2.734771e-07, 2.735906e-07, 2.741406e-07, 2.735118e-07, 
    2.748873e-07, 2.739547e-07, 2.756861e-07, 2.747556e-07, 2.757443e-07, 
    2.75565e-07, 2.758619e-07, 2.761276e-07, 2.764621e-07, 2.770781e-07, 
    2.769356e-07, 2.774505e-07, 2.721705e-07, 2.724882e-07, 2.724604e-07, 
    2.727928e-07, 2.730386e-07, 2.735711e-07, 2.74424e-07, 2.741035e-07, 
    2.74692e-07, 2.748101e-07, 2.739159e-07, 2.744649e-07, 2.727009e-07, 
    2.72986e-07, 2.728164e-07, 2.721955e-07, 2.741771e-07, 2.731608e-07, 
    2.750365e-07, 2.744868e-07, 2.760897e-07, 2.752929e-07, 2.76857e-07, 
    2.77524e-07, 2.781518e-07, 2.788838e-07, 2.726617e-07, 2.724459e-07, 
    2.728324e-07, 2.733665e-07, 2.738622e-07, 2.745203e-07, 2.745877e-07, 
    2.747109e-07, 2.7503e-07, 2.752981e-07, 2.747497e-07, 2.753653e-07, 
    2.730518e-07, 2.742653e-07, 2.723641e-07, 2.72937e-07, 2.733351e-07, 
    2.731607e-07, 2.740668e-07, 2.742802e-07, 2.751464e-07, 2.746988e-07, 
    2.773593e-07, 2.761835e-07, 2.794411e-07, 2.785324e-07, 2.723704e-07, 
    2.726611e-07, 2.736713e-07, 2.731908e-07, 2.745643e-07, 2.749019e-07, 
    2.751763e-07, 2.755268e-07, 2.755647e-07, 2.757722e-07, 2.754321e-07, 
    2.757589e-07, 2.745217e-07, 2.750749e-07, 2.735561e-07, 2.73926e-07, 
    2.737559e-07, 2.735692e-07, 2.741453e-07, 2.747583e-07, 2.747716e-07, 
    2.74968e-07, 2.755206e-07, 2.745699e-07, 2.775104e-07, 2.756955e-07, 
    2.729778e-07, 2.735366e-07, 2.736167e-07, 2.734002e-07, 2.748681e-07, 
    2.743365e-07, 2.757672e-07, 2.753809e-07, 2.760138e-07, 2.756993e-07, 
    2.756531e-07, 2.75249e-07, 2.749973e-07, 2.743609e-07, 2.738427e-07, 
    2.734317e-07, 2.735273e-07, 2.739787e-07, 2.747958e-07, 2.75568e-07, 
    2.753989e-07, 2.759657e-07, 2.744648e-07, 2.750944e-07, 2.748511e-07, 
    2.754855e-07, 2.740949e-07, 2.752785e-07, 2.737919e-07, 2.739224e-07, 
    2.74326e-07, 2.75137e-07, 2.753166e-07, 2.755079e-07, 2.7539e-07, 
    2.748166e-07, 2.747227e-07, 2.743162e-07, 2.742039e-07, 2.73894e-07, 
    2.736373e-07, 2.738718e-07, 2.74118e-07, 2.748169e-07, 2.754461e-07, 
    2.761314e-07, 2.762991e-07, 2.770981e-07, 2.764475e-07, 2.775204e-07, 
    2.766078e-07, 2.78187e-07, 2.753474e-07, 2.765815e-07, 2.743444e-07, 
    2.745859e-07, 2.75022e-07, 2.760218e-07, 2.754825e-07, 2.761133e-07, 
    2.74719e-07, 2.739942e-07, 2.738068e-07, 2.734566e-07, 2.738148e-07, 
    2.737857e-07, 2.741283e-07, 2.740183e-07, 2.748401e-07, 2.743988e-07, 
    2.756518e-07, 2.761084e-07, 2.773965e-07, 2.781846e-07, 2.789861e-07, 
    2.793395e-07, 2.794471e-07, 2.79492e-07,
  2.348912e-07, 2.357843e-07, 2.356108e-07, 2.363306e-07, 2.359315e-07, 
    2.364027e-07, 2.350724e-07, 2.358197e-07, 2.353428e-07, 2.349718e-07, 
    2.377259e-07, 2.363628e-07, 2.391405e-07, 2.382725e-07, 2.404518e-07, 
    2.390054e-07, 2.407432e-07, 2.404103e-07, 2.414124e-07, 2.411254e-07, 
    2.424057e-07, 2.415448e-07, 2.430689e-07, 2.422003e-07, 2.423362e-07, 
    2.415164e-07, 2.366374e-07, 2.375562e-07, 2.365829e-07, 2.36714e-07, 
    2.366552e-07, 2.359396e-07, 2.355787e-07, 2.34823e-07, 2.349603e-07, 
    2.355154e-07, 2.367729e-07, 2.363463e-07, 2.374214e-07, 2.373972e-07, 
    2.385926e-07, 2.380538e-07, 2.40061e-07, 2.39491e-07, 2.411374e-07, 
    2.407236e-07, 2.41118e-07, 2.409984e-07, 2.411195e-07, 2.405125e-07, 
    2.407726e-07, 2.402384e-07, 2.381547e-07, 2.387675e-07, 2.369386e-07, 
    2.35837e-07, 2.351052e-07, 2.345854e-07, 2.346589e-07, 2.347989e-07, 
    2.355186e-07, 2.36195e-07, 2.367101e-07, 2.370545e-07, 2.373937e-07, 
    2.384193e-07, 2.389621e-07, 2.401761e-07, 2.399573e-07, 2.403281e-07, 
    2.406824e-07, 2.412768e-07, 2.41179e-07, 2.414407e-07, 2.403185e-07, 
    2.410644e-07, 2.398326e-07, 2.401697e-07, 2.374853e-07, 2.364615e-07, 
    2.360255e-07, 2.356442e-07, 2.347154e-07, 2.353568e-07, 2.35104e-07, 
    2.357055e-07, 2.360875e-07, 2.358986e-07, 2.370639e-07, 2.36611e-07, 
    2.389943e-07, 2.379684e-07, 2.406411e-07, 2.400022e-07, 2.407942e-07, 
    2.403902e-07, 2.410823e-07, 2.404594e-07, 2.415382e-07, 2.41773e-07, 
    2.416125e-07, 2.422287e-07, 2.404249e-07, 2.411179e-07, 2.358933e-07, 
    2.359241e-07, 2.360676e-07, 2.354364e-07, 2.353978e-07, 2.348193e-07, 
    2.353342e-07, 2.355533e-07, 2.361096e-07, 2.364385e-07, 2.36751e-07, 
    2.374378e-07, 2.382042e-07, 2.39275e-07, 2.400437e-07, 2.405586e-07, 
    2.402429e-07, 2.405216e-07, 2.4021e-07, 2.40064e-07, 2.41685e-07, 
    2.40775e-07, 2.421401e-07, 2.420646e-07, 2.414469e-07, 2.420731e-07, 
    2.359457e-07, 2.357684e-07, 2.351525e-07, 2.356346e-07, 2.347562e-07, 
    2.352479e-07, 2.355305e-07, 2.366203e-07, 2.368597e-07, 2.370815e-07, 
    2.375196e-07, 2.380814e-07, 2.390661e-07, 2.399221e-07, 2.407031e-07, 
    2.406459e-07, 2.40666e-07, 2.408403e-07, 2.404084e-07, 2.409112e-07, 
    2.409955e-07, 2.40775e-07, 2.420545e-07, 2.416892e-07, 2.42063e-07, 
    2.418252e-07, 2.358261e-07, 2.361244e-07, 2.359632e-07, 2.362662e-07, 
    2.360527e-07, 2.370016e-07, 2.37286e-07, 2.386156e-07, 2.380703e-07, 
    2.389382e-07, 2.381585e-07, 2.382967e-07, 2.389662e-07, 2.382007e-07, 
    2.398749e-07, 2.387399e-07, 2.408471e-07, 2.397146e-07, 2.40918e-07, 
    2.406997e-07, 2.410612e-07, 2.413847e-07, 2.417919e-07, 2.425422e-07, 
    2.423685e-07, 2.429958e-07, 2.365689e-07, 2.369555e-07, 2.369216e-07, 
    2.37326e-07, 2.37625e-07, 2.382728e-07, 2.393109e-07, 2.389207e-07, 
    2.39637e-07, 2.397807e-07, 2.386925e-07, 2.393607e-07, 2.372142e-07, 
    2.375612e-07, 2.373547e-07, 2.365994e-07, 2.390105e-07, 2.377737e-07, 
    2.400564e-07, 2.393873e-07, 2.413386e-07, 2.403686e-07, 2.422729e-07, 
    2.430854e-07, 2.4385e-07, 2.44742e-07, 2.371665e-07, 2.369039e-07, 
    2.373741e-07, 2.380241e-07, 2.386271e-07, 2.394281e-07, 2.395101e-07, 
    2.3966e-07, 2.400484e-07, 2.403748e-07, 2.397073e-07, 2.404566e-07, 
    2.376414e-07, 2.391178e-07, 2.368045e-07, 2.375015e-07, 2.379859e-07, 
    2.377735e-07, 2.388761e-07, 2.391358e-07, 2.401901e-07, 2.396453e-07, 
    2.428848e-07, 2.414529e-07, 2.45421e-07, 2.443138e-07, 2.368121e-07, 
    2.371656e-07, 2.383949e-07, 2.378102e-07, 2.394816e-07, 2.398925e-07, 
    2.402265e-07, 2.406532e-07, 2.406993e-07, 2.40952e-07, 2.405379e-07, 
    2.409357e-07, 2.394298e-07, 2.40103e-07, 2.382546e-07, 2.387048e-07, 
    2.384977e-07, 2.382705e-07, 2.389716e-07, 2.397178e-07, 2.397339e-07, 
    2.39973e-07, 2.406462e-07, 2.394884e-07, 2.430691e-07, 2.40859e-07, 
    2.37551e-07, 2.382311e-07, 2.383284e-07, 2.38065e-07, 2.398513e-07, 
    2.392044e-07, 2.409459e-07, 2.404756e-07, 2.412461e-07, 2.408632e-07, 
    2.408069e-07, 2.40315e-07, 2.400086e-07, 2.392341e-07, 2.386035e-07, 
    2.381032e-07, 2.382196e-07, 2.38769e-07, 2.397635e-07, 2.407034e-07, 
    2.404976e-07, 2.411875e-07, 2.393605e-07, 2.40127e-07, 2.398307e-07, 
    2.40603e-07, 2.389103e-07, 2.403513e-07, 2.385416e-07, 2.387004e-07, 
    2.391916e-07, 2.401788e-07, 2.403973e-07, 2.406303e-07, 2.404866e-07, 
    2.397887e-07, 2.396744e-07, 2.391797e-07, 2.39043e-07, 2.386658e-07, 
    2.383534e-07, 2.386388e-07, 2.389384e-07, 2.397891e-07, 2.40555e-07, 
    2.413893e-07, 2.415935e-07, 2.425668e-07, 2.417744e-07, 2.430814e-07, 
    2.419699e-07, 2.438933e-07, 2.40435e-07, 2.419376e-07, 2.39214e-07, 
    2.395078e-07, 2.400388e-07, 2.412561e-07, 2.405993e-07, 2.413674e-07, 
    2.3967e-07, 2.387879e-07, 2.385597e-07, 2.381336e-07, 2.385695e-07, 
    2.38534e-07, 2.389509e-07, 2.38817e-07, 2.398173e-07, 2.392801e-07, 
    2.408054e-07, 2.413614e-07, 2.4293e-07, 2.4389e-07, 2.448666e-07, 
    2.452972e-07, 2.454283e-07, 2.454831e-07,
  2.200482e-07, 2.210231e-07, 2.208336e-07, 2.216195e-07, 2.211837e-07, 
    2.216982e-07, 2.202459e-07, 2.210617e-07, 2.20541e-07, 2.201361e-07, 
    2.231434e-07, 2.216546e-07, 2.24689e-07, 2.237405e-07, 2.261223e-07, 
    2.245414e-07, 2.264409e-07, 2.260769e-07, 2.271727e-07, 2.268588e-07, 
    2.282594e-07, 2.273175e-07, 2.28985e-07, 2.280346e-07, 2.281832e-07, 
    2.272864e-07, 2.219544e-07, 2.229581e-07, 2.218949e-07, 2.220381e-07, 
    2.219739e-07, 2.211926e-07, 2.207987e-07, 2.199737e-07, 2.201236e-07, 
    2.207295e-07, 2.221025e-07, 2.216366e-07, 2.228107e-07, 2.227842e-07, 
    2.240902e-07, 2.235014e-07, 2.25695e-07, 2.250719e-07, 2.268719e-07, 
    2.264194e-07, 2.268507e-07, 2.267199e-07, 2.268524e-07, 2.261887e-07, 
    2.26473e-07, 2.258889e-07, 2.236117e-07, 2.242813e-07, 2.222834e-07, 
    2.210807e-07, 2.202817e-07, 2.197144e-07, 2.197946e-07, 2.199475e-07, 
    2.20733e-07, 2.214714e-07, 2.220338e-07, 2.224099e-07, 2.227804e-07, 
    2.23901e-07, 2.24494e-07, 2.258209e-07, 2.255816e-07, 2.259871e-07, 
    2.263744e-07, 2.270244e-07, 2.269174e-07, 2.272037e-07, 2.259764e-07, 
    2.267921e-07, 2.254453e-07, 2.258138e-07, 2.228807e-07, 2.217623e-07, 
    2.212864e-07, 2.2087e-07, 2.198563e-07, 2.205564e-07, 2.202804e-07, 
    2.20937e-07, 2.21354e-07, 2.211478e-07, 2.224201e-07, 2.219256e-07, 
    2.245292e-07, 2.234082e-07, 2.263292e-07, 2.256308e-07, 2.264966e-07, 
    2.260549e-07, 2.268117e-07, 2.261306e-07, 2.273102e-07, 2.27567e-07, 
    2.273915e-07, 2.280655e-07, 2.260928e-07, 2.268506e-07, 2.21142e-07, 
    2.211756e-07, 2.213323e-07, 2.206433e-07, 2.206012e-07, 2.199696e-07, 
    2.205316e-07, 2.207709e-07, 2.213782e-07, 2.217372e-07, 2.220785e-07, 
    2.228285e-07, 2.236658e-07, 2.248359e-07, 2.256761e-07, 2.26239e-07, 
    2.258938e-07, 2.261985e-07, 2.258579e-07, 2.256982e-07, 2.274708e-07, 
    2.264757e-07, 2.279686e-07, 2.27886e-07, 2.272105e-07, 2.278953e-07, 
    2.211992e-07, 2.210057e-07, 2.203334e-07, 2.208595e-07, 2.199008e-07, 
    2.204375e-07, 2.207459e-07, 2.219358e-07, 2.221972e-07, 2.224395e-07, 
    2.229179e-07, 2.235316e-07, 2.246076e-07, 2.255432e-07, 2.263969e-07, 
    2.263344e-07, 2.263564e-07, 2.26547e-07, 2.260748e-07, 2.266246e-07, 
    2.267168e-07, 2.264756e-07, 2.27875e-07, 2.274754e-07, 2.278843e-07, 
    2.276241e-07, 2.210686e-07, 2.213943e-07, 2.212183e-07, 2.215492e-07, 
    2.21316e-07, 2.223523e-07, 2.226628e-07, 2.241153e-07, 2.235195e-07, 
    2.244678e-07, 2.236159e-07, 2.237668e-07, 2.244985e-07, 2.236619e-07, 
    2.254916e-07, 2.242512e-07, 2.265544e-07, 2.253165e-07, 2.26632e-07, 
    2.263933e-07, 2.267885e-07, 2.271424e-07, 2.275877e-07, 2.284086e-07, 
    2.282185e-07, 2.289048e-07, 2.218797e-07, 2.223018e-07, 2.222647e-07, 
    2.227064e-07, 2.23033e-07, 2.237408e-07, 2.248751e-07, 2.244487e-07, 
    2.252315e-07, 2.253886e-07, 2.241993e-07, 2.249296e-07, 2.225843e-07, 
    2.229634e-07, 2.227378e-07, 2.219129e-07, 2.245468e-07, 2.231956e-07, 
    2.256899e-07, 2.249586e-07, 2.27092e-07, 2.260313e-07, 2.281139e-07, 
    2.29003e-07, 2.298397e-07, 2.308165e-07, 2.225323e-07, 2.222454e-07, 
    2.22759e-07, 2.234691e-07, 2.241279e-07, 2.250032e-07, 2.250928e-07, 
    2.252567e-07, 2.256812e-07, 2.26038e-07, 2.253084e-07, 2.261275e-07, 
    2.230512e-07, 2.246641e-07, 2.221369e-07, 2.228983e-07, 2.234273e-07, 
    2.231953e-07, 2.243999e-07, 2.246837e-07, 2.258362e-07, 2.252406e-07, 
    2.287836e-07, 2.272171e-07, 2.3156e-07, 2.303476e-07, 2.221452e-07, 
    2.225313e-07, 2.238742e-07, 2.232354e-07, 2.250617e-07, 2.255108e-07, 
    2.25876e-07, 2.263425e-07, 2.263929e-07, 2.266692e-07, 2.262163e-07, 
    2.266513e-07, 2.250051e-07, 2.25741e-07, 2.237208e-07, 2.242127e-07, 
    2.239864e-07, 2.237382e-07, 2.245043e-07, 2.253199e-07, 2.253374e-07, 
    2.255989e-07, 2.26335e-07, 2.250691e-07, 2.289854e-07, 2.265678e-07, 
    2.229522e-07, 2.236952e-07, 2.238015e-07, 2.235137e-07, 2.254658e-07, 
    2.247588e-07, 2.266625e-07, 2.261482e-07, 2.269907e-07, 2.265721e-07, 
    2.265105e-07, 2.259727e-07, 2.256377e-07, 2.247912e-07, 2.24102e-07, 
    2.235554e-07, 2.236825e-07, 2.242829e-07, 2.253698e-07, 2.263974e-07, 
    2.261723e-07, 2.269267e-07, 2.249293e-07, 2.257671e-07, 2.254433e-07, 
    2.262875e-07, 2.244373e-07, 2.260126e-07, 2.240344e-07, 2.242079e-07, 
    2.247447e-07, 2.258239e-07, 2.260627e-07, 2.263174e-07, 2.261603e-07, 
    2.253974e-07, 2.252724e-07, 2.247317e-07, 2.245823e-07, 2.241701e-07, 
    2.238288e-07, 2.241406e-07, 2.244681e-07, 2.253978e-07, 2.262351e-07, 
    2.271474e-07, 2.273707e-07, 2.284356e-07, 2.275687e-07, 2.289988e-07, 
    2.277828e-07, 2.298873e-07, 2.26104e-07, 2.277473e-07, 2.247692e-07, 
    2.250903e-07, 2.256708e-07, 2.270018e-07, 2.262835e-07, 2.271236e-07, 
    2.252675e-07, 2.243036e-07, 2.240542e-07, 2.235886e-07, 2.240649e-07, 
    2.240261e-07, 2.244817e-07, 2.243353e-07, 2.254286e-07, 2.248415e-07, 
    2.265089e-07, 2.27117e-07, 2.288329e-07, 2.298837e-07, 2.309527e-07, 
    2.314243e-07, 2.315679e-07, 2.316279e-07,
  2.107057e-07, 2.117065e-07, 2.11512e-07, 2.12319e-07, 2.118714e-07, 
    2.123998e-07, 2.109087e-07, 2.117462e-07, 2.112116e-07, 2.107959e-07, 
    2.13885e-07, 2.123551e-07, 2.154741e-07, 2.144986e-07, 2.16949e-07, 
    2.153223e-07, 2.17277e-07, 2.169021e-07, 2.180304e-07, 2.177072e-07, 
    2.1915e-07, 2.181795e-07, 2.198978e-07, 2.189183e-07, 2.190715e-07, 
    2.181475e-07, 2.12663e-07, 2.136945e-07, 2.126019e-07, 2.12749e-07, 
    2.12683e-07, 2.118806e-07, 2.114762e-07, 2.106293e-07, 2.10783e-07, 
    2.114051e-07, 2.128151e-07, 2.123365e-07, 2.135427e-07, 2.135155e-07, 
    2.148581e-07, 2.142528e-07, 2.165091e-07, 2.158679e-07, 2.177206e-07, 
    2.172547e-07, 2.176988e-07, 2.175641e-07, 2.177005e-07, 2.170172e-07, 
    2.1731e-07, 2.167087e-07, 2.143662e-07, 2.150547e-07, 2.13001e-07, 
    2.117658e-07, 2.109454e-07, 2.103631e-07, 2.104454e-07, 2.106024e-07, 
    2.114087e-07, 2.121668e-07, 2.127445e-07, 2.131309e-07, 2.135116e-07, 
    2.146637e-07, 2.152735e-07, 2.166387e-07, 2.163924e-07, 2.168097e-07, 
    2.172084e-07, 2.178776e-07, 2.177675e-07, 2.180623e-07, 2.167987e-07, 
    2.176385e-07, 2.162521e-07, 2.166313e-07, 2.136149e-07, 2.124657e-07, 
    2.11977e-07, 2.115493e-07, 2.105087e-07, 2.112274e-07, 2.109441e-07, 
    2.11618e-07, 2.120463e-07, 2.118345e-07, 2.131415e-07, 2.126334e-07, 
    2.153097e-07, 2.14157e-07, 2.171619e-07, 2.16443e-07, 2.173342e-07, 
    2.168794e-07, 2.176586e-07, 2.169574e-07, 2.181721e-07, 2.184366e-07, 
    2.182558e-07, 2.189501e-07, 2.169185e-07, 2.176987e-07, 2.118285e-07, 
    2.118631e-07, 2.12024e-07, 2.113166e-07, 2.112733e-07, 2.10625e-07, 
    2.112019e-07, 2.114475e-07, 2.120711e-07, 2.124399e-07, 2.127904e-07, 
    2.135612e-07, 2.144218e-07, 2.156251e-07, 2.164896e-07, 2.170689e-07, 
    2.167137e-07, 2.170273e-07, 2.166767e-07, 2.165124e-07, 2.183375e-07, 
    2.173127e-07, 2.188503e-07, 2.187652e-07, 2.180693e-07, 2.187748e-07, 
    2.118873e-07, 2.116886e-07, 2.109984e-07, 2.115385e-07, 2.105544e-07, 
    2.111053e-07, 2.11422e-07, 2.12644e-07, 2.129124e-07, 2.131613e-07, 
    2.136529e-07, 2.142838e-07, 2.153903e-07, 2.163529e-07, 2.172316e-07, 
    2.171672e-07, 2.171899e-07, 2.173861e-07, 2.169e-07, 2.17466e-07, 
    2.175609e-07, 2.173126e-07, 2.187538e-07, 2.183421e-07, 2.187634e-07, 
    2.184954e-07, 2.117532e-07, 2.120876e-07, 2.119069e-07, 2.122467e-07, 
    2.120073e-07, 2.130718e-07, 2.133909e-07, 2.148841e-07, 2.142714e-07, 
    2.152465e-07, 2.143704e-07, 2.145257e-07, 2.152782e-07, 2.144178e-07, 
    2.162998e-07, 2.150239e-07, 2.173938e-07, 2.161197e-07, 2.174736e-07, 
    2.172278e-07, 2.176348e-07, 2.179992e-07, 2.184578e-07, 2.193037e-07, 
    2.191078e-07, 2.198152e-07, 2.125862e-07, 2.130199e-07, 2.129818e-07, 
    2.134357e-07, 2.137713e-07, 2.144988e-07, 2.156655e-07, 2.152268e-07, 
    2.160321e-07, 2.161938e-07, 2.149703e-07, 2.157215e-07, 2.133102e-07, 
    2.136998e-07, 2.134679e-07, 2.126204e-07, 2.153278e-07, 2.139385e-07, 
    2.165038e-07, 2.157514e-07, 2.179473e-07, 2.168553e-07, 2.19e-07, 
    2.199166e-07, 2.207792e-07, 2.21787e-07, 2.132567e-07, 2.12962e-07, 
    2.134897e-07, 2.142196e-07, 2.148969e-07, 2.157972e-07, 2.158894e-07, 
    2.16058e-07, 2.164949e-07, 2.168621e-07, 2.161113e-07, 2.169542e-07, 
    2.137901e-07, 2.154484e-07, 2.128505e-07, 2.136329e-07, 2.141766e-07, 
    2.139381e-07, 2.151767e-07, 2.154685e-07, 2.166544e-07, 2.160414e-07, 
    2.196903e-07, 2.180762e-07, 2.225543e-07, 2.213032e-07, 2.12859e-07, 
    2.132557e-07, 2.14636e-07, 2.139793e-07, 2.158574e-07, 2.163195e-07, 
    2.166953e-07, 2.171755e-07, 2.172274e-07, 2.175119e-07, 2.170457e-07, 
    2.174935e-07, 2.157992e-07, 2.165564e-07, 2.144783e-07, 2.149841e-07, 
    2.147514e-07, 2.144962e-07, 2.15284e-07, 2.161231e-07, 2.161411e-07, 
    2.164101e-07, 2.171682e-07, 2.15865e-07, 2.198985e-07, 2.174077e-07, 
    2.136882e-07, 2.144521e-07, 2.145612e-07, 2.142653e-07, 2.162732e-07, 
    2.155457e-07, 2.17505e-07, 2.169755e-07, 2.17843e-07, 2.17412e-07, 
    2.173485e-07, 2.167949e-07, 2.164501e-07, 2.155791e-07, 2.148703e-07, 
    2.143083e-07, 2.14439e-07, 2.150564e-07, 2.161745e-07, 2.172321e-07, 
    2.170004e-07, 2.177771e-07, 2.157212e-07, 2.165833e-07, 2.162501e-07, 
    2.171189e-07, 2.152151e-07, 2.168362e-07, 2.148007e-07, 2.149792e-07, 
    2.155313e-07, 2.166418e-07, 2.168875e-07, 2.171497e-07, 2.169879e-07, 
    2.162028e-07, 2.160742e-07, 2.155179e-07, 2.153643e-07, 2.149403e-07, 
    2.145893e-07, 2.1491e-07, 2.152468e-07, 2.162032e-07, 2.17065e-07, 
    2.180044e-07, 2.182343e-07, 2.193317e-07, 2.184384e-07, 2.199124e-07, 
    2.186592e-07, 2.208285e-07, 2.169302e-07, 2.186224e-07, 2.155564e-07, 
    2.158868e-07, 2.164843e-07, 2.178545e-07, 2.171148e-07, 2.179799e-07, 
    2.160692e-07, 2.150776e-07, 2.148211e-07, 2.143424e-07, 2.148321e-07, 
    2.147923e-07, 2.152608e-07, 2.151102e-07, 2.16235e-07, 2.156308e-07, 
    2.173469e-07, 2.179731e-07, 2.197411e-07, 2.208246e-07, 2.219274e-07, 
    2.224142e-07, 2.225624e-07, 2.226243e-07,
  2.033617e-07, 2.043102e-07, 2.041257e-07, 2.048911e-07, 2.044665e-07, 
    2.049677e-07, 2.03554e-07, 2.043479e-07, 2.03841e-07, 2.034471e-07, 
    2.063778e-07, 2.049253e-07, 2.078882e-07, 2.069606e-07, 2.09292e-07, 
    2.077438e-07, 2.096044e-07, 2.092473e-07, 2.103224e-07, 2.100143e-07, 
    2.113905e-07, 2.104646e-07, 2.121045e-07, 2.111694e-07, 2.113156e-07, 
    2.104341e-07, 2.052174e-07, 2.061969e-07, 2.051594e-07, 2.05299e-07, 
    2.052364e-07, 2.044753e-07, 2.040919e-07, 2.032892e-07, 2.034349e-07, 
    2.040244e-07, 2.053618e-07, 2.049077e-07, 2.060525e-07, 2.060266e-07, 
    2.073023e-07, 2.06727e-07, 2.088731e-07, 2.082627e-07, 2.100272e-07, 
    2.095832e-07, 2.100063e-07, 2.09878e-07, 2.10008e-07, 2.093569e-07, 
    2.096358e-07, 2.090631e-07, 2.068347e-07, 2.074892e-07, 2.055382e-07, 
    2.043665e-07, 2.035888e-07, 2.030372e-07, 2.031151e-07, 2.032638e-07, 
    2.040279e-07, 2.047467e-07, 2.052948e-07, 2.056615e-07, 2.060229e-07, 
    2.071177e-07, 2.076974e-07, 2.089965e-07, 2.08762e-07, 2.091593e-07, 
    2.095391e-07, 2.101769e-07, 2.100719e-07, 2.103529e-07, 2.091488e-07, 
    2.09949e-07, 2.086284e-07, 2.089894e-07, 2.061213e-07, 2.050302e-07, 
    2.045668e-07, 2.041612e-07, 2.031751e-07, 2.03856e-07, 2.035875e-07, 
    2.042263e-07, 2.046323e-07, 2.044315e-07, 2.056715e-07, 2.051893e-07, 
    2.077318e-07, 2.06636e-07, 2.094948e-07, 2.088101e-07, 2.096589e-07, 
    2.092257e-07, 2.099681e-07, 2.092999e-07, 2.104576e-07, 2.107098e-07, 
    2.105374e-07, 2.111997e-07, 2.092629e-07, 2.100063e-07, 2.044259e-07, 
    2.044586e-07, 2.046112e-07, 2.039406e-07, 2.038996e-07, 2.032853e-07, 
    2.038318e-07, 2.040647e-07, 2.046559e-07, 2.050057e-07, 2.053384e-07, 
    2.0607e-07, 2.068877e-07, 2.080318e-07, 2.088545e-07, 2.094062e-07, 
    2.090678e-07, 2.093666e-07, 2.090326e-07, 2.088762e-07, 2.106153e-07, 
    2.096385e-07, 2.111044e-07, 2.110232e-07, 2.103596e-07, 2.110324e-07, 
    2.044816e-07, 2.042931e-07, 2.03639e-07, 2.041509e-07, 2.032184e-07, 
    2.037403e-07, 2.040405e-07, 2.051994e-07, 2.054541e-07, 2.056904e-07, 
    2.061572e-07, 2.067564e-07, 2.078084e-07, 2.087244e-07, 2.095612e-07, 
    2.094998e-07, 2.095214e-07, 2.097084e-07, 2.092453e-07, 2.097845e-07, 
    2.09875e-07, 2.096383e-07, 2.110124e-07, 2.106197e-07, 2.110215e-07, 
    2.107658e-07, 2.043544e-07, 2.046716e-07, 2.045002e-07, 2.048225e-07, 
    2.045954e-07, 2.056055e-07, 2.059084e-07, 2.073271e-07, 2.067447e-07, 
    2.076717e-07, 2.068388e-07, 2.069863e-07, 2.07702e-07, 2.068838e-07, 
    2.086739e-07, 2.0746e-07, 2.097157e-07, 2.085025e-07, 2.097918e-07, 
    2.095575e-07, 2.099453e-07, 2.102928e-07, 2.1073e-07, 2.115372e-07, 
    2.113502e-07, 2.120255e-07, 2.051445e-07, 2.055562e-07, 2.055199e-07, 
    2.059508e-07, 2.062696e-07, 2.069608e-07, 2.080702e-07, 2.076529e-07, 
    2.08419e-07, 2.085729e-07, 2.074089e-07, 2.081235e-07, 2.058318e-07, 
    2.062018e-07, 2.059814e-07, 2.05177e-07, 2.07749e-07, 2.064285e-07, 
    2.088681e-07, 2.081519e-07, 2.102432e-07, 2.092027e-07, 2.112473e-07, 
    2.121224e-07, 2.129465e-07, 2.139104e-07, 2.057809e-07, 2.055011e-07, 
    2.060021e-07, 2.066955e-07, 2.073392e-07, 2.081955e-07, 2.082832e-07, 
    2.084437e-07, 2.088595e-07, 2.092092e-07, 2.084944e-07, 2.092969e-07, 
    2.062876e-07, 2.078637e-07, 2.053954e-07, 2.061382e-07, 2.066546e-07, 
    2.06428e-07, 2.076052e-07, 2.078828e-07, 2.090115e-07, 2.084279e-07, 
    2.119064e-07, 2.103662e-07, 2.146447e-07, 2.134476e-07, 2.054034e-07, 
    2.057799e-07, 2.070912e-07, 2.064671e-07, 2.082527e-07, 2.086926e-07, 
    2.090503e-07, 2.095078e-07, 2.095571e-07, 2.098283e-07, 2.09384e-07, 
    2.098107e-07, 2.081974e-07, 2.089181e-07, 2.069413e-07, 2.074221e-07, 
    2.072009e-07, 2.069583e-07, 2.077072e-07, 2.085057e-07, 2.085227e-07, 
    2.087789e-07, 2.09501e-07, 2.0826e-07, 2.121054e-07, 2.097292e-07, 
    2.061906e-07, 2.069165e-07, 2.070201e-07, 2.067389e-07, 2.086485e-07, 
    2.079563e-07, 2.098216e-07, 2.093172e-07, 2.101438e-07, 2.09733e-07, 
    2.096726e-07, 2.091452e-07, 2.088169e-07, 2.07988e-07, 2.073139e-07, 
    2.067797e-07, 2.069039e-07, 2.074908e-07, 2.085546e-07, 2.095616e-07, 
    2.09341e-07, 2.10081e-07, 2.081232e-07, 2.089438e-07, 2.086265e-07, 
    2.094538e-07, 2.076418e-07, 2.091848e-07, 2.072477e-07, 2.074174e-07, 
    2.079425e-07, 2.089995e-07, 2.092334e-07, 2.094832e-07, 2.09329e-07, 
    2.085816e-07, 2.084591e-07, 2.079298e-07, 2.077836e-07, 2.073805e-07, 
    2.070468e-07, 2.073517e-07, 2.076719e-07, 2.085819e-07, 2.094025e-07, 
    2.102977e-07, 2.105169e-07, 2.11564e-07, 2.107116e-07, 2.121186e-07, 
    2.109224e-07, 2.129939e-07, 2.092742e-07, 2.108872e-07, 2.079664e-07, 
    2.082807e-07, 2.088495e-07, 2.101549e-07, 2.094499e-07, 2.102744e-07, 
    2.084543e-07, 2.075111e-07, 2.072671e-07, 2.068122e-07, 2.072776e-07, 
    2.072397e-07, 2.076852e-07, 2.07542e-07, 2.086121e-07, 2.080372e-07, 
    2.096711e-07, 2.102679e-07, 2.119547e-07, 2.1299e-07, 2.140447e-07, 
    2.145106e-07, 2.146525e-07, 2.147118e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.215762e-08, 6.243169e-08, 6.237841e-08, 6.259947e-08, 6.247685e-08, 
    6.26216e-08, 6.221319e-08, 6.244257e-08, 6.229614e-08, 6.21823e-08, 
    6.302847e-08, 6.260934e-08, 6.346394e-08, 6.319659e-08, 6.386823e-08, 
    6.342233e-08, 6.395815e-08, 6.385538e-08, 6.416472e-08, 6.40761e-08, 
    6.447177e-08, 6.420563e-08, 6.46769e-08, 6.440823e-08, 6.445025e-08, 
    6.419685e-08, 6.269369e-08, 6.297628e-08, 6.267695e-08, 6.271725e-08, 
    6.269916e-08, 6.247938e-08, 6.236861e-08, 6.213668e-08, 6.217878e-08, 
    6.234914e-08, 6.273537e-08, 6.260426e-08, 6.29347e-08, 6.292724e-08, 
    6.329513e-08, 6.312926e-08, 6.374764e-08, 6.357188e-08, 6.40798e-08, 
    6.395206e-08, 6.40738e-08, 6.403688e-08, 6.407428e-08, 6.388693e-08, 
    6.39672e-08, 6.380235e-08, 6.316031e-08, 6.334899e-08, 6.278628e-08, 
    6.244793e-08, 6.222324e-08, 6.20638e-08, 6.208634e-08, 6.212931e-08, 
    6.235014e-08, 6.255778e-08, 6.271602e-08, 6.282187e-08, 6.292617e-08, 
    6.324185e-08, 6.340898e-08, 6.378317e-08, 6.371565e-08, 6.383004e-08, 
    6.393935e-08, 6.412285e-08, 6.409265e-08, 6.417349e-08, 6.382704e-08, 
    6.405729e-08, 6.367719e-08, 6.378114e-08, 6.295448e-08, 6.263964e-08, 
    6.250578e-08, 6.238865e-08, 6.210367e-08, 6.230047e-08, 6.222289e-08, 
    6.240747e-08, 6.252476e-08, 6.246675e-08, 6.282476e-08, 6.268557e-08, 
    6.341888e-08, 6.310301e-08, 6.39266e-08, 6.372951e-08, 6.397384e-08, 
    6.384917e-08, 6.406279e-08, 6.387053e-08, 6.420358e-08, 6.427612e-08, 
    6.422655e-08, 6.441695e-08, 6.385987e-08, 6.40738e-08, 6.246512e-08, 
    6.247458e-08, 6.251866e-08, 6.232491e-08, 6.231306e-08, 6.213552e-08, 
    6.229349e-08, 6.236077e-08, 6.253156e-08, 6.263257e-08, 6.27286e-08, 
    6.293975e-08, 6.317556e-08, 6.350534e-08, 6.374228e-08, 6.390112e-08, 
    6.380372e-08, 6.388971e-08, 6.379359e-08, 6.374854e-08, 6.424895e-08, 
    6.396795e-08, 6.438957e-08, 6.436624e-08, 6.417542e-08, 6.436887e-08, 
    6.248122e-08, 6.242679e-08, 6.223777e-08, 6.238569e-08, 6.211619e-08, 
    6.226703e-08, 6.235377e-08, 6.268847e-08, 6.276202e-08, 6.283021e-08, 
    6.296489e-08, 6.313774e-08, 6.344097e-08, 6.370482e-08, 6.394571e-08, 
    6.392806e-08, 6.393427e-08, 6.398808e-08, 6.385479e-08, 6.400997e-08, 
    6.403601e-08, 6.396792e-08, 6.436311e-08, 6.425022e-08, 6.436574e-08, 
    6.429224e-08, 6.244449e-08, 6.253608e-08, 6.248658e-08, 6.257967e-08, 
    6.251409e-08, 6.280568e-08, 6.289311e-08, 6.330224e-08, 6.313434e-08, 
    6.340156e-08, 6.316149e-08, 6.320403e-08, 6.341026e-08, 6.317446e-08, 
    6.369027e-08, 6.334054e-08, 6.399017e-08, 6.36409e-08, 6.401206e-08, 
    6.394467e-08, 6.405626e-08, 6.415619e-08, 6.428195e-08, 6.451393e-08, 
    6.446022e-08, 6.465423e-08, 6.267265e-08, 6.279146e-08, 6.278102e-08, 
    6.290536e-08, 6.299733e-08, 6.319667e-08, 6.35164e-08, 6.339616e-08, 
    6.361689e-08, 6.366121e-08, 6.332587e-08, 6.353175e-08, 6.2871e-08, 
    6.297773e-08, 6.291419e-08, 6.268202e-08, 6.342385e-08, 6.304312e-08, 
    6.37462e-08, 6.353994e-08, 6.414194e-08, 6.384253e-08, 6.443064e-08, 
    6.468203e-08, 6.491868e-08, 6.51952e-08, 6.285632e-08, 6.277559e-08, 
    6.292016e-08, 6.312016e-08, 6.330577e-08, 6.355251e-08, 6.357777e-08, 
    6.362399e-08, 6.374373e-08, 6.384442e-08, 6.363859e-08, 6.386966e-08, 
    6.300247e-08, 6.345691e-08, 6.274506e-08, 6.295939e-08, 6.310837e-08, 
    6.304303e-08, 6.338242e-08, 6.346242e-08, 6.378748e-08, 6.361945e-08, 
    6.461998e-08, 6.417729e-08, 6.540579e-08, 6.506244e-08, 6.274738e-08, 
    6.285605e-08, 6.323427e-08, 6.305431e-08, 6.356899e-08, 6.369568e-08, 
    6.379868e-08, 6.393034e-08, 6.394456e-08, 6.402257e-08, 6.389474e-08, 
    6.401752e-08, 6.355304e-08, 6.37606e-08, 6.319105e-08, 6.332966e-08, 
    6.326589e-08, 6.319594e-08, 6.341183e-08, 6.364183e-08, 6.364677e-08, 
    6.372051e-08, 6.392831e-08, 6.357108e-08, 6.467708e-08, 6.399399e-08, 
    6.297455e-08, 6.318386e-08, 6.321378e-08, 6.313269e-08, 6.368298e-08, 
    6.348358e-08, 6.402067e-08, 6.387551e-08, 6.411335e-08, 6.399516e-08, 
    6.397777e-08, 6.382598e-08, 6.373148e-08, 6.349272e-08, 6.329847e-08, 
    6.314445e-08, 6.318027e-08, 6.334945e-08, 6.365591e-08, 6.394584e-08, 
    6.388233e-08, 6.409527e-08, 6.353167e-08, 6.376798e-08, 6.367664e-08, 
    6.391483e-08, 6.339297e-08, 6.383731e-08, 6.327939e-08, 6.332831e-08, 
    6.347963e-08, 6.378401e-08, 6.385137e-08, 6.392327e-08, 6.387891e-08, 
    6.366369e-08, 6.362843e-08, 6.347595e-08, 6.343384e-08, 6.331766e-08, 
    6.322146e-08, 6.330935e-08, 6.340164e-08, 6.366378e-08, 6.390003e-08, 
    6.415761e-08, 6.422066e-08, 6.452161e-08, 6.427662e-08, 6.468089e-08, 
    6.433715e-08, 6.493221e-08, 6.386308e-08, 6.432707e-08, 6.348652e-08, 
    6.357706e-08, 6.374083e-08, 6.41165e-08, 6.39137e-08, 6.415087e-08, 
    6.362706e-08, 6.335529e-08, 6.328499e-08, 6.315381e-08, 6.328799e-08, 
    6.327708e-08, 6.340547e-08, 6.336422e-08, 6.367249e-08, 6.35069e-08, 
    6.397733e-08, 6.414901e-08, 6.463389e-08, 6.493114e-08, 6.523376e-08, 
    6.536735e-08, 6.540802e-08, 6.542501e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  9.690869e-13, 9.717061e-13, 9.711974e-13, 9.733079e-13, 9.721376e-13, 
    9.735191e-13, 9.696185e-13, 9.718098e-13, 9.704114e-13, 9.693234e-13, 
    9.773974e-13, 9.734021e-13, 9.815437e-13, 9.790004e-13, 9.853853e-13, 
    9.811477e-13, 9.86239e-13, 9.852641e-13, 9.881991e-13, 9.873587e-13, 
    9.911072e-13, 9.885869e-13, 9.93049e-13, 9.90506e-13, 9.909036e-13, 
    9.885037e-13, 9.742074e-13, 9.769001e-13, 9.740476e-13, 9.744318e-13, 
    9.742596e-13, 9.721616e-13, 9.711031e-13, 9.688872e-13, 9.692898e-13, 
    9.709175e-13, 9.746046e-13, 9.733541e-13, 9.765059e-13, 9.764349e-13, 
    9.799384e-13, 9.783593e-13, 9.842408e-13, 9.825708e-13, 9.873939e-13, 
    9.861817e-13, 9.873367e-13, 9.869868e-13, 9.873413e-13, 9.855635e-13, 
    9.863253e-13, 9.847605e-13, 9.78655e-13, 9.804507e-13, 9.750905e-13, 
    9.718604e-13, 9.697145e-13, 9.6819e-13, 9.684057e-13, 9.688164e-13, 
    9.70927e-13, 9.729104e-13, 9.744206e-13, 9.754301e-13, 9.764246e-13, 
    9.7943e-13, 9.810209e-13, 9.845779e-13, 9.83937e-13, 9.85023e-13, 
    9.860612e-13, 9.87802e-13, 9.875156e-13, 9.88282e-13, 9.84995e-13, 
    9.871798e-13, 9.835717e-13, 9.845591e-13, 9.766921e-13, 9.736917e-13, 
    9.724129e-13, 9.712951e-13, 9.685714e-13, 9.704525e-13, 9.69711e-13, 
    9.714752e-13, 9.725951e-13, 9.720413e-13, 9.754578e-13, 9.741301e-13, 
    9.811151e-13, 9.78109e-13, 9.859402e-13, 9.840686e-13, 9.863886e-13, 
    9.852052e-13, 9.872322e-13, 9.85408e-13, 9.885674e-13, 9.892546e-13, 
    9.887849e-13, 9.90589e-13, 9.853068e-13, 9.873365e-13, 9.720257e-13, 
    9.721161e-13, 9.725369e-13, 9.70686e-13, 9.705728e-13, 9.68876e-13, 
    9.703861e-13, 9.710287e-13, 9.726602e-13, 9.736242e-13, 9.745404e-13, 
    9.765538e-13, 9.787998e-13, 9.819377e-13, 9.841899e-13, 9.856984e-13, 
    9.847737e-13, 9.855901e-13, 9.846774e-13, 9.842496e-13, 9.88997e-13, 
    9.863322e-13, 9.903297e-13, 9.901088e-13, 9.883002e-13, 9.901336e-13, 
    9.721795e-13, 9.716597e-13, 9.698534e-13, 9.712671e-13, 9.686912e-13, 
    9.70133e-13, 9.709616e-13, 9.741572e-13, 9.748594e-13, 9.755095e-13, 
    9.767935e-13, 9.784401e-13, 9.813257e-13, 9.838339e-13, 9.861217e-13, 
    9.859542e-13, 9.860131e-13, 9.865236e-13, 9.852585e-13, 9.867312e-13, 
    9.869781e-13, 9.863323e-13, 9.900791e-13, 9.890094e-13, 9.90104e-13, 
    9.894077e-13, 9.718287e-13, 9.727034e-13, 9.722308e-13, 9.731192e-13, 
    9.72493e-13, 9.752751e-13, 9.761085e-13, 9.800055e-13, 9.784076e-13, 
    9.809508e-13, 9.786663e-13, 9.790711e-13, 9.810325e-13, 9.7879e-13, 
    9.836951e-13, 9.803696e-13, 9.865434e-13, 9.832255e-13, 9.867512e-13, 
    9.861118e-13, 9.871705e-13, 9.88118e-13, 9.893101e-13, 9.915069e-13, 
    9.909985e-13, 9.928348e-13, 9.740068e-13, 9.751398e-13, 9.750406e-13, 
    9.762262e-13, 9.771025e-13, 9.790014e-13, 9.820431e-13, 9.808999e-13, 
    9.829987e-13, 9.834197e-13, 9.802312e-13, 9.821889e-13, 9.758982e-13, 
    9.769152e-13, 9.763101e-13, 9.740959e-13, 9.811626e-13, 9.775383e-13, 
    9.842271e-13, 9.82267e-13, 9.879829e-13, 9.851415e-13, 9.907185e-13, 
    9.930969e-13, 9.953354e-13, 9.979456e-13, 9.757585e-13, 9.749889e-13, 
    9.763673e-13, 9.782722e-13, 9.800396e-13, 9.823865e-13, 9.826268e-13, 
    9.830661e-13, 9.842039e-13, 9.8516e-13, 9.832044e-13, 9.853997e-13, 
    9.771499e-13, 9.814773e-13, 9.746973e-13, 9.767403e-13, 9.781602e-13, 
    9.775379e-13, 9.807693e-13, 9.815302e-13, 9.84619e-13, 9.83023e-13, 
    9.925097e-13, 9.883174e-13, 9.999327e-13, 9.966926e-13, 9.747198e-13, 
    9.757562e-13, 9.793588e-13, 9.776454e-13, 9.825434e-13, 9.837473e-13, 
    9.847259e-13, 9.859754e-13, 9.861106e-13, 9.868507e-13, 9.856378e-13, 
    9.86803e-13, 9.823915e-13, 9.84364e-13, 9.789479e-13, 9.80267e-13, 
    9.796605e-13, 9.789946e-13, 9.81049e-13, 9.832351e-13, 9.832826e-13, 
    9.839829e-13, 9.859539e-13, 9.825632e-13, 9.930485e-13, 9.865775e-13, 
    9.768857e-13, 9.788785e-13, 9.79164e-13, 9.783922e-13, 9.836265e-13, 
    9.817312e-13, 9.868328e-13, 9.854553e-13, 9.87712e-13, 9.865908e-13, 
    9.864258e-13, 9.84985e-13, 9.840873e-13, 9.818179e-13, 9.799701e-13, 
    9.785043e-13, 9.788453e-13, 9.804552e-13, 9.833689e-13, 9.861225e-13, 
    9.855195e-13, 9.875406e-13, 9.821886e-13, 9.844338e-13, 9.83566e-13, 
    9.858284e-13, 9.808694e-13, 9.850903e-13, 9.797888e-13, 9.802544e-13, 
    9.816936e-13, 9.845855e-13, 9.852261e-13, 9.859084e-13, 9.854876e-13, 
    9.834429e-13, 9.831082e-13, 9.816588e-13, 9.81258e-13, 9.801531e-13, 
    9.792375e-13, 9.800739e-13, 9.809516e-13, 9.834441e-13, 9.856877e-13, 
    9.881313e-13, 9.887294e-13, 9.915783e-13, 9.892584e-13, 9.930844e-13, 
    9.898302e-13, 9.954612e-13, 9.853359e-13, 9.897361e-13, 9.817593e-13, 
    9.826202e-13, 9.841756e-13, 9.877409e-13, 9.858178e-13, 9.880671e-13, 
    9.830951e-13, 9.805104e-13, 9.798422e-13, 9.785933e-13, 9.798707e-13, 
    9.797668e-13, 9.809886e-13, 9.805961e-13, 9.835268e-13, 9.819531e-13, 
    9.864214e-13, 9.880496e-13, 9.926422e-13, 9.954523e-13, 9.983104e-13, 
    9.995705e-13, 9.99954e-13, 1.000114e-12 ;

 LITR1C =
  3.066825e-05, 3.066813e-05, 3.066816e-05, 3.066806e-05, 3.066811e-05, 
    3.066805e-05, 3.066823e-05, 3.066813e-05, 3.066819e-05, 3.066824e-05, 
    3.066787e-05, 3.066806e-05, 3.066769e-05, 3.06678e-05, 3.066751e-05, 
    3.066771e-05, 3.066747e-05, 3.066752e-05, 3.066739e-05, 3.066742e-05, 
    3.066726e-05, 3.066737e-05, 3.066716e-05, 3.066728e-05, 3.066726e-05, 
    3.066737e-05, 3.066802e-05, 3.06679e-05, 3.066803e-05, 3.066801e-05, 
    3.066802e-05, 3.066811e-05, 3.066816e-05, 3.066826e-05, 3.066824e-05, 
    3.066817e-05, 3.0668e-05, 3.066806e-05, 3.066791e-05, 3.066792e-05, 
    3.066776e-05, 3.066783e-05, 3.066756e-05, 3.066764e-05, 3.066742e-05, 
    3.066748e-05, 3.066743e-05, 3.066744e-05, 3.066743e-05, 3.066751e-05, 
    3.066747e-05, 3.066754e-05, 3.066782e-05, 3.066774e-05, 3.066798e-05, 
    3.066812e-05, 3.066822e-05, 3.066829e-05, 3.066828e-05, 3.066826e-05, 
    3.066817e-05, 3.066808e-05, 3.066801e-05, 3.066796e-05, 3.066792e-05, 
    3.066778e-05, 3.066771e-05, 3.066755e-05, 3.066758e-05, 3.066753e-05, 
    3.066748e-05, 3.06674e-05, 3.066742e-05, 3.066738e-05, 3.066753e-05, 
    3.066743e-05, 3.066759e-05, 3.066755e-05, 3.066791e-05, 3.066804e-05, 
    3.06681e-05, 3.066815e-05, 3.066827e-05, 3.066819e-05, 3.066822e-05, 
    3.066814e-05, 3.066809e-05, 3.066812e-05, 3.066796e-05, 3.066802e-05, 
    3.066771e-05, 3.066784e-05, 3.066749e-05, 3.066757e-05, 3.066747e-05, 
    3.066752e-05, 3.066743e-05, 3.066751e-05, 3.066737e-05, 3.066734e-05, 
    3.066736e-05, 3.066728e-05, 3.066752e-05, 3.066743e-05, 3.066812e-05, 
    3.066811e-05, 3.06681e-05, 3.066818e-05, 3.066818e-05, 3.066826e-05, 
    3.066819e-05, 3.066816e-05, 3.066809e-05, 3.066804e-05, 3.0668e-05, 
    3.066791e-05, 3.066781e-05, 3.066767e-05, 3.066757e-05, 3.06675e-05, 
    3.066754e-05, 3.06675e-05, 3.066755e-05, 3.066756e-05, 3.066735e-05, 
    3.066747e-05, 3.066729e-05, 3.06673e-05, 3.066738e-05, 3.06673e-05, 
    3.066811e-05, 3.066814e-05, 3.066822e-05, 3.066815e-05, 3.066827e-05, 
    3.06682e-05, 3.066817e-05, 3.066802e-05, 3.066799e-05, 3.066796e-05, 
    3.06679e-05, 3.066783e-05, 3.06677e-05, 3.066758e-05, 3.066748e-05, 
    3.066749e-05, 3.066748e-05, 3.066746e-05, 3.066752e-05, 3.066745e-05, 
    3.066744e-05, 3.066747e-05, 3.06673e-05, 3.066735e-05, 3.06673e-05, 
    3.066733e-05, 3.066813e-05, 3.066809e-05, 3.066811e-05, 3.066807e-05, 
    3.06681e-05, 3.066797e-05, 3.066793e-05, 3.066776e-05, 3.066783e-05, 
    3.066771e-05, 3.066782e-05, 3.06678e-05, 3.066771e-05, 3.066781e-05, 
    3.066759e-05, 3.066774e-05, 3.066746e-05, 3.066761e-05, 3.066745e-05, 
    3.066748e-05, 3.066743e-05, 3.066739e-05, 3.066734e-05, 3.066724e-05, 
    3.066726e-05, 3.066718e-05, 3.066803e-05, 3.066798e-05, 3.066798e-05, 
    3.066793e-05, 3.066789e-05, 3.06678e-05, 3.066767e-05, 3.066772e-05, 
    3.066762e-05, 3.06676e-05, 3.066775e-05, 3.066766e-05, 3.066794e-05, 
    3.06679e-05, 3.066792e-05, 3.066803e-05, 3.06677e-05, 3.066787e-05, 
    3.066756e-05, 3.066766e-05, 3.06674e-05, 3.066752e-05, 3.066727e-05, 
    3.066716e-05, 3.066706e-05, 3.066694e-05, 3.066795e-05, 3.066798e-05, 
    3.066792e-05, 3.066783e-05, 3.066775e-05, 3.066765e-05, 3.066764e-05, 
    3.066762e-05, 3.066757e-05, 3.066752e-05, 3.066761e-05, 3.066751e-05, 
    3.066788e-05, 3.066769e-05, 3.0668e-05, 3.066791e-05, 3.066784e-05, 
    3.066787e-05, 3.066772e-05, 3.066769e-05, 3.066755e-05, 3.066762e-05, 
    3.066719e-05, 3.066738e-05, 3.066686e-05, 3.0667e-05, 3.0668e-05, 
    3.066795e-05, 3.066779e-05, 3.066786e-05, 3.066764e-05, 3.066759e-05, 
    3.066754e-05, 3.066749e-05, 3.066748e-05, 3.066745e-05, 3.06675e-05, 
    3.066745e-05, 3.066765e-05, 3.066756e-05, 3.06678e-05, 3.066775e-05, 
    3.066777e-05, 3.06678e-05, 3.066771e-05, 3.066761e-05, 3.066761e-05, 
    3.066758e-05, 3.066749e-05, 3.066764e-05, 3.066716e-05, 3.066746e-05, 
    3.06679e-05, 3.066781e-05, 3.066779e-05, 3.066783e-05, 3.066759e-05, 
    3.066768e-05, 3.066745e-05, 3.066751e-05, 3.066741e-05, 3.066746e-05, 
    3.066747e-05, 3.066753e-05, 3.066757e-05, 3.066767e-05, 3.066776e-05, 
    3.066783e-05, 3.066781e-05, 3.066774e-05, 3.06676e-05, 3.066748e-05, 
    3.066751e-05, 3.066742e-05, 3.066766e-05, 3.066756e-05, 3.06676e-05, 
    3.066749e-05, 3.066772e-05, 3.066753e-05, 3.066777e-05, 3.066775e-05, 
    3.066768e-05, 3.066755e-05, 3.066752e-05, 3.066749e-05, 3.066751e-05, 
    3.06676e-05, 3.066762e-05, 3.066768e-05, 3.06677e-05, 3.066775e-05, 
    3.066779e-05, 3.066775e-05, 3.066771e-05, 3.06676e-05, 3.06675e-05, 
    3.066739e-05, 3.066736e-05, 3.066723e-05, 3.066734e-05, 3.066716e-05, 
    3.066731e-05, 3.066706e-05, 3.066752e-05, 3.066732e-05, 3.066768e-05, 
    3.066764e-05, 3.066757e-05, 3.066741e-05, 3.06675e-05, 3.066739e-05, 
    3.066762e-05, 3.066774e-05, 3.066776e-05, 3.066782e-05, 3.066776e-05, 
    3.066777e-05, 3.066771e-05, 3.066773e-05, 3.06676e-05, 3.066767e-05, 
    3.066747e-05, 3.066739e-05, 3.066719e-05, 3.066706e-05, 3.066693e-05, 
    3.066687e-05, 3.066685e-05, 3.066684e-05 ;

 LITR1C_TO_SOIL1C =
  6.454541e-13, 6.471983e-13, 6.468595e-13, 6.482649e-13, 6.474856e-13, 
    6.484055e-13, 6.458081e-13, 6.472672e-13, 6.463361e-13, 6.456115e-13, 
    6.509882e-13, 6.483276e-13, 6.537493e-13, 6.520556e-13, 6.563074e-13, 
    6.534855e-13, 6.568759e-13, 6.562266e-13, 6.581812e-13, 6.576216e-13, 
    6.601176e-13, 6.584394e-13, 6.614108e-13, 6.597173e-13, 6.599822e-13, 
    6.583839e-13, 6.488639e-13, 6.50657e-13, 6.487575e-13, 6.490133e-13, 
    6.488987e-13, 6.475015e-13, 6.467967e-13, 6.453211e-13, 6.455892e-13, 
    6.466731e-13, 6.491284e-13, 6.482957e-13, 6.503945e-13, 6.503472e-13, 
    6.526802e-13, 6.516287e-13, 6.555452e-13, 6.544332e-13, 6.576449e-13, 
    6.568378e-13, 6.576069e-13, 6.573738e-13, 6.5761e-13, 6.564261e-13, 
    6.569334e-13, 6.558914e-13, 6.518256e-13, 6.530214e-13, 6.494519e-13, 
    6.47301e-13, 6.45872e-13, 6.448569e-13, 6.450004e-13, 6.452739e-13, 
    6.466794e-13, 6.480002e-13, 6.490059e-13, 6.496782e-13, 6.503404e-13, 
    6.523417e-13, 6.534011e-13, 6.557698e-13, 6.55343e-13, 6.560662e-13, 
    6.567575e-13, 6.579167e-13, 6.57726e-13, 6.582364e-13, 6.560475e-13, 
    6.575024e-13, 6.550998e-13, 6.557572e-13, 6.505185e-13, 6.485205e-13, 
    6.476689e-13, 6.469245e-13, 6.451108e-13, 6.463634e-13, 6.458697e-13, 
    6.470445e-13, 6.477903e-13, 6.474215e-13, 6.496966e-13, 6.488124e-13, 
    6.534639e-13, 6.51462e-13, 6.566769e-13, 6.554306e-13, 6.569755e-13, 
    6.561875e-13, 6.575373e-13, 6.563225e-13, 6.584264e-13, 6.58884e-13, 
    6.585713e-13, 6.597727e-13, 6.562552e-13, 6.576067e-13, 6.474111e-13, 
    6.474712e-13, 6.477515e-13, 6.465189e-13, 6.464436e-13, 6.453136e-13, 
    6.463193e-13, 6.467471e-13, 6.478336e-13, 6.484756e-13, 6.490857e-13, 
    6.504264e-13, 6.51922e-13, 6.540117e-13, 6.555115e-13, 6.565159e-13, 
    6.559001e-13, 6.564438e-13, 6.55836e-13, 6.555511e-13, 6.587125e-13, 
    6.56938e-13, 6.595999e-13, 6.594529e-13, 6.582485e-13, 6.594694e-13, 
    6.475135e-13, 6.471674e-13, 6.459645e-13, 6.469059e-13, 6.451906e-13, 
    6.461507e-13, 6.467024e-13, 6.488305e-13, 6.492981e-13, 6.49731e-13, 
    6.505861e-13, 6.516825e-13, 6.536041e-13, 6.552743e-13, 6.567978e-13, 
    6.566862e-13, 6.567255e-13, 6.570654e-13, 6.56223e-13, 6.572037e-13, 
    6.57368e-13, 6.56938e-13, 6.594331e-13, 6.587207e-13, 6.594497e-13, 
    6.58986e-13, 6.472799e-13, 6.478623e-13, 6.475476e-13, 6.481393e-13, 
    6.477223e-13, 6.495749e-13, 6.501299e-13, 6.527249e-13, 6.516609e-13, 
    6.533544e-13, 6.518331e-13, 6.521027e-13, 6.534089e-13, 6.519155e-13, 
    6.551819e-13, 6.529674e-13, 6.570787e-13, 6.548692e-13, 6.57217e-13, 
    6.567912e-13, 6.574962e-13, 6.581272e-13, 6.589209e-13, 6.603839e-13, 
    6.600453e-13, 6.612682e-13, 6.487303e-13, 6.494848e-13, 6.494187e-13, 
    6.502082e-13, 6.507918e-13, 6.520563e-13, 6.540818e-13, 6.533206e-13, 
    6.547182e-13, 6.549985e-13, 6.528752e-13, 6.541789e-13, 6.499898e-13, 
    6.50667e-13, 6.502641e-13, 6.487897e-13, 6.534955e-13, 6.51082e-13, 
    6.555362e-13, 6.542309e-13, 6.580372e-13, 6.561451e-13, 6.598588e-13, 
    6.614426e-13, 6.629333e-13, 6.646714e-13, 6.498968e-13, 6.493843e-13, 
    6.503022e-13, 6.515706e-13, 6.527477e-13, 6.543105e-13, 6.544705e-13, 
    6.54763e-13, 6.555207e-13, 6.561574e-13, 6.548551e-13, 6.56317e-13, 
    6.508234e-13, 6.53705e-13, 6.491902e-13, 6.505506e-13, 6.514961e-13, 
    6.510817e-13, 6.532336e-13, 6.537402e-13, 6.557971e-13, 6.547344e-13, 
    6.610516e-13, 6.5826e-13, 6.659947e-13, 6.638371e-13, 6.492051e-13, 
    6.498952e-13, 6.522943e-13, 6.511533e-13, 6.544149e-13, 6.552166e-13, 
    6.558683e-13, 6.567004e-13, 6.567904e-13, 6.572832e-13, 6.564756e-13, 
    6.572515e-13, 6.543138e-13, 6.556273e-13, 6.520206e-13, 6.528991e-13, 
    6.524951e-13, 6.520517e-13, 6.534199e-13, 6.548755e-13, 6.549072e-13, 
    6.553735e-13, 6.566861e-13, 6.544282e-13, 6.614105e-13, 6.571013e-13, 
    6.506474e-13, 6.519745e-13, 6.521646e-13, 6.516506e-13, 6.551362e-13, 
    6.538741e-13, 6.572713e-13, 6.56354e-13, 6.578568e-13, 6.571102e-13, 
    6.570003e-13, 6.560408e-13, 6.55443e-13, 6.539319e-13, 6.527014e-13, 
    6.517253e-13, 6.519523e-13, 6.530245e-13, 6.549647e-13, 6.567983e-13, 
    6.563968e-13, 6.577426e-13, 6.541787e-13, 6.556738e-13, 6.550959e-13, 
    6.566024e-13, 6.533002e-13, 6.56111e-13, 6.525807e-13, 6.528907e-13, 
    6.53849e-13, 6.557748e-13, 6.562014e-13, 6.566557e-13, 6.563755e-13, 
    6.55014e-13, 6.547911e-13, 6.538259e-13, 6.53559e-13, 6.528232e-13, 
    6.522135e-13, 6.527705e-13, 6.53355e-13, 6.550148e-13, 6.565088e-13, 
    6.581361e-13, 6.585343e-13, 6.604315e-13, 6.588865e-13, 6.614343e-13, 
    6.592673e-13, 6.630171e-13, 6.562746e-13, 6.592047e-13, 6.538928e-13, 
    6.544661e-13, 6.555019e-13, 6.57876e-13, 6.565954e-13, 6.580933e-13, 
    6.547824e-13, 6.530612e-13, 6.526161e-13, 6.517845e-13, 6.526352e-13, 
    6.52566e-13, 6.533796e-13, 6.531182e-13, 6.550699e-13, 6.540219e-13, 
    6.569974e-13, 6.580816e-13, 6.611399e-13, 6.630111e-13, 6.649144e-13, 
    6.657535e-13, 6.660089e-13, 6.661156e-13 ;

 LITR1C_vr =
  0.001751189, 0.001751182, 0.001751183, 0.001751178, 0.001751181, 
    0.001751177, 0.001751187, 0.001751182, 0.001751185, 0.001751188, 
    0.001751167, 0.001751178, 0.001751157, 0.001751163, 0.001751147, 
    0.001751158, 0.001751145, 0.001751147, 0.001751139, 0.001751142, 
    0.001751132, 0.001751138, 0.001751127, 0.001751133, 0.001751132, 
    0.001751139, 0.001751176, 0.001751169, 0.001751176, 0.001751175, 
    0.001751175, 0.001751181, 0.001751184, 0.001751189, 0.001751188, 
    0.001751184, 0.001751175, 0.001751178, 0.00175117, 0.00175117, 
    0.001751161, 0.001751165, 0.00175115, 0.001751154, 0.001751142, 
    0.001751145, 0.001751142, 0.001751143, 0.001751142, 0.001751146, 
    0.001751144, 0.001751148, 0.001751164, 0.001751159, 0.001751173, 
    0.001751182, 0.001751187, 0.001751191, 0.001751191, 0.00175119, 
    0.001751184, 0.001751179, 0.001751175, 0.001751172, 0.00175117, 
    0.001751162, 0.001751158, 0.001751149, 0.00175115, 0.001751148, 
    0.001751145, 0.00175114, 0.001751141, 0.001751139, 0.001751148, 
    0.001751142, 0.001751151, 0.001751149, 0.001751169, 0.001751177, 
    0.00175118, 0.001751183, 0.00175119, 0.001751185, 0.001751187, 
    0.001751183, 0.00175118, 0.001751181, 0.001751172, 0.001751176, 
    0.001751158, 0.001751165, 0.001751145, 0.00175115, 0.001751144, 
    0.001751147, 0.001751142, 0.001751147, 0.001751138, 0.001751137, 
    0.001751138, 0.001751133, 0.001751147, 0.001751142, 0.001751181, 
    0.001751181, 0.00175118, 0.001751185, 0.001751185, 0.001751189, 
    0.001751186, 0.001751184, 0.00175118, 0.001751177, 0.001751175, 
    0.00175117, 0.001751164, 0.001751156, 0.00175115, 0.001751146, 
    0.001751148, 0.001751146, 0.001751148, 0.00175115, 0.001751137, 
    0.001751144, 0.001751134, 0.001751135, 0.001751139, 0.001751134, 
    0.001751181, 0.001751182, 0.001751187, 0.001751183, 0.00175119, 
    0.001751186, 0.001751184, 0.001751176, 0.001751174, 0.001751172, 
    0.001751169, 0.001751165, 0.001751157, 0.001751151, 0.001751145, 
    0.001751145, 0.001751145, 0.001751144, 0.001751147, 0.001751143, 
    0.001751143, 0.001751144, 0.001751135, 0.001751137, 0.001751135, 
    0.001751136, 0.001751182, 0.00175118, 0.001751181, 0.001751178, 
    0.00175118, 0.001751173, 0.001751171, 0.001751161, 0.001751165, 
    0.001751158, 0.001751164, 0.001751163, 0.001751158, 0.001751164, 
    0.001751151, 0.00175116, 0.001751144, 0.001751152, 0.001751143, 
    0.001751145, 0.001751142, 0.00175114, 0.001751137, 0.001751131, 
    0.001751132, 0.001751127, 0.001751176, 0.001751173, 0.001751174, 
    0.00175117, 0.001751168, 0.001751163, 0.001751155, 0.001751158, 
    0.001751153, 0.001751152, 0.00175116, 0.001751155, 0.001751171, 
    0.001751169, 0.00175117, 0.001751176, 0.001751158, 0.001751167, 
    0.00175115, 0.001751155, 0.00175114, 0.001751147, 0.001751133, 
    0.001751127, 0.001751121, 0.001751114, 0.001751172, 0.001751174, 
    0.00175117, 0.001751165, 0.00175116, 0.001751154, 0.001751154, 
    0.001751153, 0.00175115, 0.001751147, 0.001751152, 0.001751147, 
    0.001751168, 0.001751157, 0.001751174, 0.001751169, 0.001751165, 
    0.001751167, 0.001751159, 0.001751157, 0.001751149, 0.001751153, 
    0.001751128, 0.001751139, 0.001751109, 0.001751117, 0.001751174, 
    0.001751172, 0.001751162, 0.001751167, 0.001751154, 0.001751151, 
    0.001751148, 0.001751145, 0.001751145, 0.001751143, 0.001751146, 
    0.001751143, 0.001751154, 0.001751149, 0.001751163, 0.00175116, 
    0.001751162, 0.001751163, 0.001751158, 0.001751152, 0.001751152, 
    0.00175115, 0.001751145, 0.001751154, 0.001751127, 0.001751144, 
    0.001751169, 0.001751164, 0.001751163, 0.001751165, 0.001751151, 
    0.001751156, 0.001751143, 0.001751147, 0.001751141, 0.001751144, 
    0.001751144, 0.001751148, 0.00175115, 0.001751156, 0.001751161, 
    0.001751165, 0.001751164, 0.001751159, 0.001751152, 0.001751145, 
    0.001751146, 0.001751141, 0.001751155, 0.001751149, 0.001751151, 
    0.001751146, 0.001751158, 0.001751147, 0.001751161, 0.00175116, 
    0.001751156, 0.001751149, 0.001751147, 0.001751145, 0.001751146, 
    0.001751152, 0.001751153, 0.001751156, 0.001751157, 0.00175116, 
    0.001751163, 0.00175116, 0.001751158, 0.001751152, 0.001751146, 
    0.00175114, 0.001751138, 0.001751131, 0.001751137, 0.001751127, 
    0.001751135, 0.001751121, 0.001751147, 0.001751135, 0.001751156, 
    0.001751154, 0.00175115, 0.001751141, 0.001751146, 0.00175114, 
    0.001751153, 0.001751159, 0.001751161, 0.001751164, 0.001751161, 
    0.001751161, 0.001751158, 0.001751159, 0.001751152, 0.001751156, 
    0.001751144, 0.00175114, 0.001751128, 0.001751121, 0.001751113, 
    0.00175111, 0.001751109, 0.001751109,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.732964e-07, 9.732926e-07, 9.732934e-07, 9.732903e-07, 9.73292e-07, 
    9.732901e-07, 9.732956e-07, 9.732925e-07, 9.732945e-07, 9.732961e-07, 
    9.732845e-07, 9.732902e-07, 9.732785e-07, 9.732821e-07, 9.732729e-07, 
    9.73279e-07, 9.732718e-07, 9.732731e-07, 9.732689e-07, 9.732701e-07, 
    9.732647e-07, 9.732684e-07, 9.73262e-07, 9.732656e-07, 9.732651e-07, 
    9.732685e-07, 9.73289e-07, 9.732852e-07, 9.732893e-07, 9.732887e-07, 
    9.732889e-07, 9.73292e-07, 9.732935e-07, 9.732967e-07, 9.732961e-07, 
    9.732937e-07, 9.732885e-07, 9.732903e-07, 9.732858e-07, 9.732859e-07, 
    9.732807e-07, 9.73283e-07, 9.732746e-07, 9.73277e-07, 9.732701e-07, 
    9.732718e-07, 9.732702e-07, 9.732706e-07, 9.732702e-07, 9.732727e-07, 
    9.732717e-07, 9.732738e-07, 9.732827e-07, 9.732801e-07, 9.732878e-07, 
    9.732925e-07, 9.732955e-07, 9.732977e-07, 9.732973e-07, 9.732968e-07, 
    9.732937e-07, 9.732909e-07, 9.732887e-07, 9.732872e-07, 9.732859e-07, 
    9.732815e-07, 9.732793e-07, 9.732742e-07, 9.732751e-07, 9.732735e-07, 
    9.73272e-07, 9.732695e-07, 9.732699e-07, 9.732688e-07, 9.732735e-07, 
    9.732704e-07, 9.732755e-07, 9.732742e-07, 9.732854e-07, 9.732897e-07, 
    9.732917e-07, 9.732933e-07, 9.732971e-07, 9.732944e-07, 9.732955e-07, 
    9.732929e-07, 9.732913e-07, 9.732921e-07, 9.732872e-07, 9.732892e-07, 
    9.73279e-07, 9.732834e-07, 9.732721e-07, 9.732748e-07, 9.732715e-07, 
    9.732732e-07, 9.732703e-07, 9.732729e-07, 9.732684e-07, 9.732674e-07, 
    9.73268e-07, 9.732655e-07, 9.73273e-07, 9.732702e-07, 9.732921e-07, 
    9.73292e-07, 9.732914e-07, 9.73294e-07, 9.732943e-07, 9.732967e-07, 
    9.732945e-07, 9.732936e-07, 9.732912e-07, 9.732898e-07, 9.732886e-07, 
    9.732856e-07, 9.732825e-07, 9.732779e-07, 9.732747e-07, 9.732724e-07, 
    9.732738e-07, 9.732727e-07, 9.732739e-07, 9.732746e-07, 9.732678e-07, 
    9.732715e-07, 9.732659e-07, 9.732662e-07, 9.732688e-07, 9.732661e-07, 
    9.732919e-07, 9.732927e-07, 9.732953e-07, 9.732933e-07, 9.73297e-07, 
    9.732948e-07, 9.732937e-07, 9.73289e-07, 9.732881e-07, 9.732871e-07, 
    9.732853e-07, 9.732829e-07, 9.732788e-07, 9.732752e-07, 9.732719e-07, 
    9.732721e-07, 9.732721e-07, 9.732713e-07, 9.732731e-07, 9.73271e-07, 
    9.732706e-07, 9.732715e-07, 9.732662e-07, 9.732678e-07, 9.732662e-07, 
    9.732672e-07, 9.732925e-07, 9.732912e-07, 9.732919e-07, 9.732906e-07, 
    9.732915e-07, 9.732875e-07, 9.732863e-07, 9.732807e-07, 9.73283e-07, 
    9.732794e-07, 9.732826e-07, 9.73282e-07, 9.732793e-07, 9.732825e-07, 
    9.732754e-07, 9.732802e-07, 9.732713e-07, 9.732761e-07, 9.73271e-07, 
    9.732719e-07, 9.732704e-07, 9.73269e-07, 9.732673e-07, 9.732642e-07, 
    9.732648e-07, 9.732622e-07, 9.732893e-07, 9.732877e-07, 9.732878e-07, 
    9.732861e-07, 9.732848e-07, 9.732821e-07, 9.732778e-07, 9.732794e-07, 
    9.732764e-07, 9.732757e-07, 9.732804e-07, 9.732776e-07, 9.732865e-07, 
    9.732852e-07, 9.73286e-07, 9.732892e-07, 9.73279e-07, 9.732843e-07, 
    9.732746e-07, 9.732775e-07, 9.732693e-07, 9.732734e-07, 9.732653e-07, 
    9.732619e-07, 9.732587e-07, 9.732549e-07, 9.732868e-07, 9.732879e-07, 
    9.73286e-07, 9.732831e-07, 9.732806e-07, 9.732772e-07, 9.732769e-07, 
    9.732763e-07, 9.732746e-07, 9.732732e-07, 9.732761e-07, 9.732729e-07, 
    9.732848e-07, 9.732786e-07, 9.732884e-07, 9.732854e-07, 9.732834e-07, 
    9.732843e-07, 9.732796e-07, 9.732785e-07, 9.73274e-07, 9.732763e-07, 
    9.732627e-07, 9.732687e-07, 9.73252e-07, 9.732566e-07, 9.732883e-07, 
    9.732868e-07, 9.732817e-07, 9.73284e-07, 9.73277e-07, 9.732753e-07, 
    9.732739e-07, 9.732721e-07, 9.732719e-07, 9.732709e-07, 9.732726e-07, 
    9.73271e-07, 9.732772e-07, 9.732744e-07, 9.732822e-07, 9.732803e-07, 
    9.732812e-07, 9.732821e-07, 9.732792e-07, 9.732761e-07, 9.73276e-07, 
    9.73275e-07, 9.732721e-07, 9.73277e-07, 9.73262e-07, 9.732712e-07, 
    9.732852e-07, 9.732823e-07, 9.732819e-07, 9.73283e-07, 9.732755e-07, 
    9.732782e-07, 9.732709e-07, 9.732729e-07, 9.732696e-07, 9.732712e-07, 
    9.732714e-07, 9.732736e-07, 9.732748e-07, 9.732781e-07, 9.732807e-07, 
    9.732828e-07, 9.732823e-07, 9.732801e-07, 9.732759e-07, 9.732719e-07, 
    9.732728e-07, 9.732698e-07, 9.732776e-07, 9.732743e-07, 9.732755e-07, 
    9.732723e-07, 9.732795e-07, 9.732734e-07, 9.73281e-07, 9.732803e-07, 
    9.732782e-07, 9.732742e-07, 9.732731e-07, 9.732722e-07, 9.732728e-07, 
    9.732757e-07, 9.732762e-07, 9.732784e-07, 9.732789e-07, 9.732805e-07, 
    9.732818e-07, 9.732806e-07, 9.732794e-07, 9.732757e-07, 9.732726e-07, 
    9.73269e-07, 9.732681e-07, 9.73264e-07, 9.732673e-07, 9.732619e-07, 
    9.732665e-07, 9.732585e-07, 9.73273e-07, 9.732667e-07, 9.732781e-07, 
    9.732769e-07, 9.732747e-07, 9.732696e-07, 9.732723e-07, 9.732692e-07, 
    9.732762e-07, 9.7328e-07, 9.73281e-07, 9.732827e-07, 9.732809e-07, 
    9.732811e-07, 9.732793e-07, 9.732798e-07, 9.732756e-07, 9.732779e-07, 
    9.732714e-07, 9.732692e-07, 9.732626e-07, 9.732585e-07, 9.732544e-07, 
    9.732526e-07, 9.73252e-07, 9.732518e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  1.225453e-25, 2.794032e-25, -1.519561e-25, 1.56858e-25, -5.882173e-26, 
    1.960724e-26, -5.293956e-25, -5.784137e-25, -1.81367e-25, 4.999847e-25, 
    -5.931191e-25, 7.156644e-25, -3.137159e-25, 1.274471e-25, -4.803775e-25, 
    1.862688e-25, -1.470543e-25, 8.82326e-26, 5.931191e-25, -4.068503e-25, 
    -1.960724e-25, 3.774394e-25, 6.862535e-26, 5.097883e-25, -7.352717e-25, 
    1.764652e-25, 4.901811e-26, -4.999847e-25, -3.431268e-25, -2.352869e-25, 
    -4.313593e-25, 1.960724e-26, 6.078246e-25, -1.176435e-25, 4.901811e-26, 
    2.941087e-26, 1.960724e-26, 4.019485e-25, 4.999847e-25, -1.0833e-24, 
    -1.666616e-25, 7.058608e-25, 3.529304e-25, 7.058608e-25, 6.862535e-26, 
    7.499771e-25, 3.921449e-26, 1.372507e-25, 1.960724e-25, -5.490028e-25, 
    -9.803622e-27, -8.431115e-25, 6.862535e-26, -2.892069e-25, -5.882173e-26, 
    4.607703e-25, -1.764652e-25, 5.391992e-26, 1.176435e-25, -3.284213e-25, 
    -2.352869e-25, -6.862535e-26, -5.588064e-25, -1.078398e-25, 6.568427e-25, 
    -6.078246e-25, -1.911706e-25, 7.352717e-25, 2.695996e-25, 5.097883e-25, 
    2.254833e-25, 4.509666e-25, -4.607703e-25, 1.24506e-24, -1.666616e-25, 
    -4.117521e-25, 1.862688e-25, 2.548942e-25, -1.078398e-25, -3.823413e-25, 
    -5.686101e-25, -8.235043e-25, 5.097883e-25, -1.960724e-26, -6.519409e-25, 
    6.372354e-25, -9.803622e-27, 2.941087e-25, 2.107779e-25, 3.921449e-26, 
    2.745014e-25, 1.132318e-24, 2.254833e-25, 3.088141e-25, 2.548942e-25, 
    7.107626e-25, 9.803622e-26, -5.391992e-26, -4.607703e-25, -2.254833e-25, 
    1.02938e-25, -5.19592e-25, -8.235043e-25, -3.235195e-25, 6.568427e-25, 
    -7.842898e-26, -4.754757e-25, -1.960724e-26, 2.450905e-26, -1.81367e-25, 
    1.058791e-24, -2.058761e-25, 1.274471e-25, 3.333231e-25, 7.744861e-25, 
    3.823413e-25, -3.921449e-25, 6.862535e-26, -3.039123e-25, 1.274471e-25, 
    6.568427e-25, -1.176435e-25, 3.431268e-25, -1.274471e-25, -1.470543e-25, 
    1.078398e-25, 4.901811e-26, 2.058761e-25, -9.803622e-27, -9.803622e-27, 
    6.176282e-25, 3.235195e-25, 7.842898e-26, -6.617445e-25, -7.842898e-26, 
    7.450753e-25, 8.627187e-25, -1.960724e-25, 4.754757e-25, 1.274471e-25, 
    2.646978e-25, -2.156797e-25, -3.431268e-25, 2.303851e-25, 4.901811e-25, 
    1.274471e-25, 3.725376e-25, 3.235195e-25, 2.794032e-25, 5.391992e-25, 
    -4.950829e-25, 3.431268e-25, -2.058761e-25, 4.607703e-25, -5.784137e-25, 
    -3.284213e-25, -9.803622e-26, 5.391992e-26, 5.833155e-25, 2.009742e-25, 
    1.960724e-26, 8.333079e-25, 1.519561e-25, 6.862535e-26, -1.960724e-25, 
    1.274471e-25, 4.558684e-25, 2.548942e-25, -5.931191e-25, 7.352717e-25, 
    7.989952e-25, 1.372507e-25, -5.686101e-25, -4.264576e-25, -7.352717e-26, 
    -3.137159e-25, 3.578322e-25, 1.470543e-25, 4.803775e-25, 1.470543e-25, 
    -5.882173e-25, -8.186024e-25, -7.842898e-26, -1.960724e-25, 2.303851e-25, 
    -4.41163e-26, 5.784137e-25, -1.862688e-25, 3.235195e-25, -1.56858e-25, 
    7.842898e-26, 2.843051e-25, 2.548942e-25, -6.764499e-25, -7.352717e-26, 
    6.078246e-25, -3.578322e-25, 1.176435e-25, -7.00959e-25, 3.137159e-25, 
    4.803775e-25, -4.215557e-25, -5.097883e-25, 4.901811e-26, 2.59796e-25, 
    -2.941087e-26, 3.62734e-25, -9.117368e-25, -3.62734e-25, 3.872431e-25, 
    9.803622e-27, -3.284213e-25, 1.56858e-25, -1.357802e-24, -2.548942e-25, 
    -5.44101e-25, -7.891916e-25, 4.558684e-25, -3.921449e-26, 9.509513e-25, 
    3.333231e-25, 6.862535e-26, 1.13722e-24, 2.941087e-26, 9.803622e-27, 
    2.745014e-25, -4.803775e-25, -2.156797e-25, -1.323489e-25, -6.862535e-25, 
    7.842898e-25, -4.901811e-25, -2.352869e-25, 7.695843e-25, -1.117613e-24, 
    -3.088141e-25, -2.156797e-25, -9.803622e-27, 4.41163e-25, -5.588064e-25, 
    6.568427e-25, -1.764652e-25, -9.803622e-27, 4.558684e-25, -2.695996e-25, 
    -3.725376e-25, 9.803622e-26, -4.117521e-25, 7.646825e-25, 3.529304e-25, 
    6.078246e-25, -9.803622e-26, -1.960724e-26, 4.607703e-25, -2.59796e-25, 
    4.41163e-25, 1.56858e-25, 5.882173e-26, -3.529304e-25, 9.901658e-25, 
    1.078398e-25, 6.47039e-25, 1.078398e-25, -5.588064e-25, 2.892069e-25, 
    1.470543e-25, 7.842898e-26, -2.646978e-25, 4.313593e-25, 3.62734e-25, 
    -3.137159e-25, -4.705739e-25, 5.342974e-25, -9.803622e-26, 6.862535e-26, 
    8.333079e-26, 1.176435e-25, 8.82326e-26, -2.794032e-25, 4.509666e-25, 
    -1.176435e-25, -9.313441e-26, 4.362612e-25, 3.529304e-25, -4.607703e-25, 
    2.941087e-26, 7.156644e-25, -1.323489e-25, -4.41163e-26, -3.921449e-26, 
    1.372507e-25, 3.921449e-25, -9.803622e-26, -7.25468e-25, 2.352869e-25, 
    -4.901811e-26, 5.19592e-25, 1.009773e-24, 6.47039e-25, -1.56858e-25, 
    -3.333231e-25, -8.82326e-26, 1.764652e-25, 4.803775e-25, -7.303698e-25, 
    6.176282e-25, 6.372354e-25, -7.744861e-25, 1.127417e-25, -3.921449e-25, 
    8.676206e-25, 6.372354e-26, 9.313441e-26, -5.98021e-25, 5.882173e-26, 
    2.499924e-25, -1.56858e-25, -9.60755e-25, 6.029227e-25, 3.62734e-25, 
    2.548942e-25, 1.200944e-24, 3.333231e-25, -1.470543e-25, -9.803622e-27, 
    5.588064e-25, 2.745014e-25, 5.490028e-25, -3.921449e-26, 9.803622e-26, 
    -3.088141e-25, 1.470543e-25, 7.25468e-25, 2.745014e-25, -1.421525e-25, 
    7.842898e-26, 5.882173e-25, -3.333231e-25,
  9.436804e-32, 9.436766e-32, 9.436773e-32, 9.436743e-32, 9.43676e-32, 
    9.43674e-32, 9.436796e-32, 9.436765e-32, 9.436785e-32, 9.4368e-32, 
    9.436684e-32, 9.436742e-32, 9.436624e-32, 9.436661e-32, 9.436569e-32, 
    9.43663e-32, 9.436557e-32, 9.436571e-32, 9.436528e-32, 9.43654e-32, 
    9.436486e-32, 9.436522e-32, 9.436458e-32, 9.436495e-32, 9.436489e-32, 
    9.436524e-32, 9.43673e-32, 9.436691e-32, 9.436732e-32, 9.436727e-32, 
    9.436729e-32, 9.43676e-32, 9.436775e-32, 9.436807e-32, 9.436801e-32, 
    9.436778e-32, 9.436725e-32, 9.436742e-32, 9.436697e-32, 9.436698e-32, 
    9.436647e-32, 9.43667e-32, 9.436585e-32, 9.436609e-32, 9.43654e-32, 
    9.436557e-32, 9.436541e-32, 9.436545e-32, 9.43654e-32, 9.436566e-32, 
    9.436555e-32, 9.436578e-32, 9.436666e-32, 9.43664e-32, 9.436718e-32, 
    9.436764e-32, 9.436795e-32, 9.436817e-32, 9.436814e-32, 9.436808e-32, 
    9.436778e-32, 9.436749e-32, 9.436727e-32, 9.436712e-32, 9.436698e-32, 
    9.436655e-32, 9.436632e-32, 9.43658e-32, 9.436589e-32, 9.436574e-32, 
    9.436559e-32, 9.436534e-32, 9.436538e-32, 9.436527e-32, 9.436574e-32, 
    9.436542e-32, 9.436595e-32, 9.436581e-32, 9.436694e-32, 9.436738e-32, 
    9.436756e-32, 9.436772e-32, 9.436812e-32, 9.436785e-32, 9.436795e-32, 
    9.436769e-32, 9.436753e-32, 9.436762e-32, 9.436712e-32, 9.436731e-32, 
    9.436631e-32, 9.436674e-32, 9.436561e-32, 9.436588e-32, 9.436554e-32, 
    9.436571e-32, 9.436542e-32, 9.436568e-32, 9.436522e-32, 9.436512e-32, 
    9.43652e-32, 9.436494e-32, 9.436569e-32, 9.436541e-32, 9.436762e-32, 
    9.436761e-32, 9.436754e-32, 9.436781e-32, 9.436783e-32, 9.436807e-32, 
    9.436785e-32, 9.436776e-32, 9.436752e-32, 9.436739e-32, 9.436725e-32, 
    9.436696e-32, 9.436664e-32, 9.436618e-32, 9.436586e-32, 9.436564e-32, 
    9.436578e-32, 9.436566e-32, 9.436579e-32, 9.436585e-32, 9.436517e-32, 
    9.436555e-32, 9.436497e-32, 9.4365e-32, 9.436527e-32, 9.4365e-32, 
    9.436759e-32, 9.436767e-32, 9.436793e-32, 9.436773e-32, 9.43681e-32, 
    9.436789e-32, 9.436777e-32, 9.436731e-32, 9.436721e-32, 9.436711e-32, 
    9.436693e-32, 9.436669e-32, 9.436627e-32, 9.436591e-32, 9.436558e-32, 
    9.436561e-32, 9.436559e-32, 9.436552e-32, 9.436571e-32, 9.436549e-32, 
    9.436545e-32, 9.436555e-32, 9.436501e-32, 9.436516e-32, 9.436501e-32, 
    9.436511e-32, 9.436765e-32, 9.436752e-32, 9.436759e-32, 9.436746e-32, 
    9.436755e-32, 9.436715e-32, 9.436703e-32, 9.436646e-32, 9.436669e-32, 
    9.436633e-32, 9.436666e-32, 9.43666e-32, 9.436632e-32, 9.436664e-32, 
    9.436593e-32, 9.436641e-32, 9.436552e-32, 9.4366e-32, 9.436549e-32, 
    9.436558e-32, 9.436543e-32, 9.436529e-32, 9.436512e-32, 9.43648e-32, 
    9.436488e-32, 9.436461e-32, 9.436733e-32, 9.436716e-32, 9.436718e-32, 
    9.436701e-32, 9.436688e-32, 9.436661e-32, 9.436617e-32, 9.436634e-32, 
    9.436603e-32, 9.436597e-32, 9.436643e-32, 9.436615e-32, 9.436706e-32, 
    9.436691e-32, 9.4367e-32, 9.436732e-32, 9.436629e-32, 9.436682e-32, 
    9.436585e-32, 9.436614e-32, 9.436531e-32, 9.436572e-32, 9.436491e-32, 
    9.436457e-32, 9.436425e-32, 9.436387e-32, 9.436708e-32, 9.436719e-32, 
    9.436699e-32, 9.436671e-32, 9.436646e-32, 9.436612e-32, 9.436608e-32, 
    9.436602e-32, 9.436586e-32, 9.436572e-32, 9.4366e-32, 9.436568e-32, 
    9.436688e-32, 9.436625e-32, 9.436723e-32, 9.436693e-32, 9.436673e-32, 
    9.436682e-32, 9.436635e-32, 9.436624e-32, 9.436579e-32, 9.436603e-32, 
    9.436465e-32, 9.436526e-32, 9.436358e-32, 9.436406e-32, 9.436723e-32, 
    9.436708e-32, 9.436656e-32, 9.436681e-32, 9.436609e-32, 9.436592e-32, 
    9.436578e-32, 9.43656e-32, 9.436558e-32, 9.436548e-32, 9.436565e-32, 
    9.436548e-32, 9.436612e-32, 9.436584e-32, 9.436662e-32, 9.436642e-32, 
    9.436651e-32, 9.436661e-32, 9.436631e-32, 9.436599e-32, 9.436599e-32, 
    9.436589e-32, 9.436561e-32, 9.436609e-32, 9.436458e-32, 9.436551e-32, 
    9.436691e-32, 9.436662e-32, 9.436658e-32, 9.436669e-32, 9.436594e-32, 
    9.436621e-32, 9.436548e-32, 9.436568e-32, 9.436535e-32, 9.436551e-32, 
    9.436554e-32, 9.436574e-32, 9.436587e-32, 9.43662e-32, 9.436647e-32, 
    9.436668e-32, 9.436663e-32, 9.43664e-32, 9.436598e-32, 9.436558e-32, 
    9.436567e-32, 9.436538e-32, 9.436615e-32, 9.436582e-32, 9.436595e-32, 
    9.436562e-32, 9.436634e-32, 9.436573e-32, 9.436649e-32, 9.436643e-32, 
    9.436622e-32, 9.43658e-32, 9.436571e-32, 9.436561e-32, 9.436567e-32, 
    9.436597e-32, 9.436602e-32, 9.436622e-32, 9.436628e-32, 9.436644e-32, 
    9.436658e-32, 9.436645e-32, 9.436633e-32, 9.436597e-32, 9.436564e-32, 
    9.436529e-32, 9.43652e-32, 9.436479e-32, 9.436512e-32, 9.436457e-32, 
    9.436504e-32, 9.436423e-32, 9.436569e-32, 9.436506e-32, 9.436621e-32, 
    9.436609e-32, 9.436586e-32, 9.436535e-32, 9.436562e-32, 9.43653e-32, 
    9.436602e-32, 9.436639e-32, 9.436649e-32, 9.436666e-32, 9.436648e-32, 
    9.43665e-32, 9.436632e-32, 9.436638e-32, 9.436595e-32, 9.436618e-32, 
    9.436554e-32, 9.43653e-32, 9.436464e-32, 9.436423e-32, 9.436382e-32, 
    9.436364e-32, 9.436358e-32, 9.436356e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.552066e-14, 4.564366e-14, 4.561977e-14, 4.571889e-14, 4.566393e-14, 
    4.57288e-14, 4.554562e-14, 4.564853e-14, 4.558285e-14, 4.553176e-14, 
    4.591094e-14, 4.572331e-14, 4.610567e-14, 4.598623e-14, 4.628609e-14, 
    4.608707e-14, 4.632618e-14, 4.628039e-14, 4.641824e-14, 4.637876e-14, 
    4.65548e-14, 4.643645e-14, 4.6646e-14, 4.652657e-14, 4.654525e-14, 
    4.643253e-14, 4.576113e-14, 4.588759e-14, 4.575363e-14, 4.577167e-14, 
    4.576358e-14, 4.566505e-14, 4.561534e-14, 4.551127e-14, 4.553018e-14, 
    4.560663e-14, 4.577979e-14, 4.572106e-14, 4.586908e-14, 4.586574e-14, 
    4.603028e-14, 4.595612e-14, 4.623233e-14, 4.615391e-14, 4.638041e-14, 
    4.632349e-14, 4.637773e-14, 4.636129e-14, 4.637795e-14, 4.629445e-14, 
    4.633023e-14, 4.625674e-14, 4.597001e-14, 4.605434e-14, 4.58026e-14, 
    4.565091e-14, 4.555013e-14, 4.547854e-14, 4.548866e-14, 4.550795e-14, 
    4.560707e-14, 4.570022e-14, 4.577114e-14, 4.581856e-14, 4.586526e-14, 
    4.60064e-14, 4.608112e-14, 4.624816e-14, 4.621807e-14, 4.626907e-14, 
    4.631783e-14, 4.639958e-14, 4.638613e-14, 4.642213e-14, 4.626775e-14, 
    4.637036e-14, 4.620092e-14, 4.624728e-14, 4.587783e-14, 4.573691e-14, 
    4.567685e-14, 4.562436e-14, 4.549644e-14, 4.558479e-14, 4.554997e-14, 
    4.563282e-14, 4.568541e-14, 4.565941e-14, 4.581985e-14, 4.57575e-14, 
    4.608554e-14, 4.594436e-14, 4.631214e-14, 4.622425e-14, 4.63332e-14, 
    4.627762e-14, 4.637282e-14, 4.628715e-14, 4.643553e-14, 4.64678e-14, 
    4.644574e-14, 4.653047e-14, 4.62824e-14, 4.637772e-14, 4.565867e-14, 
    4.566291e-14, 4.568268e-14, 4.559575e-14, 4.559044e-14, 4.551075e-14, 
    4.558167e-14, 4.561185e-14, 4.568847e-14, 4.573374e-14, 4.577677e-14, 
    4.587133e-14, 4.597681e-14, 4.612418e-14, 4.622995e-14, 4.630079e-14, 
    4.625736e-14, 4.62957e-14, 4.625284e-14, 4.623275e-14, 4.64557e-14, 
    4.633056e-14, 4.651829e-14, 4.650792e-14, 4.642298e-14, 4.650908e-14, 
    4.566589e-14, 4.564148e-14, 4.555665e-14, 4.562304e-14, 4.550207e-14, 
    4.556979e-14, 4.56087e-14, 4.575877e-14, 4.579175e-14, 4.582228e-14, 
    4.588259e-14, 4.595992e-14, 4.609543e-14, 4.621323e-14, 4.632067e-14, 
    4.63128e-14, 4.631557e-14, 4.633955e-14, 4.628013e-14, 4.63493e-14, 
    4.636089e-14, 4.633056e-14, 4.650653e-14, 4.645629e-14, 4.65077e-14, 
    4.647499e-14, 4.564942e-14, 4.56905e-14, 4.56683e-14, 4.571002e-14, 
    4.568062e-14, 4.581127e-14, 4.585042e-14, 4.603343e-14, 4.595839e-14, 
    4.607783e-14, 4.597053e-14, 4.598955e-14, 4.608167e-14, 4.597635e-14, 
    4.620671e-14, 4.605054e-14, 4.634048e-14, 4.618466e-14, 4.635023e-14, 
    4.63202e-14, 4.636993e-14, 4.641442e-14, 4.647041e-14, 4.657358e-14, 
    4.65497e-14, 4.663594e-14, 4.575171e-14, 4.580492e-14, 4.580026e-14, 
    4.585594e-14, 4.589709e-14, 4.598627e-14, 4.612912e-14, 4.607543e-14, 
    4.617401e-14, 4.619378e-14, 4.604403e-14, 4.613597e-14, 4.584054e-14, 
    4.58883e-14, 4.585988e-14, 4.575589e-14, 4.608778e-14, 4.591756e-14, 
    4.623169e-14, 4.613964e-14, 4.640808e-14, 4.627464e-14, 4.653655e-14, 
    4.664825e-14, 4.675338e-14, 4.687596e-14, 4.583398e-14, 4.579783e-14, 
    4.586257e-14, 4.595203e-14, 4.603503e-14, 4.614525e-14, 4.615654e-14, 
    4.617716e-14, 4.62306e-14, 4.62755e-14, 4.618366e-14, 4.628676e-14, 
    4.589932e-14, 4.610255e-14, 4.578414e-14, 4.588009e-14, 4.594676e-14, 
    4.591754e-14, 4.606931e-14, 4.610503e-14, 4.62501e-14, 4.617514e-14, 
    4.662067e-14, 4.642379e-14, 4.696928e-14, 4.681712e-14, 4.578519e-14, 
    4.583386e-14, 4.600306e-14, 4.592259e-14, 4.615262e-14, 4.620915e-14, 
    4.625511e-14, 4.63138e-14, 4.632015e-14, 4.63549e-14, 4.629795e-14, 
    4.635267e-14, 4.614549e-14, 4.623812e-14, 4.598376e-14, 4.604571e-14, 
    4.601723e-14, 4.598595e-14, 4.608244e-14, 4.61851e-14, 4.618733e-14, 
    4.622022e-14, 4.631279e-14, 4.615355e-14, 4.664598e-14, 4.634207e-14, 
    4.588691e-14, 4.598051e-14, 4.599391e-14, 4.595766e-14, 4.620349e-14, 
    4.611448e-14, 4.635406e-14, 4.628937e-14, 4.639536e-14, 4.63427e-14, 
    4.633495e-14, 4.626728e-14, 4.622513e-14, 4.611855e-14, 4.603177e-14, 
    4.596293e-14, 4.597894e-14, 4.605455e-14, 4.619139e-14, 4.632071e-14, 
    4.629239e-14, 4.638731e-14, 4.613596e-14, 4.62414e-14, 4.620065e-14, 
    4.630689e-14, 4.6074e-14, 4.627223e-14, 4.602326e-14, 4.604512e-14, 
    4.611271e-14, 4.624852e-14, 4.627861e-14, 4.631065e-14, 4.629089e-14, 
    4.619487e-14, 4.617915e-14, 4.611107e-14, 4.609225e-14, 4.604036e-14, 
    4.599737e-14, 4.603664e-14, 4.607787e-14, 4.619492e-14, 4.630029e-14, 
    4.641505e-14, 4.644313e-14, 4.657694e-14, 4.646798e-14, 4.664766e-14, 
    4.649483e-14, 4.675928e-14, 4.628377e-14, 4.649042e-14, 4.61158e-14, 
    4.615623e-14, 4.622927e-14, 4.639671e-14, 4.630639e-14, 4.641203e-14, 
    4.617853e-14, 4.605714e-14, 4.602576e-14, 4.596711e-14, 4.60271e-14, 
    4.602222e-14, 4.60796e-14, 4.606117e-14, 4.619881e-14, 4.61249e-14, 
    4.633475e-14, 4.641121e-14, 4.662689e-14, 4.675886e-14, 4.689309e-14, 
    4.695227e-14, 4.697028e-14, 4.697781e-14 ;

 LITR1N_vr =
  5.557623e-05, 5.557602e-05, 5.557606e-05, 5.557588e-05, 5.557598e-05, 
    5.557587e-05, 5.557619e-05, 5.557601e-05, 5.557612e-05, 5.557621e-05, 
    5.557555e-05, 5.557587e-05, 5.557521e-05, 5.557542e-05, 5.557489e-05, 
    5.557524e-05, 5.557482e-05, 5.55749e-05, 5.557466e-05, 5.557473e-05, 
    5.557442e-05, 5.557463e-05, 5.557426e-05, 5.557447e-05, 5.557444e-05, 
    5.557463e-05, 5.557581e-05, 5.557559e-05, 5.557582e-05, 5.557579e-05, 
    5.557581e-05, 5.557598e-05, 5.557606e-05, 5.557625e-05, 5.557621e-05, 
    5.557608e-05, 5.557578e-05, 5.557588e-05, 5.557562e-05, 5.557563e-05, 
    5.557534e-05, 5.557547e-05, 5.557499e-05, 5.557512e-05, 5.557473e-05, 
    5.557483e-05, 5.557473e-05, 5.557476e-05, 5.557473e-05, 5.557488e-05, 
    5.557482e-05, 5.557494e-05, 5.557545e-05, 5.55753e-05, 5.557574e-05, 
    5.5576e-05, 5.557618e-05, 5.55763e-05, 5.557629e-05, 5.557625e-05, 
    5.557608e-05, 5.557591e-05, 5.557579e-05, 5.557571e-05, 5.557563e-05, 
    5.557538e-05, 5.557525e-05, 5.557496e-05, 5.557501e-05, 5.557492e-05, 
    5.557484e-05, 5.557469e-05, 5.557472e-05, 5.557465e-05, 5.557492e-05, 
    5.557474e-05, 5.557504e-05, 5.557496e-05, 5.557561e-05, 5.557585e-05, 
    5.557596e-05, 5.557605e-05, 5.557627e-05, 5.557612e-05, 5.557618e-05, 
    5.557603e-05, 5.557594e-05, 5.557599e-05, 5.557571e-05, 5.557582e-05, 
    5.557524e-05, 5.557549e-05, 5.557484e-05, 5.5575e-05, 5.557481e-05, 
    5.557491e-05, 5.557474e-05, 5.557489e-05, 5.557463e-05, 5.557458e-05, 
    5.557461e-05, 5.557446e-05, 5.55749e-05, 5.557473e-05, 5.557599e-05, 
    5.557598e-05, 5.557595e-05, 5.55761e-05, 5.557611e-05, 5.557625e-05, 
    5.557612e-05, 5.557607e-05, 5.557594e-05, 5.557586e-05, 5.557578e-05, 
    5.557562e-05, 5.557543e-05, 5.557518e-05, 5.557499e-05, 5.557487e-05, 
    5.557494e-05, 5.557487e-05, 5.557495e-05, 5.557498e-05, 5.557459e-05, 
    5.557481e-05, 5.557448e-05, 5.55745e-05, 5.557465e-05, 5.55745e-05, 
    5.557598e-05, 5.557602e-05, 5.557617e-05, 5.557605e-05, 5.557626e-05, 
    5.557614e-05, 5.557607e-05, 5.557581e-05, 5.557575e-05, 5.55757e-05, 
    5.55756e-05, 5.557546e-05, 5.557522e-05, 5.557502e-05, 5.557483e-05, 
    5.557484e-05, 5.557484e-05, 5.55748e-05, 5.55749e-05, 5.557478e-05, 
    5.557476e-05, 5.557481e-05, 5.557451e-05, 5.557459e-05, 5.55745e-05, 
    5.557456e-05, 5.557601e-05, 5.557593e-05, 5.557597e-05, 5.55759e-05, 
    5.557595e-05, 5.557572e-05, 5.557565e-05, 5.557533e-05, 5.557546e-05, 
    5.557526e-05, 5.557545e-05, 5.557541e-05, 5.557525e-05, 5.557543e-05, 
    5.557503e-05, 5.55753e-05, 5.55748e-05, 5.557507e-05, 5.557478e-05, 
    5.557483e-05, 5.557475e-05, 5.557467e-05, 5.557457e-05, 5.557439e-05, 
    5.557443e-05, 5.557428e-05, 5.557583e-05, 5.557573e-05, 5.557574e-05, 
    5.557565e-05, 5.557557e-05, 5.557542e-05, 5.557516e-05, 5.557526e-05, 
    5.557509e-05, 5.557505e-05, 5.557531e-05, 5.557515e-05, 5.557567e-05, 
    5.557559e-05, 5.557564e-05, 5.557582e-05, 5.557524e-05, 5.557554e-05, 
    5.557499e-05, 5.557515e-05, 5.557468e-05, 5.557491e-05, 5.557445e-05, 
    5.557426e-05, 5.557407e-05, 5.557386e-05, 5.557568e-05, 5.557574e-05, 
    5.557563e-05, 5.557547e-05, 5.557533e-05, 5.557514e-05, 5.557512e-05, 
    5.557508e-05, 5.557499e-05, 5.557491e-05, 5.557507e-05, 5.557489e-05, 
    5.557557e-05, 5.557521e-05, 5.557577e-05, 5.55756e-05, 5.557549e-05, 
    5.557554e-05, 5.557527e-05, 5.557521e-05, 5.557495e-05, 5.557508e-05, 
    5.557431e-05, 5.557465e-05, 5.55737e-05, 5.557396e-05, 5.557577e-05, 
    5.557568e-05, 5.557539e-05, 5.557553e-05, 5.557512e-05, 5.557503e-05, 
    5.557495e-05, 5.557484e-05, 5.557483e-05, 5.557477e-05, 5.557487e-05, 
    5.557478e-05, 5.557514e-05, 5.557498e-05, 5.557542e-05, 5.557531e-05, 
    5.557536e-05, 5.557542e-05, 5.557525e-05, 5.557507e-05, 5.557506e-05, 
    5.557501e-05, 5.557484e-05, 5.557512e-05, 5.557426e-05, 5.557479e-05, 
    5.557559e-05, 5.557543e-05, 5.55754e-05, 5.557547e-05, 5.557504e-05, 
    5.557519e-05, 5.557477e-05, 5.557488e-05, 5.55747e-05, 5.557479e-05, 
    5.55748e-05, 5.557492e-05, 5.5575e-05, 5.557518e-05, 5.557534e-05, 
    5.557546e-05, 5.557543e-05, 5.55753e-05, 5.557506e-05, 5.557483e-05, 
    5.557488e-05, 5.557471e-05, 5.557515e-05, 5.557497e-05, 5.557504e-05, 
    5.557486e-05, 5.557526e-05, 5.557492e-05, 5.557535e-05, 5.557531e-05, 
    5.557519e-05, 5.557496e-05, 5.55749e-05, 5.557485e-05, 5.557488e-05, 
    5.557505e-05, 5.557508e-05, 5.55752e-05, 5.557523e-05, 5.557532e-05, 
    5.55754e-05, 5.557533e-05, 5.557526e-05, 5.557505e-05, 5.557487e-05, 
    5.557467e-05, 5.557462e-05, 5.557438e-05, 5.557457e-05, 5.557426e-05, 
    5.557453e-05, 5.557406e-05, 5.55749e-05, 5.557454e-05, 5.557519e-05, 
    5.557512e-05, 5.557499e-05, 5.55747e-05, 5.557486e-05, 5.557467e-05, 
    5.557508e-05, 5.557529e-05, 5.557535e-05, 5.557545e-05, 5.557534e-05, 
    5.557535e-05, 5.557525e-05, 5.557528e-05, 5.557504e-05, 5.557517e-05, 
    5.55748e-05, 5.557467e-05, 5.55743e-05, 5.557407e-05, 5.557383e-05, 
    5.557373e-05, 5.55737e-05, 5.557368e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  7.888883e-13, 7.910201e-13, 7.90606e-13, 7.923238e-13, 7.913713e-13, 
    7.924956e-13, 7.89321e-13, 7.911044e-13, 7.899663e-13, 7.890807e-13, 
    7.956522e-13, 7.924004e-13, 7.990269e-13, 7.969568e-13, 8.021535e-13, 
    7.987045e-13, 8.028483e-13, 8.020548e-13, 8.044437e-13, 8.037597e-13, 
    8.068105e-13, 8.047593e-13, 8.083909e-13, 8.063212e-13, 8.066449e-13, 
    8.046915e-13, 7.930559e-13, 7.952474e-13, 7.929258e-13, 7.932385e-13, 
    7.930984e-13, 7.913908e-13, 7.905293e-13, 7.887257e-13, 7.890534e-13, 
    7.903782e-13, 7.933791e-13, 7.923614e-13, 7.949266e-13, 7.948688e-13, 
    7.977203e-13, 7.964351e-13, 8.01222e-13, 7.998628e-13, 8.037882e-13, 
    8.028017e-13, 8.037418e-13, 8.034569e-13, 8.037455e-13, 8.022985e-13, 
    8.029186e-13, 8.016449e-13, 7.966757e-13, 7.981373e-13, 7.937746e-13, 
    7.911456e-13, 7.893991e-13, 7.881584e-13, 7.883339e-13, 7.886682e-13, 
    7.90386e-13, 7.920003e-13, 7.932294e-13, 7.940511e-13, 7.948604e-13, 
    7.973065e-13, 7.986014e-13, 8.014963e-13, 8.009748e-13, 8.018587e-13, 
    8.027036e-13, 8.041204e-13, 8.038873e-13, 8.045111e-13, 8.018358e-13, 
    8.036141e-13, 8.006775e-13, 8.014811e-13, 7.950782e-13, 7.926361e-13, 
    7.915954e-13, 7.906856e-13, 7.884687e-13, 7.899997e-13, 7.893963e-13, 
    7.908321e-13, 7.917436e-13, 7.91293e-13, 7.940735e-13, 7.929929e-13, 
    7.986781e-13, 7.962314e-13, 8.026051e-13, 8.010819e-13, 8.0297e-13, 
    8.020069e-13, 8.036567e-13, 8.02172e-13, 8.047434e-13, 8.053027e-13, 
    8.049205e-13, 8.063888e-13, 8.020896e-13, 8.037416e-13, 7.912802e-13, 
    7.913537e-13, 7.916964e-13, 7.901897e-13, 7.900977e-13, 7.887166e-13, 
    7.899457e-13, 7.904687e-13, 7.917966e-13, 7.925812e-13, 7.933269e-13, 
    7.949655e-13, 7.967936e-13, 7.993476e-13, 8.011806e-13, 8.024083e-13, 
    8.016557e-13, 8.023202e-13, 8.015773e-13, 8.012292e-13, 8.05093e-13, 
    8.029242e-13, 8.061777e-13, 8.059979e-13, 8.045259e-13, 8.060182e-13, 
    7.914054e-13, 7.909823e-13, 7.895122e-13, 7.906628e-13, 7.885663e-13, 
    7.897398e-13, 7.904141e-13, 7.93015e-13, 7.935866e-13, 7.941156e-13, 
    7.951608e-13, 7.965009e-13, 7.988494e-13, 8.008908e-13, 8.027528e-13, 
    8.026165e-13, 8.026645e-13, 8.0308e-13, 8.020503e-13, 8.03249e-13, 
    8.034499e-13, 8.029242e-13, 8.059738e-13, 8.051032e-13, 8.059941e-13, 
    8.054273e-13, 7.911199e-13, 7.918317e-13, 7.914471e-13, 7.921702e-13, 
    7.916606e-13, 7.939249e-13, 7.946032e-13, 7.977749e-13, 7.964744e-13, 
    7.985443e-13, 7.966849e-13, 7.970144e-13, 7.986109e-13, 7.967856e-13, 
    8.007779e-13, 7.980714e-13, 8.030961e-13, 8.003957e-13, 8.032652e-13, 
    8.027448e-13, 8.036065e-13, 8.043777e-13, 8.053479e-13, 8.071358e-13, 
    8.06722e-13, 8.082167e-13, 7.928926e-13, 7.938148e-13, 7.93734e-13, 
    7.946989e-13, 7.954122e-13, 7.969577e-13, 7.994333e-13, 7.985029e-13, 
    8.002111e-13, 8.005537e-13, 7.979586e-13, 7.99552e-13, 7.94432e-13, 
    7.952597e-13, 7.947672e-13, 7.929651e-13, 7.987168e-13, 7.957669e-13, 
    8.012108e-13, 7.996156e-13, 8.042677e-13, 8.019551e-13, 8.064941e-13, 
    8.084299e-13, 8.102518e-13, 8.123763e-13, 7.943183e-13, 7.936919e-13, 
    7.948138e-13, 7.963641e-13, 7.978027e-13, 7.997128e-13, 7.999084e-13, 
    8.002659e-13, 8.01192e-13, 8.019701e-13, 8.003785e-13, 8.021652e-13, 
    7.954508e-13, 7.989728e-13, 7.934546e-13, 7.951173e-13, 7.96273e-13, 
    7.957666e-13, 7.983966e-13, 7.990158e-13, 8.015298e-13, 8.002309e-13, 
    8.07952e-13, 8.045399e-13, 8.139935e-13, 8.113565e-13, 7.934729e-13, 
    7.943164e-13, 7.972486e-13, 7.958541e-13, 7.998405e-13, 8.008203e-13, 
    8.016167e-13, 8.026338e-13, 8.027439e-13, 8.033462e-13, 8.02359e-13, 
    8.033073e-13, 7.997169e-13, 8.013223e-13, 7.969141e-13, 7.979878e-13, 
    7.974941e-13, 7.969521e-13, 7.986242e-13, 8.004034e-13, 8.004421e-13, 
    8.010121e-13, 8.026163e-13, 7.998567e-13, 8.083906e-13, 8.031238e-13, 
    7.952357e-13, 7.968577e-13, 7.970901e-13, 7.964619e-13, 8.007221e-13, 
    7.991795e-13, 8.033316e-13, 8.022105e-13, 8.040472e-13, 8.031347e-13, 
    8.030004e-13, 8.018277e-13, 8.010971e-13, 7.992501e-13, 7.977461e-13, 
    7.965531e-13, 7.968306e-13, 7.98141e-13, 8.005124e-13, 8.027535e-13, 
    8.022628e-13, 8.039077e-13, 7.995517e-13, 8.013791e-13, 8.006728e-13, 
    8.025141e-13, 7.98478e-13, 8.019134e-13, 7.975986e-13, 7.979775e-13, 
    7.991488e-13, 8.015025e-13, 8.02024e-13, 8.025792e-13, 8.022367e-13, 
    8.005727e-13, 8.003002e-13, 7.991205e-13, 7.987944e-13, 7.978951e-13, 
    7.971499e-13, 7.978306e-13, 7.98545e-13, 8.005736e-13, 8.023996e-13, 
    8.043885e-13, 8.048752e-13, 8.07194e-13, 8.053057e-13, 8.084197e-13, 
    8.057712e-13, 8.103542e-13, 8.021134e-13, 8.056946e-13, 7.992023e-13, 
    7.99903e-13, 8.01169e-13, 8.040707e-13, 8.025055e-13, 8.043362e-13, 
    8.002896e-13, 7.981858e-13, 7.97642e-13, 7.966255e-13, 7.976652e-13, 
    7.975807e-13, 7.985751e-13, 7.982556e-13, 8.00641e-13, 7.9936e-13, 
    8.029968e-13, 8.043219e-13, 8.080598e-13, 8.10347e-13, 8.126732e-13, 
    8.136988e-13, 8.140109e-13, 8.141413e-13 ;

 LITR2C =
  1.939604e-05, 1.939602e-05, 1.939602e-05, 1.9396e-05, 1.939601e-05, 
    1.9396e-05, 1.939603e-05, 1.939601e-05, 1.939603e-05, 1.939603e-05, 
    1.939597e-05, 1.9396e-05, 1.939594e-05, 1.939596e-05, 1.939591e-05, 
    1.939594e-05, 1.939591e-05, 1.939591e-05, 1.939589e-05, 1.93959e-05, 
    1.939587e-05, 1.939589e-05, 1.939585e-05, 1.939587e-05, 1.939587e-05, 
    1.939589e-05, 1.9396e-05, 1.939598e-05, 1.9396e-05, 1.939599e-05, 
    1.9396e-05, 1.939601e-05, 1.939602e-05, 1.939604e-05, 1.939603e-05, 
    1.939602e-05, 1.939599e-05, 1.9396e-05, 1.939598e-05, 1.939598e-05, 
    1.939595e-05, 1.939597e-05, 1.939592e-05, 1.939593e-05, 1.93959e-05, 
    1.939591e-05, 1.93959e-05, 1.93959e-05, 1.93959e-05, 1.939591e-05, 
    1.939591e-05, 1.939592e-05, 1.939596e-05, 1.939595e-05, 1.939599e-05, 
    1.939601e-05, 1.939603e-05, 1.939604e-05, 1.939604e-05, 1.939604e-05, 
    1.939602e-05, 1.939601e-05, 1.9396e-05, 1.939599e-05, 1.939598e-05, 
    1.939596e-05, 1.939595e-05, 1.939592e-05, 1.939592e-05, 1.939591e-05, 
    1.939591e-05, 1.939589e-05, 1.93959e-05, 1.939589e-05, 1.939591e-05, 
    1.93959e-05, 1.939593e-05, 1.939592e-05, 1.939598e-05, 1.9396e-05, 
    1.939601e-05, 1.939602e-05, 1.939604e-05, 1.939603e-05, 1.939603e-05, 
    1.939602e-05, 1.939601e-05, 1.939601e-05, 1.939599e-05, 1.9396e-05, 
    1.939595e-05, 1.939597e-05, 1.939591e-05, 1.939592e-05, 1.939591e-05, 
    1.939591e-05, 1.93959e-05, 1.939591e-05, 1.939589e-05, 1.939588e-05, 
    1.939589e-05, 1.939587e-05, 1.939591e-05, 1.93959e-05, 1.939601e-05, 
    1.939601e-05, 1.939601e-05, 1.939602e-05, 1.939603e-05, 1.939604e-05, 
    1.939603e-05, 1.939602e-05, 1.939601e-05, 1.9396e-05, 1.939599e-05, 
    1.939598e-05, 1.939596e-05, 1.939594e-05, 1.939592e-05, 1.939591e-05, 
    1.939592e-05, 1.939591e-05, 1.939592e-05, 1.939592e-05, 1.939589e-05, 
    1.939591e-05, 1.939587e-05, 1.939588e-05, 1.939589e-05, 1.939588e-05, 
    1.939601e-05, 1.939602e-05, 1.939603e-05, 1.939602e-05, 1.939604e-05, 
    1.939603e-05, 1.939602e-05, 1.9396e-05, 1.939599e-05, 1.939599e-05, 
    1.939598e-05, 1.939597e-05, 1.939594e-05, 1.939592e-05, 1.939591e-05, 
    1.939591e-05, 1.939591e-05, 1.93959e-05, 1.939591e-05, 1.93959e-05, 
    1.93959e-05, 1.939591e-05, 1.939588e-05, 1.939589e-05, 1.939588e-05, 
    1.939588e-05, 1.939601e-05, 1.939601e-05, 1.939601e-05, 1.939601e-05, 
    1.939601e-05, 1.939599e-05, 1.939598e-05, 1.939595e-05, 1.939597e-05, 
    1.939595e-05, 1.939596e-05, 1.939596e-05, 1.939595e-05, 1.939596e-05, 
    1.939593e-05, 1.939595e-05, 1.93959e-05, 1.939593e-05, 1.93959e-05, 
    1.939591e-05, 1.93959e-05, 1.939589e-05, 1.939588e-05, 1.939587e-05, 
    1.939587e-05, 1.939586e-05, 1.9396e-05, 1.939599e-05, 1.939599e-05, 
    1.939598e-05, 1.939597e-05, 1.939596e-05, 1.939594e-05, 1.939595e-05, 
    1.939593e-05, 1.939593e-05, 1.939595e-05, 1.939594e-05, 1.939598e-05, 
    1.939598e-05, 1.939598e-05, 1.9396e-05, 1.939594e-05, 1.939597e-05, 
    1.939592e-05, 1.939594e-05, 1.939589e-05, 1.939591e-05, 1.939587e-05, 
    1.939585e-05, 1.939584e-05, 1.939582e-05, 1.939599e-05, 1.939599e-05, 
    1.939598e-05, 1.939597e-05, 1.939595e-05, 1.939593e-05, 1.939593e-05, 
    1.939593e-05, 1.939592e-05, 1.939591e-05, 1.939593e-05, 1.939591e-05, 
    1.939597e-05, 1.939594e-05, 1.939599e-05, 1.939598e-05, 1.939597e-05, 
    1.939597e-05, 1.939595e-05, 1.939594e-05, 1.939592e-05, 1.939593e-05, 
    1.939586e-05, 1.939589e-05, 1.93958e-05, 1.939583e-05, 1.939599e-05, 
    1.939599e-05, 1.939596e-05, 1.939597e-05, 1.939593e-05, 1.939593e-05, 
    1.939592e-05, 1.939591e-05, 1.939591e-05, 1.93959e-05, 1.939591e-05, 
    1.93959e-05, 1.939593e-05, 1.939592e-05, 1.939596e-05, 1.939595e-05, 
    1.939596e-05, 1.939596e-05, 1.939595e-05, 1.939593e-05, 1.939593e-05, 
    1.939592e-05, 1.939591e-05, 1.939593e-05, 1.939585e-05, 1.93959e-05, 
    1.939598e-05, 1.939596e-05, 1.939596e-05, 1.939597e-05, 1.939593e-05, 
    1.939594e-05, 1.93959e-05, 1.939591e-05, 1.939589e-05, 1.93959e-05, 
    1.93959e-05, 1.939591e-05, 1.939592e-05, 1.939594e-05, 1.939595e-05, 
    1.939596e-05, 1.939596e-05, 1.939595e-05, 1.939593e-05, 1.939591e-05, 
    1.939591e-05, 1.93959e-05, 1.939594e-05, 1.939592e-05, 1.939593e-05, 
    1.939591e-05, 1.939595e-05, 1.939591e-05, 1.939595e-05, 1.939595e-05, 
    1.939594e-05, 1.939592e-05, 1.939591e-05, 1.939591e-05, 1.939591e-05, 
    1.939593e-05, 1.939593e-05, 1.939594e-05, 1.939594e-05, 1.939595e-05, 
    1.939596e-05, 1.939595e-05, 1.939595e-05, 1.939593e-05, 1.939591e-05, 
    1.939589e-05, 1.939589e-05, 1.939587e-05, 1.939588e-05, 1.939585e-05, 
    1.939588e-05, 1.939584e-05, 1.939591e-05, 1.939588e-05, 1.939594e-05, 
    1.939593e-05, 1.939592e-05, 1.939589e-05, 1.939591e-05, 1.939589e-05, 
    1.939593e-05, 1.939595e-05, 1.939595e-05, 1.939596e-05, 1.939595e-05, 
    1.939595e-05, 1.939595e-05, 1.939595e-05, 1.939593e-05, 1.939594e-05, 
    1.939591e-05, 1.939589e-05, 1.939586e-05, 1.939584e-05, 1.939581e-05, 
    1.939581e-05, 1.93958e-05, 1.93958e-05 ;

 LITR2C_TO_SOIL1C =
  1.201324e-13, 1.204574e-13, 1.203942e-13, 1.206561e-13, 1.205109e-13, 
    1.206823e-13, 1.201984e-13, 1.204702e-13, 1.202967e-13, 1.201617e-13, 
    1.211635e-13, 1.206678e-13, 1.216779e-13, 1.213624e-13, 1.221545e-13, 
    1.216288e-13, 1.222605e-13, 1.221395e-13, 1.225037e-13, 1.223994e-13, 
    1.228644e-13, 1.225518e-13, 1.231054e-13, 1.227899e-13, 1.228392e-13, 
    1.225414e-13, 1.207677e-13, 1.211018e-13, 1.207479e-13, 1.207955e-13, 
    1.207742e-13, 1.205139e-13, 1.203825e-13, 1.201076e-13, 1.201576e-13, 
    1.203595e-13, 1.20817e-13, 1.206618e-13, 1.210529e-13, 1.21044e-13, 
    1.214787e-13, 1.212828e-13, 1.220125e-13, 1.218053e-13, 1.224037e-13, 
    1.222533e-13, 1.223967e-13, 1.223532e-13, 1.223972e-13, 1.221766e-13, 
    1.222712e-13, 1.22077e-13, 1.213195e-13, 1.215423e-13, 1.208773e-13, 
    1.204765e-13, 1.202103e-13, 1.200211e-13, 1.200479e-13, 1.200988e-13, 
    1.203607e-13, 1.206068e-13, 1.207941e-13, 1.209194e-13, 1.210428e-13, 
    1.214157e-13, 1.21613e-13, 1.220544e-13, 1.219748e-13, 1.221096e-13, 
    1.222384e-13, 1.224544e-13, 1.224188e-13, 1.225139e-13, 1.221061e-13, 
    1.223772e-13, 1.219295e-13, 1.22052e-13, 1.21076e-13, 1.207037e-13, 
    1.205451e-13, 1.204064e-13, 1.200684e-13, 1.203018e-13, 1.202098e-13, 
    1.204287e-13, 1.205677e-13, 1.20499e-13, 1.209228e-13, 1.207581e-13, 
    1.216247e-13, 1.212518e-13, 1.222234e-13, 1.219912e-13, 1.22279e-13, 
    1.221322e-13, 1.223837e-13, 1.221574e-13, 1.225494e-13, 1.226346e-13, 
    1.225763e-13, 1.228002e-13, 1.221448e-13, 1.223966e-13, 1.20497e-13, 
    1.205082e-13, 1.205604e-13, 1.203308e-13, 1.203168e-13, 1.201062e-13, 
    1.202936e-13, 1.203733e-13, 1.205757e-13, 1.206953e-13, 1.20809e-13, 
    1.210588e-13, 1.213375e-13, 1.217268e-13, 1.220062e-13, 1.221934e-13, 
    1.220787e-13, 1.221799e-13, 1.220667e-13, 1.220136e-13, 1.226026e-13, 
    1.22272e-13, 1.22768e-13, 1.227406e-13, 1.225162e-13, 1.227437e-13, 
    1.205161e-13, 1.204516e-13, 1.202275e-13, 1.204029e-13, 1.200833e-13, 
    1.202622e-13, 1.20365e-13, 1.207615e-13, 1.208486e-13, 1.209292e-13, 
    1.210886e-13, 1.212928e-13, 1.216509e-13, 1.219621e-13, 1.222459e-13, 
    1.222251e-13, 1.222324e-13, 1.222958e-13, 1.221388e-13, 1.223215e-13, 
    1.223521e-13, 1.22272e-13, 1.227369e-13, 1.226042e-13, 1.2274e-13, 
    1.226536e-13, 1.204726e-13, 1.205811e-13, 1.205224e-13, 1.206327e-13, 
    1.20555e-13, 1.209002e-13, 1.210036e-13, 1.21487e-13, 1.212888e-13, 
    1.216043e-13, 1.213209e-13, 1.213711e-13, 1.216145e-13, 1.213362e-13, 
    1.219448e-13, 1.215322e-13, 1.222982e-13, 1.218866e-13, 1.22324e-13, 
    1.222447e-13, 1.22376e-13, 1.224936e-13, 1.226415e-13, 1.22914e-13, 
    1.22851e-13, 1.230788e-13, 1.207428e-13, 1.208834e-13, 1.208711e-13, 
    1.210182e-13, 1.211269e-13, 1.213625e-13, 1.217399e-13, 1.21598e-13, 
    1.218584e-13, 1.219107e-13, 1.215151e-13, 1.21758e-13, 1.209775e-13, 
    1.211036e-13, 1.210286e-13, 1.207539e-13, 1.216306e-13, 1.21181e-13, 
    1.220108e-13, 1.217677e-13, 1.224768e-13, 1.221243e-13, 1.228162e-13, 
    1.231113e-13, 1.233891e-13, 1.237129e-13, 1.209601e-13, 1.208646e-13, 
    1.210357e-13, 1.21272e-13, 1.214913e-13, 1.217825e-13, 1.218123e-13, 
    1.218668e-13, 1.22008e-13, 1.221266e-13, 1.218839e-13, 1.221563e-13, 
    1.211328e-13, 1.216697e-13, 1.208285e-13, 1.210819e-13, 1.212581e-13, 
    1.211809e-13, 1.215818e-13, 1.216762e-13, 1.220595e-13, 1.218615e-13, 
    1.230385e-13, 1.225183e-13, 1.239595e-13, 1.235575e-13, 1.208313e-13, 
    1.209598e-13, 1.214068e-13, 1.211942e-13, 1.218019e-13, 1.219513e-13, 
    1.220727e-13, 1.222277e-13, 1.222445e-13, 1.223363e-13, 1.221859e-13, 
    1.223304e-13, 1.217831e-13, 1.220278e-13, 1.213558e-13, 1.215195e-13, 
    1.214443e-13, 1.213616e-13, 1.216165e-13, 1.218878e-13, 1.218937e-13, 
    1.219805e-13, 1.222251e-13, 1.218044e-13, 1.231053e-13, 1.223025e-13, 
    1.211e-13, 1.213472e-13, 1.213827e-13, 1.212869e-13, 1.219363e-13, 
    1.217012e-13, 1.223341e-13, 1.221632e-13, 1.224432e-13, 1.223041e-13, 
    1.222836e-13, 1.221049e-13, 1.219935e-13, 1.217119e-13, 1.214827e-13, 
    1.213008e-13, 1.213431e-13, 1.215429e-13, 1.219044e-13, 1.22246e-13, 
    1.221712e-13, 1.224219e-13, 1.217579e-13, 1.220365e-13, 1.219288e-13, 
    1.222095e-13, 1.215942e-13, 1.221179e-13, 1.214602e-13, 1.215179e-13, 
    1.216965e-13, 1.220553e-13, 1.221348e-13, 1.222194e-13, 1.221672e-13, 
    1.219135e-13, 1.21872e-13, 1.216922e-13, 1.216425e-13, 1.215054e-13, 
    1.213918e-13, 1.214955e-13, 1.216045e-13, 1.219137e-13, 1.221921e-13, 
    1.224952e-13, 1.225694e-13, 1.229229e-13, 1.226351e-13, 1.231098e-13, 
    1.22706e-13, 1.234047e-13, 1.221484e-13, 1.226943e-13, 1.217046e-13, 
    1.218115e-13, 1.220044e-13, 1.224468e-13, 1.222082e-13, 1.224873e-13, 
    1.218704e-13, 1.215497e-13, 1.214668e-13, 1.213118e-13, 1.214703e-13, 
    1.214575e-13, 1.21609e-13, 1.215603e-13, 1.21924e-13, 1.217287e-13, 
    1.222831e-13, 1.224851e-13, 1.230549e-13, 1.234036e-13, 1.237582e-13, 
    1.239145e-13, 1.239621e-13, 1.23982e-13 ;

 LITR2C_vr =
  0.001107534, 0.001107533, 0.001107533, 0.001107532, 0.001107532, 
    0.001107532, 0.001107533, 0.001107533, 0.001107533, 0.001107534, 
    0.00110753, 0.001107532, 0.001107528, 0.001107529, 0.001107527, 
    0.001107528, 0.001107526, 0.001107527, 0.001107525, 0.001107526, 
    0.001107524, 0.001107525, 0.001107523, 0.001107524, 0.001107524, 
    0.001107525, 0.001107531, 0.00110753, 0.001107532, 0.001107531, 
    0.001107531, 0.001107532, 0.001107533, 0.001107534, 0.001107534, 
    0.001107533, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.001107529, 0.00110753, 0.001107527, 0.001107528, 0.001107526, 
    0.001107526, 0.001107526, 0.001107526, 0.001107526, 0.001107527, 
    0.001107526, 0.001107527, 0.00110753, 0.001107529, 0.001107531, 
    0.001107533, 0.001107533, 0.001107534, 0.001107534, 0.001107534, 
    0.001107533, 0.001107532, 0.001107531, 0.001107531, 0.001107531, 
    0.001107529, 0.001107529, 0.001107527, 0.001107527, 0.001107527, 
    0.001107526, 0.001107526, 0.001107526, 0.001107525, 0.001107527, 
    0.001107526, 0.001107527, 0.001107527, 0.00110753, 0.001107532, 
    0.001107532, 0.001107533, 0.001107534, 0.001107533, 0.001107533, 
    0.001107533, 0.001107532, 0.001107532, 0.001107531, 0.001107531, 
    0.001107528, 0.00110753, 0.001107526, 0.001107527, 0.001107526, 
    0.001107527, 0.001107526, 0.001107527, 0.001107525, 0.001107525, 
    0.001107525, 0.001107524, 0.001107527, 0.001107526, 0.001107532, 
    0.001107532, 0.001107532, 0.001107533, 0.001107533, 0.001107534, 
    0.001107533, 0.001107533, 0.001107532, 0.001107532, 0.001107531, 
    0.00110753, 0.00110753, 0.001107528, 0.001107527, 0.001107526, 
    0.001107527, 0.001107527, 0.001107527, 0.001107527, 0.001107525, 
    0.001107526, 0.001107524, 0.001107525, 0.001107525, 0.001107525, 
    0.001107532, 0.001107533, 0.001107533, 0.001107533, 0.001107534, 
    0.001107533, 0.001107533, 0.001107531, 0.001107531, 0.001107531, 
    0.00110753, 0.00110753, 0.001107528, 0.001107527, 0.001107526, 
    0.001107526, 0.001107526, 0.001107526, 0.001107527, 0.001107526, 
    0.001107526, 0.001107526, 0.001107525, 0.001107525, 0.001107525, 
    0.001107525, 0.001107533, 0.001107532, 0.001107532, 0.001107532, 
    0.001107532, 0.001107531, 0.001107531, 0.001107529, 0.00110753, 
    0.001107529, 0.00110753, 0.001107529, 0.001107529, 0.00110753, 
    0.001107527, 0.001107529, 0.001107526, 0.001107528, 0.001107526, 
    0.001107526, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107524, 0.001107523, 0.001107532, 0.001107531, 0.001107531, 
    0.001107531, 0.00110753, 0.001107529, 0.001107528, 0.001107529, 
    0.001107528, 0.001107528, 0.001107529, 0.001107528, 0.001107531, 
    0.00110753, 0.001107531, 0.001107532, 0.001107528, 0.00110753, 
    0.001107527, 0.001107528, 0.001107526, 0.001107527, 0.001107524, 
    0.001107523, 0.001107522, 0.001107521, 0.001107531, 0.001107531, 
    0.001107531, 0.00110753, 0.001107529, 0.001107528, 0.001107528, 
    0.001107528, 0.001107527, 0.001107527, 0.001107528, 0.001107527, 
    0.00110753, 0.001107528, 0.001107531, 0.00110753, 0.00110753, 0.00110753, 
    0.001107529, 0.001107528, 0.001107527, 0.001107528, 0.001107524, 
    0.001107525, 0.00110752, 0.001107522, 0.001107531, 0.001107531, 
    0.001107529, 0.00110753, 0.001107528, 0.001107527, 0.001107527, 
    0.001107526, 0.001107526, 0.001107526, 0.001107527, 0.001107526, 
    0.001107528, 0.001107527, 0.00110753, 0.001107529, 0.001107529, 
    0.001107529, 0.001107529, 0.001107528, 0.001107528, 0.001107527, 
    0.001107526, 0.001107528, 0.001107523, 0.001107526, 0.00110753, 
    0.00110753, 0.001107529, 0.00110753, 0.001107527, 0.001107528, 
    0.001107526, 0.001107527, 0.001107526, 0.001107526, 0.001107526, 
    0.001107527, 0.001107527, 0.001107528, 0.001107529, 0.00110753, 
    0.00110753, 0.001107529, 0.001107528, 0.001107526, 0.001107527, 
    0.001107526, 0.001107528, 0.001107527, 0.001107527, 0.001107526, 
    0.001107529, 0.001107527, 0.001107529, 0.001107529, 0.001107528, 
    0.001107527, 0.001107527, 0.001107526, 0.001107527, 0.001107528, 
    0.001107528, 0.001107528, 0.001107528, 0.001107529, 0.001107529, 
    0.001107529, 0.001107529, 0.001107528, 0.001107526, 0.001107525, 
    0.001107525, 0.001107524, 0.001107525, 0.001107523, 0.001107525, 
    0.001107522, 0.001107527, 0.001107525, 0.001107528, 0.001107528, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107528, 
    0.001107529, 0.001107529, 0.00110753, 0.001107529, 0.001107529, 
    0.001107529, 0.001107529, 0.001107528, 0.001107528, 0.001107526, 
    0.001107526, 0.001107524, 0.001107522, 0.001107521, 0.001107521, 
    0.00110752, 0.00110752,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684269e-07, 2.684266e-07, 2.684266e-07, 2.684264e-07, 2.684266e-07, 
    2.684264e-07, 2.684268e-07, 2.684266e-07, 2.684267e-07, 2.684268e-07, 
    2.68426e-07, 2.684264e-07, 2.684256e-07, 2.684259e-07, 2.684252e-07, 
    2.684256e-07, 2.684251e-07, 2.684252e-07, 2.684249e-07, 2.68425e-07, 
    2.684246e-07, 2.684248e-07, 2.684244e-07, 2.684246e-07, 2.684246e-07, 
    2.684249e-07, 2.684263e-07, 2.68426e-07, 2.684264e-07, 2.684263e-07, 
    2.684263e-07, 2.684266e-07, 2.684267e-07, 2.684269e-07, 2.684269e-07, 
    2.684267e-07, 2.684263e-07, 2.684264e-07, 2.684261e-07, 2.684261e-07, 
    2.684257e-07, 2.684259e-07, 2.684253e-07, 2.684255e-07, 2.68425e-07, 
    2.684251e-07, 2.68425e-07, 2.68425e-07, 2.68425e-07, 2.684251e-07, 
    2.684251e-07, 2.684252e-07, 2.684259e-07, 2.684257e-07, 2.684262e-07, 
    2.684266e-07, 2.684268e-07, 2.68427e-07, 2.68427e-07, 2.684269e-07, 
    2.684267e-07, 2.684265e-07, 2.684263e-07, 2.684262e-07, 2.684261e-07, 
    2.684258e-07, 2.684256e-07, 2.684253e-07, 2.684253e-07, 2.684252e-07, 
    2.684251e-07, 2.684249e-07, 2.684249e-07, 2.684249e-07, 2.684252e-07, 
    2.68425e-07, 2.684254e-07, 2.684253e-07, 2.684261e-07, 2.684264e-07, 
    2.684265e-07, 2.684266e-07, 2.684269e-07, 2.684267e-07, 2.684268e-07, 
    2.684266e-07, 2.684265e-07, 2.684266e-07, 2.684262e-07, 2.684264e-07, 
    2.684256e-07, 2.684259e-07, 2.684251e-07, 2.684253e-07, 2.684251e-07, 
    2.684252e-07, 2.68425e-07, 2.684252e-07, 2.684248e-07, 2.684248e-07, 
    2.684248e-07, 2.684246e-07, 2.684252e-07, 2.68425e-07, 2.684266e-07, 
    2.684266e-07, 2.684265e-07, 2.684267e-07, 2.684267e-07, 2.684269e-07, 
    2.684267e-07, 2.684267e-07, 2.684265e-07, 2.684264e-07, 2.684263e-07, 
    2.684261e-07, 2.684259e-07, 2.684255e-07, 2.684253e-07, 2.684251e-07, 
    2.684252e-07, 2.684251e-07, 2.684253e-07, 2.684253e-07, 2.684248e-07, 
    2.684251e-07, 2.684247e-07, 2.684247e-07, 2.684249e-07, 2.684247e-07, 
    2.684266e-07, 2.684266e-07, 2.684268e-07, 2.684266e-07, 2.684269e-07, 
    2.684268e-07, 2.684267e-07, 2.684264e-07, 2.684263e-07, 2.684262e-07, 
    2.684261e-07, 2.684259e-07, 2.684256e-07, 2.684253e-07, 2.684251e-07, 
    2.684251e-07, 2.684251e-07, 2.684251e-07, 2.684252e-07, 2.68425e-07, 
    2.68425e-07, 2.684251e-07, 2.684247e-07, 2.684248e-07, 2.684247e-07, 
    2.684247e-07, 2.684266e-07, 2.684265e-07, 2.684266e-07, 2.684264e-07, 
    2.684265e-07, 2.684262e-07, 2.684261e-07, 2.684257e-07, 2.684259e-07, 
    2.684256e-07, 2.684259e-07, 2.684258e-07, 2.684256e-07, 2.684259e-07, 
    2.684253e-07, 2.684257e-07, 2.684251e-07, 2.684254e-07, 2.68425e-07, 
    2.684251e-07, 2.68425e-07, 2.684249e-07, 2.684248e-07, 2.684245e-07, 
    2.684246e-07, 2.684244e-07, 2.684264e-07, 2.684262e-07, 2.684262e-07, 
    2.684261e-07, 2.68426e-07, 2.684259e-07, 2.684255e-07, 2.684257e-07, 
    2.684254e-07, 2.684254e-07, 2.684257e-07, 2.684255e-07, 2.684262e-07, 
    2.68426e-07, 2.684261e-07, 2.684264e-07, 2.684256e-07, 2.68426e-07, 
    2.684253e-07, 2.684255e-07, 2.684249e-07, 2.684252e-07, 2.684246e-07, 
    2.684244e-07, 2.684241e-07, 2.684239e-07, 2.684262e-07, 2.684262e-07, 
    2.684261e-07, 2.684259e-07, 2.684257e-07, 2.684255e-07, 2.684255e-07, 
    2.684254e-07, 2.684253e-07, 2.684252e-07, 2.684254e-07, 2.684252e-07, 
    2.68426e-07, 2.684256e-07, 2.684263e-07, 2.684261e-07, 2.684259e-07, 
    2.68426e-07, 2.684257e-07, 2.684256e-07, 2.684253e-07, 2.684254e-07, 
    2.684244e-07, 2.684249e-07, 2.684236e-07, 2.68424e-07, 2.684263e-07, 
    2.684262e-07, 2.684258e-07, 2.68426e-07, 2.684255e-07, 2.684253e-07, 
    2.684252e-07, 2.684251e-07, 2.684251e-07, 2.68425e-07, 2.684251e-07, 
    2.68425e-07, 2.684255e-07, 2.684253e-07, 2.684259e-07, 2.684257e-07, 
    2.684258e-07, 2.684259e-07, 2.684256e-07, 2.684254e-07, 2.684254e-07, 
    2.684253e-07, 2.684251e-07, 2.684255e-07, 2.684244e-07, 2.684251e-07, 
    2.68426e-07, 2.684259e-07, 2.684258e-07, 2.684259e-07, 2.684254e-07, 
    2.684256e-07, 2.68425e-07, 2.684252e-07, 2.684249e-07, 2.684251e-07, 
    2.684251e-07, 2.684252e-07, 2.684253e-07, 2.684255e-07, 2.684257e-07, 
    2.684259e-07, 2.684259e-07, 2.684257e-07, 2.684254e-07, 2.684251e-07, 
    2.684252e-07, 2.684249e-07, 2.684255e-07, 2.684253e-07, 2.684254e-07, 
    2.684251e-07, 2.684257e-07, 2.684252e-07, 2.684258e-07, 2.684257e-07, 
    2.684256e-07, 2.684253e-07, 2.684252e-07, 2.684251e-07, 2.684252e-07, 
    2.684254e-07, 2.684254e-07, 2.684256e-07, 2.684256e-07, 2.684257e-07, 
    2.684258e-07, 2.684257e-07, 2.684256e-07, 2.684254e-07, 2.684251e-07, 
    2.684249e-07, 2.684248e-07, 2.684245e-07, 2.684248e-07, 2.684244e-07, 
    2.684247e-07, 2.684241e-07, 2.684252e-07, 2.684247e-07, 2.684255e-07, 
    2.684255e-07, 2.684253e-07, 2.684249e-07, 2.684251e-07, 2.684249e-07, 
    2.684254e-07, 2.684257e-07, 2.684258e-07, 2.684259e-07, 2.684257e-07, 
    2.684258e-07, 2.684256e-07, 2.684257e-07, 2.684254e-07, 2.684255e-07, 
    2.684251e-07, 2.684249e-07, 2.684244e-07, 2.684241e-07, 2.684238e-07, 
    2.684237e-07, 2.684236e-07, 2.684236e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  -3.431268e-26, -2.450906e-27, 8.82326e-26, 2.941087e-26, 5.146902e-26, 
    1.81367e-25, 1.200944e-25, 5.637083e-26, 7.107626e-26, 9.313441e-26, 
    1.225453e-26, -6.372354e-26, 1.593089e-25, -1.691125e-25, -1.740143e-25, 
    2.32836e-25, 2.352869e-25, 3.921449e-26, -1.02938e-25, 1.838179e-25, 
    -1.078398e-25, 2.132288e-25, 7.352717e-27, 1.176435e-25, -1.421525e-25, 
    2.450906e-27, -3.431268e-26, -1.02938e-25, 1.593089e-25, 3.921449e-26, 
    -4.901811e-27, -3.921449e-26, 7.352717e-27, -7.107626e-26, 6.372354e-26, 
    -1.56858e-25, 1.176435e-25, -1.372507e-25, 5.637083e-26, -1.02938e-25, 
    -2.132288e-25, -9.803622e-26, 4.65672e-26, -3.431268e-26, 8.82326e-26, 
    -1.102908e-25, -5.882173e-26, 1.789161e-25, -1.176435e-25, 1.81367e-25, 
    1.642107e-25, 2.401887e-25, 4.166539e-26, -1.715634e-26, 1.715634e-26, 
    2.034252e-25, 1.127417e-25, 1.225453e-25, -4.901811e-27, 2.573451e-25, 
    7.107626e-26, 1.54407e-25, -9.803622e-27, 2.034252e-25, -1.764652e-25, 
    -4.901811e-26, -1.421525e-25, -1.225453e-25, -1.838179e-25, 
    -3.063632e-25, 6.372354e-26, 5.637083e-26, -7.352717e-26, -2.32836e-25, 
    -1.225453e-25, 5.391992e-26, -1.323489e-25, -2.450906e-27, 1.666616e-25, 
    1.053889e-25, -1.372507e-25, -1.470543e-26, 8.333079e-26, -4.65672e-26, 
    2.450906e-25, -7.352717e-26, -1.470543e-26, -7.597807e-26, -8.333079e-26, 
    -1.666616e-25, 2.205815e-26, 1.176435e-25, 9.313441e-26, -2.32836e-25, 
    3.431268e-26, -1.053889e-25, 6.127264e-26, 1.715634e-26, 1.176435e-25, 
    -4.901811e-27, 4.901811e-26, -1.642107e-25, 2.205815e-26, -1.225453e-26, 
    1.225453e-25, 3.676358e-26, 8.82326e-26, 7.597807e-26, 8.578169e-26, 
    1.421525e-25, 1.495052e-25, -9.313441e-26, -4.901811e-27, -3.186177e-26, 
    1.249962e-25, 1.151926e-25, 7.352717e-26, -1.642107e-25, -2.695996e-26, 
    -3.676358e-26, -2.695996e-26, 5.391992e-26, -4.215557e-25, 1.200944e-25, 
    -3.235195e-25, -1.691125e-25, -1.740143e-25, -1.470543e-25, 8.82326e-26, 
    -7.842898e-26, -9.558531e-26, -1.715634e-26, 2.32836e-25, 7.352717e-27, 
    -2.450905e-26, 1.530638e-41, -5.882173e-26, 2.646978e-25, 2.892069e-25, 
    -1.078398e-25, -4.65672e-26, 8.087988e-26, -1.470543e-25, -2.401887e-25, 
    -1.495052e-25, -1.102908e-25, -1.176435e-25, -9.558531e-26, 8.578169e-26, 
    1.176435e-25, -8.087988e-26, -2.745014e-25, 0, -6.372354e-26, 
    2.32836e-25, 8.333079e-26, 1.887197e-25, 1.519561e-25, 2.622469e-25, 
    -1.519561e-25, 2.548942e-25, 2.058761e-25, 6.617445e-26, 1.715634e-25, 
    -1.421525e-25, 2.254833e-25, -2.450905e-26, 1.470543e-26, -1.519561e-25, 
    1.593089e-25, -1.225453e-26, -4.65672e-26, -1.642107e-25, -2.941087e-26, 
    -1.323489e-25, -7.842898e-26, 7.597807e-26, 7.597807e-26, 2.941087e-26, 
    5.146902e-26, -6.372354e-26, -4.41163e-26, -7.842898e-26, -9.803622e-27, 
    2.548942e-25, 1.838179e-25, -3.676358e-26, -3.186177e-26, -6.372354e-26, 
    2.401887e-25, 1.838179e-25, 6.127264e-26, -2.058761e-25, 1.666616e-25, 
    -6.372354e-26, 1.81367e-25, -1.323489e-25, -3.921449e-26, -1.274471e-25, 
    -2.156797e-25, 8.82326e-26, 7.842898e-26, -7.597807e-26, -1.151926e-25, 
    9.558531e-26, 7.352717e-27, -1.666616e-25, -7.352717e-26, -2.475414e-25, 
    1.225453e-26, -2.156797e-25, 3.921449e-26, -2.205815e-26, 8.333079e-26, 
    -6.127264e-26, -8.578169e-26, 1.519561e-25, 1.397016e-25, -1.176435e-25, 
    1.29898e-25, 9.068351e-26, 4.166539e-26, 2.695996e-26, 0, 4.901811e-27, 
    -2.941087e-26, -6.862535e-26, 1.960724e-25, 2.450905e-26, 1.960724e-26, 
    -2.646978e-25, -1.102908e-25, -1.372507e-25, -1.372507e-25, 
    -5.391992e-26, 6.372354e-26, -6.617445e-26, 1.274471e-25, -2.205815e-26, 
    1.764652e-25, -2.058761e-25, -6.372354e-26, 0, 7.842898e-26, 
    -3.039123e-25, -3.088141e-25, -2.205815e-26, -4.901811e-27, 1.789161e-25, 
    1.004871e-25, 2.32836e-25, 1.053889e-25, 2.205815e-26, 1.446034e-25, 
    -2.450906e-27, -7.842898e-26, 3.921449e-26, 8.82326e-26, 1.470543e-25, 
    -4.901811e-27, 1.81367e-25, -2.009742e-25, -9.558531e-26, 3.578322e-25, 
    1.02938e-25, 3.186177e-26, 2.254833e-25, -6.127264e-26, -3.480286e-25, 
    -7.352717e-27, -5.882173e-26, -6.862535e-26, 6.127264e-26, 1.053889e-25, 
    1.274471e-25, 1.715634e-26, 1.176435e-25, 1.29898e-25, 7.352717e-26, 
    1.54407e-25, -1.397016e-25, -9.803622e-26, -5.146902e-26, -4.166539e-26, 
    1.715634e-25, 4.901811e-26, -1.81367e-25, 1.960724e-26, 2.08327e-25, 
    -5.146902e-26, -1.446034e-25, -5.391992e-26, 8.82326e-26, 7.352717e-27, 
    2.401887e-25, 3.431268e-26, 1.789161e-25, -3.186177e-26, -6.372354e-26, 
    -7.352717e-27, -1.470543e-26, 2.034252e-25, 2.205815e-25, -3.676358e-26, 
    -9.803622e-26, -5.882173e-26, -1.985233e-25, 1.225453e-26, -7.352717e-27, 
    -8.578169e-26, -2.058761e-25, 1.29898e-25, 5.882173e-26, 1.470543e-26, 
    -1.54407e-25, 4.901811e-27, -6.862535e-26, -2.08327e-25, -1.421525e-25, 
    3.161668e-25, -1.715634e-25, -1.053889e-25, -1.495052e-25, -7.107626e-26, 
    2.941087e-26, -2.499924e-25, -7.107626e-26, 3.284213e-25, 2.377378e-25, 
    -1.078398e-25, 1.530638e-41, -3.186177e-26, -1.078398e-25, 6.127264e-26, 
    -1.715634e-26, 8.087988e-26, -1.225453e-25, 6.372354e-26,
  2.676255e-32, 2.676252e-32, 2.676253e-32, 2.676251e-32, 2.676252e-32, 
    2.67625e-32, 2.676254e-32, 2.676252e-32, 2.676254e-32, 2.676255e-32, 
    2.676246e-32, 2.676251e-32, 2.676242e-32, 2.676244e-32, 2.676238e-32, 
    2.676242e-32, 2.676237e-32, 2.676238e-32, 2.676235e-32, 2.676236e-32, 
    2.676232e-32, 2.676234e-32, 2.67623e-32, 2.676232e-32, 2.676232e-32, 
    2.676234e-32, 2.67625e-32, 2.676247e-32, 2.67625e-32, 2.676249e-32, 
    2.676249e-32, 2.676252e-32, 2.676253e-32, 2.676255e-32, 2.676255e-32, 
    2.676253e-32, 2.676249e-32, 2.676251e-32, 2.676247e-32, 2.676247e-32, 
    2.676244e-32, 2.676245e-32, 2.676239e-32, 2.676241e-32, 2.676236e-32, 
    2.676237e-32, 2.676236e-32, 2.676236e-32, 2.676236e-32, 2.676238e-32, 
    2.676237e-32, 2.676239e-32, 2.676245e-32, 2.676243e-32, 2.676249e-32, 
    2.676252e-32, 2.676254e-32, 2.676256e-32, 2.676256e-32, 2.676255e-32, 
    2.676253e-32, 2.676251e-32, 2.676249e-32, 2.676248e-32, 2.676247e-32, 
    2.676244e-32, 2.676242e-32, 2.676239e-32, 2.676239e-32, 2.676238e-32, 
    2.676237e-32, 2.676235e-32, 2.676236e-32, 2.676235e-32, 2.676238e-32, 
    2.676236e-32, 2.67624e-32, 2.676239e-32, 2.676247e-32, 2.67625e-32, 
    2.676252e-32, 2.676253e-32, 2.676256e-32, 2.676254e-32, 2.676254e-32, 
    2.676252e-32, 2.676251e-32, 2.676252e-32, 2.676248e-32, 2.67625e-32, 
    2.676242e-32, 2.676246e-32, 2.676237e-32, 2.676239e-32, 2.676237e-32, 
    2.676238e-32, 2.676236e-32, 2.676238e-32, 2.676234e-32, 2.676234e-32, 
    2.676234e-32, 2.676232e-32, 2.676238e-32, 2.676236e-32, 2.676252e-32, 
    2.676252e-32, 2.676252e-32, 2.676253e-32, 2.676254e-32, 2.676255e-32, 
    2.676254e-32, 2.676253e-32, 2.676251e-32, 2.67625e-32, 2.676249e-32, 
    2.676247e-32, 2.676245e-32, 2.676242e-32, 2.676239e-32, 2.676237e-32, 
    2.676239e-32, 2.676238e-32, 2.676239e-32, 2.676239e-32, 2.676234e-32, 
    2.676237e-32, 2.676233e-32, 2.676233e-32, 2.676235e-32, 2.676233e-32, 
    2.676252e-32, 2.676252e-32, 2.676254e-32, 2.676253e-32, 2.676255e-32, 
    2.676254e-32, 2.676253e-32, 2.67625e-32, 2.676249e-32, 2.676248e-32, 
    2.676247e-32, 2.676245e-32, 2.676242e-32, 2.676239e-32, 2.676237e-32, 
    2.676237e-32, 2.676237e-32, 2.676237e-32, 2.676238e-32, 2.676237e-32, 
    2.676236e-32, 2.676237e-32, 2.676233e-32, 2.676234e-32, 2.676233e-32, 
    2.676234e-32, 2.676252e-32, 2.676251e-32, 2.676252e-32, 2.676251e-32, 
    2.676252e-32, 2.676249e-32, 2.676248e-32, 2.676244e-32, 2.676245e-32, 
    2.676242e-32, 2.676245e-32, 2.676244e-32, 2.676242e-32, 2.676245e-32, 
    2.67624e-32, 2.676243e-32, 2.676237e-32, 2.67624e-32, 2.676237e-32, 
    2.676237e-32, 2.676236e-32, 2.676235e-32, 2.676234e-32, 2.676232e-32, 
    2.676232e-32, 2.67623e-32, 2.67625e-32, 2.676249e-32, 2.676249e-32, 
    2.676247e-32, 2.676247e-32, 2.676244e-32, 2.676242e-32, 2.676243e-32, 
    2.67624e-32, 2.67624e-32, 2.676243e-32, 2.676241e-32, 2.676248e-32, 
    2.676247e-32, 2.676247e-32, 2.67625e-32, 2.676242e-32, 2.676246e-32, 
    2.676239e-32, 2.676241e-32, 2.676235e-32, 2.676238e-32, 2.676232e-32, 
    2.67623e-32, 2.676227e-32, 2.676224e-32, 2.676248e-32, 2.676249e-32, 
    2.676247e-32, 2.676245e-32, 2.676244e-32, 2.676241e-32, 2.676241e-32, 
    2.67624e-32, 2.676239e-32, 2.676238e-32, 2.67624e-32, 2.676238e-32, 
    2.676247e-32, 2.676242e-32, 2.676249e-32, 2.676247e-32, 2.676245e-32, 
    2.676246e-32, 2.676243e-32, 2.676242e-32, 2.676239e-32, 2.67624e-32, 
    2.67623e-32, 2.676235e-32, 2.676222e-32, 2.676226e-32, 2.676249e-32, 
    2.676248e-32, 2.676244e-32, 2.676246e-32, 2.676241e-32, 2.676239e-32, 
    2.676239e-32, 2.676237e-32, 2.676237e-32, 2.676236e-32, 2.676238e-32, 
    2.676236e-32, 2.676241e-32, 2.676239e-32, 2.676245e-32, 2.676243e-32, 
    2.676244e-32, 2.676244e-32, 2.676242e-32, 2.67624e-32, 2.67624e-32, 
    2.676239e-32, 2.676237e-32, 2.676241e-32, 2.67623e-32, 2.676237e-32, 
    2.676247e-32, 2.676245e-32, 2.676244e-32, 2.676245e-32, 2.67624e-32, 
    2.676242e-32, 2.676236e-32, 2.676238e-32, 2.676235e-32, 2.676237e-32, 
    2.676237e-32, 2.676238e-32, 2.676239e-32, 2.676242e-32, 2.676244e-32, 
    2.676245e-32, 2.676245e-32, 2.676243e-32, 2.67624e-32, 2.676237e-32, 
    2.676238e-32, 2.676236e-32, 2.676241e-32, 2.676239e-32, 2.67624e-32, 
    2.676237e-32, 2.676243e-32, 2.676238e-32, 2.676244e-32, 2.676243e-32, 
    2.676242e-32, 2.676239e-32, 2.676238e-32, 2.676237e-32, 2.676238e-32, 
    2.67624e-32, 2.67624e-32, 2.676242e-32, 2.676242e-32, 2.676243e-32, 
    2.676244e-32, 2.676244e-32, 2.676242e-32, 2.67624e-32, 2.676237e-32, 
    2.676235e-32, 2.676234e-32, 2.676231e-32, 2.676234e-32, 2.67623e-32, 
    2.676233e-32, 2.676227e-32, 2.676238e-32, 2.676233e-32, 2.676242e-32, 
    2.676241e-32, 2.676239e-32, 2.676235e-32, 2.676237e-32, 2.676235e-32, 
    2.67624e-32, 2.676243e-32, 2.676244e-32, 2.676245e-32, 2.676244e-32, 
    2.676244e-32, 2.676242e-32, 2.676243e-32, 2.67624e-32, 2.676242e-32, 
    2.676237e-32, 2.676235e-32, 2.67623e-32, 2.676227e-32, 2.676224e-32, 
    2.676223e-32, 2.676222e-32, 2.676222e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.325088e-15, 3.334083e-15, 3.332336e-15, 3.339583e-15, 3.335565e-15, 
    3.340309e-15, 3.326914e-15, 3.334439e-15, 3.329637e-15, 3.3259e-15, 
    3.353627e-15, 3.339907e-15, 3.367866e-15, 3.359131e-15, 3.381058e-15, 
    3.366506e-15, 3.38399e-15, 3.380641e-15, 3.390721e-15, 3.387835e-15, 
    3.400707e-15, 3.392053e-15, 3.407376e-15, 3.398643e-15, 3.400009e-15, 
    3.391767e-15, 3.342672e-15, 3.351919e-15, 3.342124e-15, 3.343443e-15, 
    3.342852e-15, 3.335647e-15, 3.332012e-15, 3.324403e-15, 3.325785e-15, 
    3.331375e-15, 3.344036e-15, 3.339742e-15, 3.350565e-15, 3.350321e-15, 
    3.362353e-15, 3.35693e-15, 3.377127e-15, 3.371393e-15, 3.387955e-15, 
    3.383793e-15, 3.38776e-15, 3.386557e-15, 3.387775e-15, 3.38167e-15, 
    3.384286e-15, 3.378912e-15, 3.357945e-15, 3.364112e-15, 3.345705e-15, 
    3.334612e-15, 3.327244e-15, 3.322009e-15, 3.322749e-15, 3.324159e-15, 
    3.331407e-15, 3.338218e-15, 3.343404e-15, 3.346871e-15, 3.350286e-15, 
    3.360607e-15, 3.36607e-15, 3.378285e-15, 3.376084e-15, 3.379814e-15, 
    3.383379e-15, 3.389357e-15, 3.388374e-15, 3.391006e-15, 3.379717e-15, 
    3.387221e-15, 3.37483e-15, 3.378221e-15, 3.351205e-15, 3.340901e-15, 
    3.33651e-15, 3.332671e-15, 3.323318e-15, 3.329778e-15, 3.327232e-15, 
    3.33329e-15, 3.337136e-15, 3.335234e-15, 3.346966e-15, 3.342407e-15, 
    3.366394e-15, 3.356071e-15, 3.382963e-15, 3.376536e-15, 3.384503e-15, 
    3.380439e-15, 3.3874e-15, 3.381136e-15, 3.391986e-15, 3.394345e-15, 
    3.392733e-15, 3.398928e-15, 3.380788e-15, 3.387759e-15, 3.33518e-15, 
    3.33549e-15, 3.336936e-15, 3.33058e-15, 3.330191e-15, 3.324364e-15, 
    3.32955e-15, 3.331756e-15, 3.337359e-15, 3.34067e-15, 3.343816e-15, 
    3.35073e-15, 3.358443e-15, 3.369219e-15, 3.376953e-15, 3.382133e-15, 
    3.378958e-15, 3.381761e-15, 3.378627e-15, 3.377158e-15, 3.393461e-15, 
    3.38431e-15, 3.398037e-15, 3.397279e-15, 3.391068e-15, 3.397364e-15, 
    3.335708e-15, 3.333923e-15, 3.327721e-15, 3.332575e-15, 3.32373e-15, 
    3.328681e-15, 3.331526e-15, 3.3425e-15, 3.344911e-15, 3.347144e-15, 
    3.351553e-15, 3.357208e-15, 3.367117e-15, 3.37573e-15, 3.383587e-15, 
    3.383011e-15, 3.383214e-15, 3.384967e-15, 3.380623e-15, 3.38568e-15, 
    3.386528e-15, 3.38431e-15, 3.397177e-15, 3.393503e-15, 3.397263e-15, 
    3.394871e-15, 3.334504e-15, 3.337507e-15, 3.335884e-15, 3.338935e-15, 
    3.336785e-15, 3.346339e-15, 3.349201e-15, 3.362583e-15, 3.357096e-15, 
    3.365829e-15, 3.357984e-15, 3.359374e-15, 3.36611e-15, 3.358409e-15, 
    3.375254e-15, 3.363834e-15, 3.385035e-15, 3.373641e-15, 3.385748e-15, 
    3.383553e-15, 3.387189e-15, 3.390442e-15, 3.394536e-15, 3.40208e-15, 
    3.400334e-15, 3.406641e-15, 3.341983e-15, 3.345874e-15, 3.345533e-15, 
    3.349605e-15, 3.352614e-15, 3.359135e-15, 3.36958e-15, 3.365655e-15, 
    3.372862e-15, 3.374308e-15, 3.363358e-15, 3.370081e-15, 3.348479e-15, 
    3.351971e-15, 3.349893e-15, 3.342289e-15, 3.366557e-15, 3.354111e-15, 
    3.377081e-15, 3.370349e-15, 3.389978e-15, 3.380221e-15, 3.399373e-15, 
    3.40754e-15, 3.415228e-15, 3.424192e-15, 3.347999e-15, 3.345356e-15, 
    3.350089e-15, 3.356631e-15, 3.3627e-15, 3.37076e-15, 3.371585e-15, 
    3.373093e-15, 3.377001e-15, 3.380284e-15, 3.373568e-15, 3.381108e-15, 
    3.352777e-15, 3.367637e-15, 3.344355e-15, 3.35137e-15, 3.356246e-15, 
    3.354109e-15, 3.365206e-15, 3.367819e-15, 3.378426e-15, 3.372946e-15, 
    3.405524e-15, 3.391127e-15, 3.431016e-15, 3.419889e-15, 3.344432e-15, 
    3.347991e-15, 3.360362e-15, 3.354479e-15, 3.371298e-15, 3.375433e-15, 
    3.378793e-15, 3.383084e-15, 3.383549e-15, 3.38609e-15, 3.381925e-15, 
    3.385926e-15, 3.370777e-15, 3.377551e-15, 3.358951e-15, 3.363481e-15, 
    3.361398e-15, 3.359111e-15, 3.366167e-15, 3.373674e-15, 3.373837e-15, 
    3.376242e-15, 3.383011e-15, 3.371367e-15, 3.407375e-15, 3.385152e-15, 
    3.351869e-15, 3.358713e-15, 3.359694e-15, 3.357043e-15, 3.375018e-15, 
    3.368509e-15, 3.386029e-15, 3.381298e-15, 3.389048e-15, 3.385198e-15, 
    3.384631e-15, 3.379683e-15, 3.3766e-15, 3.368807e-15, 3.362462e-15, 
    3.357428e-15, 3.358599e-15, 3.364128e-15, 3.374133e-15, 3.38359e-15, 
    3.381519e-15, 3.388459e-15, 3.37008e-15, 3.377791e-15, 3.37481e-15, 
    3.382579e-15, 3.36555e-15, 3.380045e-15, 3.361839e-15, 3.363438e-15, 
    3.36838e-15, 3.378311e-15, 3.380511e-15, 3.382854e-15, 3.381409e-15, 
    3.374388e-15, 3.373238e-15, 3.368261e-15, 3.366885e-15, 3.36309e-15, 
    3.359946e-15, 3.362818e-15, 3.365832e-15, 3.374392e-15, 3.382096e-15, 
    3.390488e-15, 3.392542e-15, 3.402326e-15, 3.394358e-15, 3.407498e-15, 
    3.396322e-15, 3.41566e-15, 3.380889e-15, 3.395999e-15, 3.368606e-15, 
    3.371562e-15, 3.376904e-15, 3.389147e-15, 3.382543e-15, 3.390268e-15, 
    3.373193e-15, 3.364317e-15, 3.362022e-15, 3.357733e-15, 3.36212e-15, 
    3.361764e-15, 3.365959e-15, 3.364611e-15, 3.374676e-15, 3.369271e-15, 
    3.384616e-15, 3.390207e-15, 3.405979e-15, 3.415629e-15, 3.425445e-15, 
    3.429772e-15, 3.431089e-15, 3.431639e-15 ;

 LITR2N_vr =
  1.532745e-05, 1.532744e-05, 1.532744e-05, 1.532743e-05, 1.532743e-05, 
    1.532742e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 1.532745e-05, 
    1.53274e-05, 1.532743e-05, 1.532738e-05, 1.532739e-05, 1.532735e-05, 
    1.532738e-05, 1.532735e-05, 1.532736e-05, 1.532734e-05, 1.532734e-05, 
    1.532732e-05, 1.532734e-05, 1.532731e-05, 1.532732e-05, 1.532732e-05, 
    1.532734e-05, 1.532742e-05, 1.53274e-05, 1.532742e-05, 1.532742e-05, 
    1.532742e-05, 1.532743e-05, 1.532744e-05, 1.532745e-05, 1.532745e-05, 
    1.532744e-05, 1.532742e-05, 1.532743e-05, 1.532741e-05, 1.532741e-05, 
    1.532739e-05, 1.53274e-05, 1.532736e-05, 1.532737e-05, 1.532734e-05, 
    1.532735e-05, 1.532734e-05, 1.532734e-05, 1.532734e-05, 1.532735e-05, 
    1.532735e-05, 1.532736e-05, 1.532739e-05, 1.532738e-05, 1.532742e-05, 
    1.532744e-05, 1.532745e-05, 1.532746e-05, 1.532746e-05, 1.532745e-05, 
    1.532744e-05, 1.532743e-05, 1.532742e-05, 1.532741e-05, 1.532741e-05, 
    1.532739e-05, 1.532738e-05, 1.532736e-05, 1.532736e-05, 1.532736e-05, 
    1.532735e-05, 1.532734e-05, 1.532734e-05, 1.532734e-05, 1.532736e-05, 
    1.532734e-05, 1.532736e-05, 1.532736e-05, 1.532741e-05, 1.532742e-05, 
    1.532743e-05, 1.532744e-05, 1.532746e-05, 1.532744e-05, 1.532745e-05, 
    1.532744e-05, 1.532743e-05, 1.532743e-05, 1.532741e-05, 1.532742e-05, 
    1.532738e-05, 1.53274e-05, 1.532735e-05, 1.532736e-05, 1.532735e-05, 
    1.532736e-05, 1.532734e-05, 1.532735e-05, 1.532734e-05, 1.532733e-05, 
    1.532733e-05, 1.532732e-05, 1.532736e-05, 1.532734e-05, 1.532743e-05, 
    1.532743e-05, 1.532743e-05, 1.532744e-05, 1.532744e-05, 1.532745e-05, 
    1.532744e-05, 1.532744e-05, 1.532743e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.532739e-05, 1.532738e-05, 1.532736e-05, 1.532735e-05, 
    1.532736e-05, 1.532735e-05, 1.532736e-05, 1.532736e-05, 1.532733e-05, 
    1.532735e-05, 1.532732e-05, 1.532733e-05, 1.532734e-05, 1.532733e-05, 
    1.532743e-05, 1.532744e-05, 1.532745e-05, 1.532744e-05, 1.532745e-05, 
    1.532745e-05, 1.532744e-05, 1.532742e-05, 1.532742e-05, 1.532741e-05, 
    1.532741e-05, 1.53274e-05, 1.532738e-05, 1.532736e-05, 1.532735e-05, 
    1.532735e-05, 1.532735e-05, 1.532735e-05, 1.532736e-05, 1.532735e-05, 
    1.532734e-05, 1.532735e-05, 1.532733e-05, 1.532733e-05, 1.532733e-05, 
    1.532733e-05, 1.532744e-05, 1.532743e-05, 1.532743e-05, 1.532743e-05, 
    1.532743e-05, 1.532742e-05, 1.532741e-05, 1.532739e-05, 1.53274e-05, 
    1.532738e-05, 1.532739e-05, 1.532739e-05, 1.532738e-05, 1.532739e-05, 
    1.532736e-05, 1.532738e-05, 1.532735e-05, 1.532737e-05, 1.532735e-05, 
    1.532735e-05, 1.532734e-05, 1.532734e-05, 1.532733e-05, 1.532732e-05, 
    1.532732e-05, 1.532731e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.53274e-05, 1.532739e-05, 1.532737e-05, 1.532738e-05, 
    1.532737e-05, 1.532737e-05, 1.532738e-05, 1.532737e-05, 1.532741e-05, 
    1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532738e-05, 1.53274e-05, 
    1.532736e-05, 1.532737e-05, 1.532734e-05, 1.532736e-05, 1.532732e-05, 
    1.532731e-05, 1.532729e-05, 1.532728e-05, 1.532741e-05, 1.532742e-05, 
    1.532741e-05, 1.53274e-05, 1.532739e-05, 1.532737e-05, 1.532737e-05, 
    1.532737e-05, 1.532736e-05, 1.532736e-05, 1.532737e-05, 1.532735e-05, 
    1.53274e-05, 1.532738e-05, 1.532742e-05, 1.532741e-05, 1.53274e-05, 
    1.53274e-05, 1.532738e-05, 1.532738e-05, 1.532736e-05, 1.532737e-05, 
    1.532731e-05, 1.532734e-05, 1.532727e-05, 1.532729e-05, 1.532742e-05, 
    1.532741e-05, 1.532739e-05, 1.53274e-05, 1.532737e-05, 1.532736e-05, 
    1.532736e-05, 1.532735e-05, 1.532735e-05, 1.532734e-05, 1.532735e-05, 
    1.532735e-05, 1.532737e-05, 1.532736e-05, 1.532739e-05, 1.532738e-05, 
    1.532739e-05, 1.532739e-05, 1.532738e-05, 1.532737e-05, 1.532737e-05, 
    1.532736e-05, 1.532735e-05, 1.532737e-05, 1.532731e-05, 1.532735e-05, 
    1.53274e-05, 1.532739e-05, 1.532739e-05, 1.53274e-05, 1.532736e-05, 
    1.532738e-05, 1.532735e-05, 1.532735e-05, 1.532734e-05, 1.532735e-05, 
    1.532735e-05, 1.532736e-05, 1.532736e-05, 1.532738e-05, 1.532739e-05, 
    1.53274e-05, 1.532739e-05, 1.532738e-05, 1.532737e-05, 1.532735e-05, 
    1.532735e-05, 1.532734e-05, 1.532737e-05, 1.532736e-05, 1.532736e-05, 
    1.532735e-05, 1.532738e-05, 1.532736e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532736e-05, 1.532736e-05, 1.532735e-05, 1.532735e-05, 
    1.532737e-05, 1.532737e-05, 1.532738e-05, 1.532738e-05, 1.532739e-05, 
    1.532739e-05, 1.532739e-05, 1.532738e-05, 1.532737e-05, 1.532735e-05, 
    1.532734e-05, 1.532733e-05, 1.532732e-05, 1.532733e-05, 1.532731e-05, 
    1.532733e-05, 1.532729e-05, 1.532735e-05, 1.532733e-05, 1.532738e-05, 
    1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532735e-05, 1.532734e-05, 
    1.532737e-05, 1.532738e-05, 1.532739e-05, 1.53274e-05, 1.532739e-05, 
    1.532739e-05, 1.532738e-05, 1.532738e-05, 1.532736e-05, 1.532738e-05, 
    1.532735e-05, 1.532734e-05, 1.532731e-05, 1.532729e-05, 1.532728e-05, 
    1.532727e-05, 1.532727e-05, 1.532727e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.201324e-13, 1.204574e-13, 1.203942e-13, 1.206561e-13, 1.205109e-13, 
    1.206823e-13, 1.201984e-13, 1.204702e-13, 1.202967e-13, 1.201617e-13, 
    1.211635e-13, 1.206678e-13, 1.216779e-13, 1.213624e-13, 1.221545e-13, 
    1.216288e-13, 1.222605e-13, 1.221395e-13, 1.225037e-13, 1.223994e-13, 
    1.228644e-13, 1.225518e-13, 1.231054e-13, 1.227899e-13, 1.228392e-13, 
    1.225414e-13, 1.207677e-13, 1.211018e-13, 1.207479e-13, 1.207955e-13, 
    1.207742e-13, 1.205139e-13, 1.203825e-13, 1.201076e-13, 1.201576e-13, 
    1.203595e-13, 1.20817e-13, 1.206618e-13, 1.210529e-13, 1.21044e-13, 
    1.214787e-13, 1.212828e-13, 1.220125e-13, 1.218053e-13, 1.224037e-13, 
    1.222533e-13, 1.223967e-13, 1.223532e-13, 1.223972e-13, 1.221766e-13, 
    1.222712e-13, 1.22077e-13, 1.213195e-13, 1.215423e-13, 1.208773e-13, 
    1.204765e-13, 1.202103e-13, 1.200211e-13, 1.200479e-13, 1.200988e-13, 
    1.203607e-13, 1.206068e-13, 1.207941e-13, 1.209194e-13, 1.210428e-13, 
    1.214157e-13, 1.21613e-13, 1.220544e-13, 1.219748e-13, 1.221096e-13, 
    1.222384e-13, 1.224544e-13, 1.224188e-13, 1.225139e-13, 1.221061e-13, 
    1.223772e-13, 1.219295e-13, 1.22052e-13, 1.21076e-13, 1.207037e-13, 
    1.205451e-13, 1.204064e-13, 1.200684e-13, 1.203018e-13, 1.202098e-13, 
    1.204287e-13, 1.205677e-13, 1.20499e-13, 1.209228e-13, 1.207581e-13, 
    1.216247e-13, 1.212518e-13, 1.222234e-13, 1.219912e-13, 1.22279e-13, 
    1.221322e-13, 1.223837e-13, 1.221574e-13, 1.225494e-13, 1.226346e-13, 
    1.225763e-13, 1.228002e-13, 1.221448e-13, 1.223966e-13, 1.20497e-13, 
    1.205082e-13, 1.205604e-13, 1.203308e-13, 1.203168e-13, 1.201062e-13, 
    1.202936e-13, 1.203733e-13, 1.205757e-13, 1.206953e-13, 1.20809e-13, 
    1.210588e-13, 1.213375e-13, 1.217268e-13, 1.220062e-13, 1.221934e-13, 
    1.220787e-13, 1.221799e-13, 1.220667e-13, 1.220136e-13, 1.226026e-13, 
    1.22272e-13, 1.22768e-13, 1.227406e-13, 1.225162e-13, 1.227437e-13, 
    1.205161e-13, 1.204516e-13, 1.202275e-13, 1.204029e-13, 1.200833e-13, 
    1.202622e-13, 1.20365e-13, 1.207615e-13, 1.208486e-13, 1.209292e-13, 
    1.210886e-13, 1.212928e-13, 1.216509e-13, 1.219621e-13, 1.222459e-13, 
    1.222251e-13, 1.222324e-13, 1.222958e-13, 1.221388e-13, 1.223215e-13, 
    1.223521e-13, 1.22272e-13, 1.227369e-13, 1.226042e-13, 1.2274e-13, 
    1.226536e-13, 1.204726e-13, 1.205811e-13, 1.205224e-13, 1.206327e-13, 
    1.20555e-13, 1.209002e-13, 1.210036e-13, 1.21487e-13, 1.212888e-13, 
    1.216043e-13, 1.213209e-13, 1.213711e-13, 1.216145e-13, 1.213362e-13, 
    1.219448e-13, 1.215322e-13, 1.222982e-13, 1.218866e-13, 1.22324e-13, 
    1.222447e-13, 1.22376e-13, 1.224936e-13, 1.226415e-13, 1.22914e-13, 
    1.22851e-13, 1.230788e-13, 1.207428e-13, 1.208834e-13, 1.208711e-13, 
    1.210182e-13, 1.211269e-13, 1.213625e-13, 1.217399e-13, 1.21598e-13, 
    1.218584e-13, 1.219107e-13, 1.215151e-13, 1.21758e-13, 1.209775e-13, 
    1.211036e-13, 1.210286e-13, 1.207539e-13, 1.216306e-13, 1.21181e-13, 
    1.220108e-13, 1.217677e-13, 1.224768e-13, 1.221243e-13, 1.228162e-13, 
    1.231113e-13, 1.233891e-13, 1.237129e-13, 1.209601e-13, 1.208646e-13, 
    1.210357e-13, 1.21272e-13, 1.214913e-13, 1.217825e-13, 1.218123e-13, 
    1.218668e-13, 1.22008e-13, 1.221266e-13, 1.218839e-13, 1.221563e-13, 
    1.211328e-13, 1.216697e-13, 1.208285e-13, 1.210819e-13, 1.212581e-13, 
    1.211809e-13, 1.215818e-13, 1.216762e-13, 1.220595e-13, 1.218615e-13, 
    1.230385e-13, 1.225183e-13, 1.239595e-13, 1.235575e-13, 1.208313e-13, 
    1.209598e-13, 1.214068e-13, 1.211942e-13, 1.218019e-13, 1.219513e-13, 
    1.220727e-13, 1.222277e-13, 1.222445e-13, 1.223363e-13, 1.221859e-13, 
    1.223304e-13, 1.217831e-13, 1.220278e-13, 1.213558e-13, 1.215195e-13, 
    1.214443e-13, 1.213616e-13, 1.216165e-13, 1.218878e-13, 1.218937e-13, 
    1.219805e-13, 1.222251e-13, 1.218044e-13, 1.231053e-13, 1.223025e-13, 
    1.211e-13, 1.213472e-13, 1.213827e-13, 1.212869e-13, 1.219363e-13, 
    1.217012e-13, 1.223341e-13, 1.221632e-13, 1.224432e-13, 1.223041e-13, 
    1.222836e-13, 1.221049e-13, 1.219935e-13, 1.217119e-13, 1.214827e-13, 
    1.213008e-13, 1.213431e-13, 1.215429e-13, 1.219044e-13, 1.22246e-13, 
    1.221712e-13, 1.224219e-13, 1.217579e-13, 1.220365e-13, 1.219288e-13, 
    1.222095e-13, 1.215942e-13, 1.221179e-13, 1.214602e-13, 1.215179e-13, 
    1.216965e-13, 1.220553e-13, 1.221348e-13, 1.222194e-13, 1.221672e-13, 
    1.219135e-13, 1.21872e-13, 1.216922e-13, 1.216425e-13, 1.215054e-13, 
    1.213918e-13, 1.214955e-13, 1.216045e-13, 1.219137e-13, 1.221921e-13, 
    1.224952e-13, 1.225694e-13, 1.229229e-13, 1.226351e-13, 1.231098e-13, 
    1.22706e-13, 1.234047e-13, 1.221484e-13, 1.226943e-13, 1.217046e-13, 
    1.218115e-13, 1.220044e-13, 1.224468e-13, 1.222082e-13, 1.224873e-13, 
    1.218704e-13, 1.215497e-13, 1.214668e-13, 1.213118e-13, 1.214703e-13, 
    1.214575e-13, 1.21609e-13, 1.215603e-13, 1.21924e-13, 1.217287e-13, 
    1.222831e-13, 1.224851e-13, 1.230549e-13, 1.234036e-13, 1.237582e-13, 
    1.239145e-13, 1.239621e-13, 1.23982e-13 ;

 LITR3C =
  9.698016e-06, 9.698006e-06, 9.698007e-06, 9.697999e-06, 9.698004e-06, 
    9.697998e-06, 9.698013e-06, 9.698005e-06, 9.69801e-06, 9.698015e-06, 
    9.697984e-06, 9.697999e-06, 9.697968e-06, 9.697977e-06, 9.697954e-06, 
    9.697969e-06, 9.69795e-06, 9.697954e-06, 9.697943e-06, 9.697946e-06, 
    9.697932e-06, 9.697941e-06, 9.697925e-06, 9.697934e-06, 9.697933e-06, 
    9.697942e-06, 9.697996e-06, 9.697986e-06, 9.697997e-06, 9.697995e-06, 
    9.697996e-06, 9.698004e-06, 9.698007e-06, 9.698016e-06, 9.698015e-06, 
    9.698008e-06, 9.697995e-06, 9.697999e-06, 9.697987e-06, 9.697987e-06, 
    9.697974e-06, 9.69798e-06, 9.697957e-06, 9.697964e-06, 9.697946e-06, 
    9.69795e-06, 9.697946e-06, 9.697947e-06, 9.697946e-06, 9.697953e-06, 
    9.69795e-06, 9.697956e-06, 9.697979e-06, 9.697972e-06, 9.697993e-06, 
    9.698005e-06, 9.698013e-06, 9.698018e-06, 9.698017e-06, 9.698017e-06, 
    9.698008e-06, 9.698001e-06, 9.697995e-06, 9.697991e-06, 9.697987e-06, 
    9.697976e-06, 9.69797e-06, 9.697957e-06, 9.697959e-06, 9.697955e-06, 
    9.697951e-06, 9.697945e-06, 9.697946e-06, 9.697943e-06, 9.697955e-06, 
    9.697947e-06, 9.69796e-06, 9.697957e-06, 9.697987e-06, 9.697997e-06, 
    9.698003e-06, 9.698007e-06, 9.698017e-06, 9.69801e-06, 9.698013e-06, 
    9.698007e-06, 9.698002e-06, 9.698004e-06, 9.697991e-06, 9.697997e-06, 
    9.697969e-06, 9.697981e-06, 9.697951e-06, 9.697958e-06, 9.697949e-06, 
    9.697954e-06, 9.697947e-06, 9.697954e-06, 9.697941e-06, 9.697938e-06, 
    9.69794e-06, 9.697934e-06, 9.697954e-06, 9.697946e-06, 9.698004e-06, 
    9.698004e-06, 9.698002e-06, 9.698009e-06, 9.698009e-06, 9.698016e-06, 
    9.69801e-06, 9.698007e-06, 9.698002e-06, 9.697998e-06, 9.697995e-06, 
    9.697987e-06, 9.697978e-06, 9.697967e-06, 9.697958e-06, 9.697952e-06, 
    9.697956e-06, 9.697953e-06, 9.697957e-06, 9.697957e-06, 9.69794e-06, 
    9.69795e-06, 9.697935e-06, 9.697936e-06, 9.697942e-06, 9.697936e-06, 
    9.698004e-06, 9.698006e-06, 9.698012e-06, 9.698007e-06, 9.698017e-06, 
    9.698011e-06, 9.698008e-06, 9.697996e-06, 9.697993e-06, 9.697991e-06, 
    9.697986e-06, 9.69798e-06, 9.697969e-06, 9.697959e-06, 9.697951e-06, 
    9.697951e-06, 9.697951e-06, 9.697949e-06, 9.697954e-06, 9.697948e-06, 
    9.697947e-06, 9.69795e-06, 9.697936e-06, 9.697939e-06, 9.697936e-06, 
    9.697938e-06, 9.698005e-06, 9.698001e-06, 9.698003e-06, 9.698e-06, 
    9.698002e-06, 9.697992e-06, 9.697988e-06, 9.697974e-06, 9.69798e-06, 
    9.69797e-06, 9.697979e-06, 9.697977e-06, 9.69797e-06, 9.697978e-06, 
    9.69796e-06, 9.697973e-06, 9.697949e-06, 9.697962e-06, 9.697948e-06, 
    9.697951e-06, 9.697947e-06, 9.697943e-06, 9.697938e-06, 9.69793e-06, 
    9.697932e-06, 9.697926e-06, 9.697997e-06, 9.697992e-06, 9.697993e-06, 
    9.697988e-06, 9.697985e-06, 9.697977e-06, 9.697967e-06, 9.69797e-06, 
    9.697963e-06, 9.697961e-06, 9.697973e-06, 9.697966e-06, 9.697989e-06, 
    9.697986e-06, 9.697987e-06, 9.697997e-06, 9.697969e-06, 9.697983e-06, 
    9.697957e-06, 9.697966e-06, 9.697944e-06, 9.697955e-06, 9.697933e-06, 
    9.697924e-06, 9.697916e-06, 9.697906e-06, 9.69799e-06, 9.697993e-06, 
    9.697987e-06, 9.69798e-06, 9.697974e-06, 9.697965e-06, 9.697964e-06, 
    9.697962e-06, 9.697958e-06, 9.697955e-06, 9.697962e-06, 9.697954e-06, 
    9.697985e-06, 9.697968e-06, 9.697994e-06, 9.697987e-06, 9.697981e-06, 
    9.697983e-06, 9.697971e-06, 9.697968e-06, 9.697957e-06, 9.697962e-06, 
    9.697927e-06, 9.697942e-06, 9.697898e-06, 9.69791e-06, 9.697994e-06, 
    9.69799e-06, 9.697977e-06, 9.697983e-06, 9.697964e-06, 9.697959e-06, 
    9.697956e-06, 9.697951e-06, 9.697951e-06, 9.697947e-06, 9.697953e-06, 
    9.697948e-06, 9.697965e-06, 9.697957e-06, 9.697977e-06, 9.697973e-06, 
    9.697975e-06, 9.697977e-06, 9.69797e-06, 9.697962e-06, 9.697961e-06, 
    9.697958e-06, 9.697951e-06, 9.697964e-06, 9.697925e-06, 9.697949e-06, 
    9.697986e-06, 9.697978e-06, 9.697977e-06, 9.69798e-06, 9.69796e-06, 
    9.697967e-06, 9.697948e-06, 9.697953e-06, 9.697945e-06, 9.697949e-06, 
    9.697949e-06, 9.697955e-06, 9.697958e-06, 9.697967e-06, 9.697974e-06, 
    9.697979e-06, 9.697978e-06, 9.697972e-06, 9.697961e-06, 9.697951e-06, 
    9.697953e-06, 9.697946e-06, 9.697966e-06, 9.697957e-06, 9.69796e-06, 
    9.697952e-06, 9.69797e-06, 9.697955e-06, 9.697975e-06, 9.697973e-06, 
    9.697967e-06, 9.697957e-06, 9.697954e-06, 9.697951e-06, 9.697953e-06, 
    9.697961e-06, 9.697962e-06, 9.697967e-06, 9.697969e-06, 9.697973e-06, 
    9.697977e-06, 9.697974e-06, 9.69797e-06, 9.697961e-06, 9.697952e-06, 
    9.697943e-06, 9.697941e-06, 9.69793e-06, 9.697938e-06, 9.697924e-06, 
    9.697937e-06, 9.697916e-06, 9.697954e-06, 9.697937e-06, 9.697967e-06, 
    9.697964e-06, 9.697958e-06, 9.697945e-06, 9.697952e-06, 9.697943e-06, 
    9.697962e-06, 9.697972e-06, 9.697975e-06, 9.697979e-06, 9.697975e-06, 
    9.697975e-06, 9.69797e-06, 9.697972e-06, 9.69796e-06, 9.697967e-06, 
    9.697949e-06, 9.697943e-06, 9.697926e-06, 9.697916e-06, 9.697905e-06, 
    9.697899e-06, 9.697898e-06, 9.697897e-06 ;

 LITR3C_TO_SOIL2C =
  6.006619e-14, 6.022866e-14, 6.019711e-14, 6.032803e-14, 6.025544e-14, 
    6.034113e-14, 6.009916e-14, 6.023509e-14, 6.014834e-14, 6.008085e-14, 
    6.058172e-14, 6.033387e-14, 6.083893e-14, 6.068116e-14, 6.107725e-14, 
    6.081437e-14, 6.113021e-14, 6.106973e-14, 6.125181e-14, 6.119968e-14, 
    6.143221e-14, 6.127587e-14, 6.155267e-14, 6.139491e-14, 6.141959e-14, 
    6.12707e-14, 6.038383e-14, 6.055087e-14, 6.037392e-14, 6.039775e-14, 
    6.038707e-14, 6.025691e-14, 6.019125e-14, 6.00538e-14, 6.007877e-14, 
    6.017974e-14, 6.040847e-14, 6.03309e-14, 6.052642e-14, 6.052201e-14, 
    6.073934e-14, 6.064139e-14, 6.100625e-14, 6.090265e-14, 6.120185e-14, 
    6.112666e-14, 6.119831e-14, 6.11766e-14, 6.119859e-14, 6.10883e-14, 
    6.113557e-14, 6.103849e-14, 6.065973e-14, 6.077113e-14, 6.043861e-14, 
    6.023823e-14, 6.010512e-14, 6.001055e-14, 6.002393e-14, 6.00494e-14, 
    6.018033e-14, 6.030337e-14, 6.039705e-14, 6.045968e-14, 6.052137e-14, 
    6.070781e-14, 6.08065e-14, 6.102716e-14, 6.098741e-14, 6.105478e-14, 
    6.111918e-14, 6.122717e-14, 6.120941e-14, 6.125695e-14, 6.105303e-14, 
    6.118858e-14, 6.096475e-14, 6.102599e-14, 6.053797e-14, 6.035184e-14, 
    6.027251e-14, 6.020316e-14, 6.00342e-14, 6.015089e-14, 6.01049e-14, 
    6.021434e-14, 6.028381e-14, 6.024946e-14, 6.046139e-14, 6.037903e-14, 
    6.081235e-14, 6.062586e-14, 6.111167e-14, 6.099557e-14, 6.113949e-14, 
    6.106607e-14, 6.119182e-14, 6.107866e-14, 6.127465e-14, 6.131728e-14, 
    6.128815e-14, 6.140007e-14, 6.107238e-14, 6.119829e-14, 6.024849e-14, 
    6.02541e-14, 6.02802e-14, 6.016538e-14, 6.015836e-14, 6.00531e-14, 
    6.014678e-14, 6.018664e-14, 6.028785e-14, 6.034766e-14, 6.040449e-14, 
    6.052939e-14, 6.066872e-14, 6.086338e-14, 6.10031e-14, 6.109668e-14, 
    6.103931e-14, 6.108995e-14, 6.103333e-14, 6.10068e-14, 6.13013e-14, 
    6.113599e-14, 6.138398e-14, 6.137027e-14, 6.125807e-14, 6.137182e-14, 
    6.025803e-14, 6.022578e-14, 6.011373e-14, 6.020143e-14, 6.004164e-14, 
    6.013108e-14, 6.018248e-14, 6.038072e-14, 6.042427e-14, 6.046461e-14, 
    6.054426e-14, 6.064641e-14, 6.082541e-14, 6.098101e-14, 6.112293e-14, 
    6.111254e-14, 6.11162e-14, 6.114786e-14, 6.106939e-14, 6.116075e-14, 
    6.117606e-14, 6.1136e-14, 6.136844e-14, 6.130207e-14, 6.136998e-14, 
    6.132678e-14, 6.023627e-14, 6.029052e-14, 6.026121e-14, 6.031632e-14, 
    6.027748e-14, 6.045006e-14, 6.050177e-14, 6.07435e-14, 6.064439e-14, 
    6.080215e-14, 6.066043e-14, 6.068555e-14, 6.080723e-14, 6.06681e-14, 
    6.09724e-14, 6.07661e-14, 6.11491e-14, 6.094327e-14, 6.116198e-14, 
    6.112232e-14, 6.1188e-14, 6.124678e-14, 6.132073e-14, 6.145701e-14, 
    6.142547e-14, 6.153939e-14, 6.037139e-14, 6.044167e-14, 6.043552e-14, 
    6.050907e-14, 6.056342e-14, 6.068122e-14, 6.086992e-14, 6.079899e-14, 
    6.09292e-14, 6.095532e-14, 6.075751e-14, 6.087896e-14, 6.048872e-14, 
    6.05518e-14, 6.051427e-14, 6.037692e-14, 6.08153e-14, 6.059046e-14, 
    6.10054e-14, 6.088381e-14, 6.123839e-14, 6.106212e-14, 6.140809e-14, 
    6.155565e-14, 6.169451e-14, 6.185644e-14, 6.048005e-14, 6.04323e-14, 
    6.051781e-14, 6.063599e-14, 6.074563e-14, 6.089122e-14, 6.090613e-14, 
    6.093338e-14, 6.100396e-14, 6.106328e-14, 6.094195e-14, 6.107814e-14, 
    6.056637e-14, 6.083481e-14, 6.041422e-14, 6.054095e-14, 6.062903e-14, 
    6.059044e-14, 6.07909e-14, 6.083809e-14, 6.102971e-14, 6.093071e-14, 
    6.151922e-14, 6.125914e-14, 6.197971e-14, 6.177871e-14, 6.041561e-14, 
    6.04799e-14, 6.07034e-14, 6.05971e-14, 6.090095e-14, 6.097563e-14, 
    6.103634e-14, 6.111385e-14, 6.112225e-14, 6.116815e-14, 6.109292e-14, 
    6.11652e-14, 6.089153e-14, 6.101389e-14, 6.06779e-14, 6.075973e-14, 
    6.07221e-14, 6.06808e-14, 6.080825e-14, 6.094386e-14, 6.094681e-14, 
    6.099025e-14, 6.111253e-14, 6.090218e-14, 6.155265e-14, 6.11512e-14, 
    6.054997e-14, 6.06736e-14, 6.069131e-14, 6.064343e-14, 6.096814e-14, 
    6.085056e-14, 6.116704e-14, 6.108159e-14, 6.122159e-14, 6.115203e-14, 
    6.11418e-14, 6.105241e-14, 6.099673e-14, 6.085595e-14, 6.074132e-14, 
    6.065038e-14, 6.067153e-14, 6.077141e-14, 6.095216e-14, 6.112298e-14, 
    6.108558e-14, 6.121095e-14, 6.087894e-14, 6.101823e-14, 6.096439e-14, 
    6.110473e-14, 6.07971e-14, 6.105895e-14, 6.073007e-14, 6.075895e-14, 
    6.084823e-14, 6.102763e-14, 6.106738e-14, 6.11097e-14, 6.108359e-14, 
    6.095675e-14, 6.093599e-14, 6.084608e-14, 6.082121e-14, 6.075267e-14, 
    6.069587e-14, 6.074775e-14, 6.080221e-14, 6.095683e-14, 6.109601e-14, 
    6.12476e-14, 6.12847e-14, 6.146144e-14, 6.131751e-14, 6.155487e-14, 
    6.1353e-14, 6.170232e-14, 6.107419e-14, 6.134715e-14, 6.085231e-14, 
    6.090571e-14, 6.100221e-14, 6.122338e-14, 6.110408e-14, 6.124362e-14, 
    6.093518e-14, 6.077483e-14, 6.073338e-14, 6.06559e-14, 6.073515e-14, 
    6.072871e-14, 6.08045e-14, 6.078015e-14, 6.096196e-14, 6.086433e-14, 
    6.114153e-14, 6.124253e-14, 6.152744e-14, 6.170177e-14, 6.187908e-14, 
    6.195725e-14, 6.198104e-14, 6.199098e-14 ;

 LITR3C_vr =
  0.0005537667, 0.0005537661, 0.0005537662, 0.0005537658, 0.000553766, 
    0.0005537657, 0.0005537666, 0.0005537661, 0.0005537664, 0.0005537666, 
    0.0005537649, 0.0005537657, 0.000553764, 0.0005537645, 0.0005537632, 
    0.0005537641, 0.000553763, 0.0005537632, 0.0005537625, 0.0005537627, 
    0.0005537619, 0.0005537625, 0.0005537615, 0.0005537621, 0.000553762, 
    0.0005537625, 0.0005537656, 0.000553765, 0.0005537656, 0.0005537655, 
    0.0005537656, 0.000553766, 0.0005537663, 0.0005537667, 0.0005537667, 
    0.0005537663, 0.0005537655, 0.0005537657, 0.0005537651, 0.0005537651, 
    0.0005537643, 0.0005537647, 0.0005537634, 0.0005537638, 0.0005537627, 
    0.000553763, 0.0005537627, 0.0005537628, 0.0005537627, 0.0005537631, 
    0.0005537629, 0.0005537633, 0.0005537646, 0.0005537642, 0.0005537654, 
    0.0005537661, 0.0005537666, 0.0005537669, 0.0005537668, 0.0005537667, 
    0.0005537663, 0.0005537659, 0.0005537656, 0.0005537653, 0.0005537651, 
    0.0005537645, 0.0005537641, 0.0005537634, 0.0005537635, 0.0005537632, 
    0.000553763, 0.0005537627, 0.0005537627, 0.0005537625, 0.0005537632, 
    0.0005537628, 0.0005537635, 0.0005537634, 0.000553765, 0.0005537657, 
    0.000553766, 0.0005537662, 0.0005537668, 0.0005537664, 0.0005537666, 
    0.0005537661, 0.0005537659, 0.000553766, 0.0005537653, 0.0005537656, 
    0.0005537641, 0.0005537648, 0.0005537631, 0.0005537635, 0.0005537629, 
    0.0005537632, 0.0005537628, 0.0005537632, 0.0005537625, 0.0005537623, 
    0.0005537624, 0.000553762, 0.0005537632, 0.0005537627, 0.000553766, 
    0.000553766, 0.000553766, 0.0005537663, 0.0005537664, 0.0005537667, 
    0.0005537664, 0.0005537663, 0.0005537659, 0.0005537657, 0.0005537655, 
    0.0005537651, 0.0005537646, 0.0005537639, 0.0005537634, 0.0005537631, 
    0.0005537633, 0.0005537631, 0.0005537633, 0.0005537634, 0.0005537624, 
    0.0005537629, 0.0005537621, 0.0005537621, 0.0005537625, 0.0005537621, 
    0.000553766, 0.0005537661, 0.0005537665, 0.0005537662, 0.0005537668, 
    0.0005537664, 0.0005537663, 0.0005537656, 0.0005537655, 0.0005537653, 
    0.000553765, 0.0005537647, 0.0005537641, 0.0005537635, 0.000553763, 
    0.0005537631, 0.000553763, 0.0005537629, 0.0005537632, 0.0005537629, 
    0.0005537628, 0.0005537629, 0.0005537621, 0.0005537624, 0.0005537621, 
    0.0005537623, 0.0005537661, 0.0005537659, 0.000553766, 0.0005537658, 
    0.000553766, 0.0005537653, 0.0005537652, 0.0005537643, 0.0005537647, 
    0.0005537641, 0.0005537646, 0.0005537645, 0.0005537641, 0.0005537646, 
    0.0005537635, 0.0005537642, 0.0005537629, 0.0005537636, 0.0005537629, 
    0.000553763, 0.0005537628, 0.0005537626, 0.0005537623, 0.0005537618, 
    0.000553762, 0.0005537616, 0.0005537656, 0.0005537654, 0.0005537654, 
    0.0005537652, 0.000553765, 0.0005537645, 0.0005537639, 0.0005537641, 
    0.0005537637, 0.0005537636, 0.0005537643, 0.0005537639, 0.0005537652, 
    0.000553765, 0.0005537651, 0.0005537656, 0.0005537641, 0.0005537649, 
    0.0005537634, 0.0005537638, 0.0005537626, 0.0005537632, 0.000553762, 
    0.0005537615, 0.000553761, 0.0005537604, 0.0005537653, 0.0005537654, 
    0.0005537651, 0.0005537647, 0.0005537643, 0.0005537638, 0.0005537638, 
    0.0005537636, 0.0005537634, 0.0005537632, 0.0005537636, 0.0005537632, 
    0.0005537649, 0.000553764, 0.0005537655, 0.000553765, 0.0005537648, 
    0.0005537649, 0.0005537642, 0.000553764, 0.0005537634, 0.0005537637, 
    0.0005537616, 0.0005537625, 0.00055376, 0.0005537607, 0.0005537655, 
    0.0005537653, 0.0005537645, 0.0005537649, 0.0005537638, 0.0005537635, 
    0.0005537633, 0.0005537631, 0.000553763, 0.0005537628, 0.0005537631, 
    0.0005537628, 0.0005537638, 0.0005537634, 0.0005537646, 0.0005537643, 
    0.0005537644, 0.0005537645, 0.0005537641, 0.0005537636, 0.0005537636, 
    0.0005537635, 0.0005537631, 0.0005537638, 0.0005537615, 0.0005537629, 
    0.000553765, 0.0005537646, 0.0005537645, 0.0005537647, 0.0005537635, 
    0.0005537639, 0.0005537628, 0.0005537631, 0.0005537627, 0.0005537629, 
    0.0005537629, 0.0005537632, 0.0005537635, 0.0005537639, 0.0005537643, 
    0.0005537646, 0.0005537646, 0.0005537642, 0.0005537636, 0.000553763, 
    0.0005537631, 0.0005537627, 0.0005537639, 0.0005537634, 0.0005537635, 
    0.0005537631, 0.0005537642, 0.0005537632, 0.0005537644, 0.0005537643, 
    0.0005537639, 0.0005537634, 0.0005537632, 0.0005537631, 0.0005537631, 
    0.0005537636, 0.0005537636, 0.000553764, 0.0005537641, 0.0005537643, 
    0.0005537645, 0.0005537643, 0.0005537641, 0.0005537636, 0.0005537631, 
    0.0005537626, 0.0005537624, 0.0005537618, 0.0005537623, 0.0005537615, 
    0.0005537622, 0.000553761, 0.0005537632, 0.0005537622, 0.0005537639, 
    0.0005537638, 0.0005537634, 0.0005537627, 0.0005537631, 0.0005537626, 
    0.0005537636, 0.0005537642, 0.0005537643, 0.0005537646, 0.0005537643, 
    0.0005537644, 0.0005537641, 0.0005537642, 0.0005537636, 0.0005537639, 
    0.0005537629, 0.0005537626, 0.0005537616, 0.000553761, 0.0005537604, 
    0.0005537601, 0.00055376, 0.00055376,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342134e-07, 1.342133e-07, 1.342133e-07, 1.342132e-07, 1.342133e-07, 
    1.342132e-07, 1.342134e-07, 1.342133e-07, 1.342134e-07, 1.342134e-07, 
    1.34213e-07, 1.342132e-07, 1.342128e-07, 1.342129e-07, 1.342126e-07, 
    1.342128e-07, 1.342125e-07, 1.342126e-07, 1.342124e-07, 1.342125e-07, 
    1.342123e-07, 1.342124e-07, 1.342122e-07, 1.342123e-07, 1.342123e-07, 
    1.342124e-07, 1.342132e-07, 1.34213e-07, 1.342132e-07, 1.342132e-07, 
    1.342132e-07, 1.342133e-07, 1.342133e-07, 1.342135e-07, 1.342134e-07, 
    1.342133e-07, 1.342131e-07, 1.342132e-07, 1.34213e-07, 1.342131e-07, 
    1.342129e-07, 1.34213e-07, 1.342126e-07, 1.342127e-07, 1.342125e-07, 
    1.342125e-07, 1.342125e-07, 1.342125e-07, 1.342125e-07, 1.342126e-07, 
    1.342125e-07, 1.342126e-07, 1.342129e-07, 1.342128e-07, 1.342131e-07, 
    1.342133e-07, 1.342134e-07, 1.342135e-07, 1.342135e-07, 1.342135e-07, 
    1.342133e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342131e-07, 
    1.342129e-07, 1.342128e-07, 1.342126e-07, 1.342127e-07, 1.342126e-07, 
    1.342125e-07, 1.342125e-07, 1.342125e-07, 1.342124e-07, 1.342126e-07, 
    1.342125e-07, 1.342127e-07, 1.342126e-07, 1.34213e-07, 1.342132e-07, 
    1.342133e-07, 1.342133e-07, 1.342135e-07, 1.342134e-07, 1.342134e-07, 
    1.342133e-07, 1.342133e-07, 1.342133e-07, 1.342131e-07, 1.342132e-07, 
    1.342128e-07, 1.34213e-07, 1.342126e-07, 1.342126e-07, 1.342125e-07, 
    1.342126e-07, 1.342125e-07, 1.342126e-07, 1.342124e-07, 1.342124e-07, 
    1.342124e-07, 1.342123e-07, 1.342126e-07, 1.342125e-07, 1.342133e-07, 
    1.342133e-07, 1.342133e-07, 1.342134e-07, 1.342134e-07, 1.342135e-07, 
    1.342134e-07, 1.342133e-07, 1.342133e-07, 1.342132e-07, 1.342132e-07, 
    1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342126e-07, 1.342126e-07, 
    1.342126e-07, 1.342126e-07, 1.342126e-07, 1.342126e-07, 1.342124e-07, 
    1.342125e-07, 1.342123e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342133e-07, 1.342133e-07, 1.342134e-07, 1.342133e-07, 1.342135e-07, 
    1.342134e-07, 1.342133e-07, 1.342132e-07, 1.342131e-07, 1.342131e-07, 
    1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342127e-07, 1.342125e-07, 
    1.342126e-07, 1.342125e-07, 1.342125e-07, 1.342126e-07, 1.342125e-07, 
    1.342125e-07, 1.342125e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342124e-07, 1.342133e-07, 1.342133e-07, 1.342133e-07, 1.342132e-07, 
    1.342133e-07, 1.342131e-07, 1.342131e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342129e-07, 1.342129e-07, 1.342128e-07, 1.342129e-07, 
    1.342127e-07, 1.342128e-07, 1.342125e-07, 1.342127e-07, 1.342125e-07, 
    1.342125e-07, 1.342125e-07, 1.342124e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342132e-07, 1.342131e-07, 1.342131e-07, 
    1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342128e-07, 
    1.342127e-07, 1.342127e-07, 1.342129e-07, 1.342127e-07, 1.342131e-07, 
    1.34213e-07, 1.342131e-07, 1.342132e-07, 1.342128e-07, 1.34213e-07, 
    1.342126e-07, 1.342127e-07, 1.342124e-07, 1.342126e-07, 1.342123e-07, 
    1.342122e-07, 1.342121e-07, 1.342119e-07, 1.342131e-07, 1.342131e-07, 
    1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342127e-07, 1.342127e-07, 
    1.342127e-07, 1.342126e-07, 1.342126e-07, 1.342127e-07, 1.342126e-07, 
    1.34213e-07, 1.342128e-07, 1.342131e-07, 1.34213e-07, 1.34213e-07, 
    1.34213e-07, 1.342128e-07, 1.342128e-07, 1.342126e-07, 1.342127e-07, 
    1.342122e-07, 1.342124e-07, 1.342118e-07, 1.34212e-07, 1.342131e-07, 
    1.342131e-07, 1.342129e-07, 1.34213e-07, 1.342127e-07, 1.342127e-07, 
    1.342126e-07, 1.342125e-07, 1.342125e-07, 1.342125e-07, 1.342126e-07, 
    1.342125e-07, 1.342127e-07, 1.342126e-07, 1.342129e-07, 1.342129e-07, 
    1.342129e-07, 1.342129e-07, 1.342128e-07, 1.342127e-07, 1.342127e-07, 
    1.342127e-07, 1.342126e-07, 1.342127e-07, 1.342122e-07, 1.342125e-07, 
    1.34213e-07, 1.342129e-07, 1.342129e-07, 1.342129e-07, 1.342127e-07, 
    1.342128e-07, 1.342125e-07, 1.342126e-07, 1.342125e-07, 1.342125e-07, 
    1.342125e-07, 1.342126e-07, 1.342126e-07, 1.342128e-07, 1.342129e-07, 
    1.342129e-07, 1.342129e-07, 1.342128e-07, 1.342127e-07, 1.342125e-07, 
    1.342126e-07, 1.342125e-07, 1.342127e-07, 1.342126e-07, 1.342127e-07, 
    1.342126e-07, 1.342128e-07, 1.342126e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342126e-07, 1.342126e-07, 1.342126e-07, 1.342126e-07, 
    1.342127e-07, 1.342127e-07, 1.342128e-07, 1.342128e-07, 1.342129e-07, 
    1.342129e-07, 1.342129e-07, 1.342128e-07, 1.342127e-07, 1.342126e-07, 
    1.342124e-07, 1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342122e-07, 
    1.342123e-07, 1.34212e-07, 1.342126e-07, 1.342124e-07, 1.342128e-07, 
    1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342126e-07, 1.342124e-07, 
    1.342127e-07, 1.342128e-07, 1.342129e-07, 1.342129e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.342128e-07, 1.342127e-07, 1.342128e-07, 
    1.342125e-07, 1.342124e-07, 1.342122e-07, 1.34212e-07, 1.342119e-07, 
    1.342118e-07, 1.342118e-07, 1.342118e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  -6.617445e-26, -5.882173e-26, -9.190896e-26, 6.4949e-26, 1.789161e-25, 
    -9.803622e-26, -5.391992e-26, -2.205815e-26, 2.32836e-26, 8.578169e-27, 
    7.352717e-26, 3.431268e-26, -1.838179e-26, 1.274471e-25, 9.803622e-27, 
    1.225453e-26, -1.347998e-26, -4.779266e-26, -4.901811e-27, -1.384762e-25, 
    -1.225453e-27, -7.475262e-26, -1.200944e-25, -6.127264e-26, 4.901811e-26, 
    6.127264e-26, 3.063632e-26, 9.803622e-27, 4.166539e-26, 9.068351e-26, 
    2.08327e-26, 4.166539e-26, -2.941087e-26, -4.901811e-27, -2.450906e-27, 
    -4.779266e-26, 7.352717e-27, 1.347998e-25, -3.798904e-26, -4.901811e-27, 
    6.73999e-26, -7.352717e-26, -3.921449e-26, 6.862535e-26, 4.289085e-26, 
    5.637083e-26, 1.225453e-27, -5.024356e-26, 1.225453e-26, 1.593089e-26, 
    4.41163e-26, 2.695996e-26, -3.186177e-26, 7.352717e-26, -1.102908e-26, 
    -1.470543e-26, 9.803622e-27, -6.127264e-26, -2.573451e-26, 0, 
    1.102908e-25, -6.98508e-26, -1.066144e-25, 7.720352e-26, -1.642107e-25, 
    6.73999e-26, 1.102908e-26, 5.882173e-26, -1.176435e-25, -4.901811e-26, 
    2.450905e-26, 6.004719e-26, -7.652491e-42, 3.308722e-26, -6.4949e-26, 
    2.450905e-26, 1.225453e-27, 7.720352e-26, 5.024356e-26, 9.068351e-26, 
    9.803622e-27, 4.166539e-26, -7.352717e-27, 7.107626e-26, 2.32836e-26, 
    2.120033e-25, 7.230172e-26, -2.450906e-27, -1.225453e-26, 6.372354e-26, 
    -3.553813e-26, -2.450905e-26, -3.921449e-26, -4.534175e-26, 
    -9.803622e-27, -2.08327e-26, 4.41163e-26, 6.98508e-26, 6.4949e-26, 
    -3.676358e-26, -3.063632e-26, -1.225453e-26, 5.391992e-26, -3.186177e-26, 
    3.921449e-26, 1.225453e-27, 2.818541e-26, -1.384762e-25, -6.249809e-26, 
    -1.593089e-26, -3.431268e-26, 3.431268e-26, 4.166539e-26, -4.901811e-27, 
    1.311234e-25, 3.063632e-26, -9.558531e-26, -4.289085e-26, -4.166539e-26, 
    2.254833e-25, 2.450905e-26, 1.225453e-27, 8.945805e-26, -3.186177e-26, 
    -1.225453e-26, -6.4949e-26, -2.205815e-26, 1.81367e-25, -1.715634e-26, 
    -5.514538e-26, -2.573451e-26, 5.514538e-26, 2.450906e-27, -5.269447e-26, 
    -1.127417e-25, 2.08327e-26, -6.127264e-27, -6.004719e-26, 8.700715e-26, 
    2.08327e-26, 5.759628e-26, 9.803622e-26, -6.4949e-26, -1.139671e-25, 
    -6.98508e-26, -3.186177e-26, -3.308722e-26, 1.850434e-25, -3.431268e-26, 
    1.102908e-26, 1.593089e-26, 7.352717e-27, 2.32836e-26, -1.090653e-25, 
    1.078398e-25, -4.779266e-26, -2.573451e-26, -1.740143e-25, 9.435986e-26, 
    1.200944e-25, 1.225453e-26, 3.676358e-26, -7.597807e-26, 2.08327e-26, 
    3.798904e-26, 1.225453e-27, -9.558531e-26, 1.347998e-26, -6.98508e-26, 
    -1.838179e-26, 3.553813e-26, 2.205815e-26, 1.397016e-25, -6.862535e-26, 
    5.637083e-26, -1.102908e-26, 6.004719e-26, 4.41163e-26, 1.078398e-25, 
    -6.98508e-26, -2.695996e-26, -9.926167e-26, -8.578169e-27, -3.431268e-26, 
    -6.73999e-26, 3.921449e-26, -3.553813e-26, -9.681077e-26, -4.779266e-26, 
    8.578169e-26, 2.32836e-26, -5.514538e-26, 6.862535e-26, 2.695996e-26, 
    1.102908e-26, -6.4949e-26, 7.720352e-26, -4.779266e-26, 3.553813e-26, 
    7.352717e-27, -7.965443e-26, 1.838179e-26, -2.695996e-26, 2.450905e-26, 
    -1.053889e-25, -1.715634e-26, -1.225453e-27, -2.32836e-26, -3.063632e-26, 
    -3.553813e-26, 1.066144e-25, -4.65672e-26, -3.063632e-26, 6.862535e-26, 
    1.372507e-25, -6.127264e-27, 6.127264e-27, -2.450906e-27, -2.08327e-26, 
    2.818541e-26, 9.681077e-26, -2.205815e-26, -4.65672e-26, 3.186177e-26, 
    -2.695996e-26, 1.470543e-25, 4.901811e-26, -1.139671e-25, 6.249809e-26, 
    -2.32836e-26, 8.210533e-26, -1.225453e-27, 2.450905e-26, -4.043994e-26, 
    -7.107626e-26, -1.960724e-26, -2.205815e-26, 2.08327e-26, -2.573451e-26, 
    9.803622e-27, 1.090653e-25, -8.578169e-26, 1.115162e-25, -4.289085e-26, 
    1.004871e-25, -1.838179e-26, 4.779266e-26, -3.431268e-26, -6.372354e-26, 
    -4.043994e-26, 1.151926e-25, 1.715634e-26, 9.803622e-26, 8.82326e-26, 
    -9.068351e-26, -6.249809e-26, -9.435986e-26, 2.941087e-26, -1.347998e-25, 
    1.347998e-26, 4.65672e-26, -4.534175e-26, -9.435986e-26, -9.803622e-27, 
    5.514538e-26, -1.225453e-26, 5.024356e-26, 1.213198e-25, 6.617445e-26, 
    -1.470543e-26, -5.391992e-26, 4.779266e-26, -9.803622e-26, 6.127264e-27, 
    -1.960724e-26, -1.041635e-25, 6.98508e-26, -1.580834e-25, -3.921449e-26, 
    -1.017126e-25, 2.205815e-26, -7.597807e-26, 8.455624e-26, -5.514538e-26, 
    2.573451e-26, 6.372354e-26, 5.882173e-26, -8.578169e-26, 9.926167e-26, 
    -2.450906e-27, 5.882173e-26, -8.333079e-26, -7.230172e-26, 7.107626e-26, 
    7.965443e-26, 1.67887e-25, -9.803622e-27, -4.289085e-26, 1.715634e-26, 
    6.004719e-26, -1.960724e-26, -7.720352e-26, 8.578169e-27, -8.578169e-27, 
    4.65672e-26, -3.676358e-27, 7.352717e-27, -5.391992e-26, 1.593089e-26, 
    9.803622e-27, -1.02938e-25, -1.397016e-25, 3.063632e-26, 2.818541e-26, 
    -3.676358e-26, -6.4949e-26, 2.450906e-27, -8.087988e-26, 4.166539e-26, 
    -3.553813e-26, 5.146902e-26, -1.531816e-25, -3.676358e-26, 6.249809e-26, 
    7.230172e-26, 7.107626e-26, 1.593089e-26, -1.593089e-26, 9.190896e-26, 
    1.225453e-27, 3.186177e-26, 2.695996e-26, -7.720352e-26, -2.941087e-26, 
    2.08327e-26, 8.578169e-26, 2.573451e-26, 3.676358e-26,
  1.338128e-32, 1.338126e-32, 1.338126e-32, 1.338125e-32, 1.338126e-32, 
    1.338125e-32, 1.338127e-32, 1.338126e-32, 1.338127e-32, 1.338127e-32, 
    1.338123e-32, 1.338125e-32, 1.338121e-32, 1.338122e-32, 1.338119e-32, 
    1.338121e-32, 1.338118e-32, 1.338119e-32, 1.338117e-32, 1.338118e-32, 
    1.338116e-32, 1.338117e-32, 1.338115e-32, 1.338116e-32, 1.338116e-32, 
    1.338117e-32, 1.338125e-32, 1.338123e-32, 1.338125e-32, 1.338125e-32, 
    1.338125e-32, 1.338126e-32, 1.338126e-32, 1.338128e-32, 1.338127e-32, 
    1.338126e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338124e-32, 
    1.338122e-32, 1.338123e-32, 1.338119e-32, 1.33812e-32, 1.338118e-32, 
    1.338118e-32, 1.338118e-32, 1.338118e-32, 1.338118e-32, 1.338119e-32, 
    1.338118e-32, 1.338119e-32, 1.338122e-32, 1.338121e-32, 1.338124e-32, 
    1.338126e-32, 1.338127e-32, 1.338128e-32, 1.338128e-32, 1.338128e-32, 
    1.338126e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338124e-32, 
    1.338122e-32, 1.338121e-32, 1.338119e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338118e-32, 1.338118e-32, 1.338117e-32, 1.338119e-32, 
    1.338118e-32, 1.33812e-32, 1.338119e-32, 1.338123e-32, 1.338125e-32, 
    1.338126e-32, 1.338126e-32, 1.338128e-32, 1.338127e-32, 1.338127e-32, 
    1.338126e-32, 1.338126e-32, 1.338126e-32, 1.338124e-32, 1.338125e-32, 
    1.338121e-32, 1.338123e-32, 1.338119e-32, 1.33812e-32, 1.338118e-32, 
    1.338119e-32, 1.338118e-32, 1.338119e-32, 1.338117e-32, 1.338117e-32, 
    1.338117e-32, 1.338116e-32, 1.338119e-32, 1.338118e-32, 1.338126e-32, 
    1.338126e-32, 1.338126e-32, 1.338127e-32, 1.338127e-32, 1.338128e-32, 
    1.338127e-32, 1.338126e-32, 1.338126e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338122e-32, 1.338121e-32, 1.338119e-32, 1.338119e-32, 
    1.338119e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 1.338117e-32, 
    1.338118e-32, 1.338116e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 
    1.338126e-32, 1.338126e-32, 1.338127e-32, 1.338126e-32, 1.338128e-32, 
    1.338127e-32, 1.338126e-32, 1.338125e-32, 1.338124e-32, 1.338124e-32, 
    1.338123e-32, 1.338123e-32, 1.338121e-32, 1.33812e-32, 1.338118e-32, 
    1.338119e-32, 1.338119e-32, 1.338118e-32, 1.338119e-32, 1.338118e-32, 
    1.338118e-32, 1.338118e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 
    1.338117e-32, 1.338126e-32, 1.338126e-32, 1.338126e-32, 1.338125e-32, 
    1.338126e-32, 1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338123e-32, 
    1.338121e-32, 1.338122e-32, 1.338122e-32, 1.338121e-32, 1.338122e-32, 
    1.33812e-32, 1.338121e-32, 1.338118e-32, 1.33812e-32, 1.338118e-32, 
    1.338118e-32, 1.338118e-32, 1.338117e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338115e-32, 1.338125e-32, 1.338124e-32, 1.338124e-32, 
    1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 1.338121e-32, 
    1.33812e-32, 1.33812e-32, 1.338122e-32, 1.338121e-32, 1.338124e-32, 
    1.338123e-32, 1.338124e-32, 1.338125e-32, 1.338121e-32, 1.338123e-32, 
    1.338119e-32, 1.33812e-32, 1.338118e-32, 1.338119e-32, 1.338116e-32, 
    1.338115e-32, 1.338114e-32, 1.338112e-32, 1.338124e-32, 1.338124e-32, 
    1.338124e-32, 1.338123e-32, 1.338122e-32, 1.33812e-32, 1.33812e-32, 
    1.33812e-32, 1.338119e-32, 1.338119e-32, 1.33812e-32, 1.338119e-32, 
    1.338123e-32, 1.338121e-32, 1.338124e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338121e-32, 1.338121e-32, 1.338119e-32, 1.33812e-32, 
    1.338115e-32, 1.338117e-32, 1.338111e-32, 1.338113e-32, 1.338124e-32, 
    1.338124e-32, 1.338122e-32, 1.338123e-32, 1.33812e-32, 1.33812e-32, 
    1.338119e-32, 1.338119e-32, 1.338119e-32, 1.338118e-32, 1.338119e-32, 
    1.338118e-32, 1.33812e-32, 1.338119e-32, 1.338122e-32, 1.338121e-32, 
    1.338122e-32, 1.338122e-32, 1.338121e-32, 1.33812e-32, 1.33812e-32, 
    1.33812e-32, 1.338119e-32, 1.33812e-32, 1.338115e-32, 1.338118e-32, 
    1.338123e-32, 1.338122e-32, 1.338122e-32, 1.338123e-32, 1.33812e-32, 
    1.338121e-32, 1.338118e-32, 1.338119e-32, 1.338118e-32, 1.338118e-32, 
    1.338118e-32, 1.338119e-32, 1.33812e-32, 1.338121e-32, 1.338122e-32, 
    1.338123e-32, 1.338122e-32, 1.338121e-32, 1.33812e-32, 1.338118e-32, 
    1.338119e-32, 1.338118e-32, 1.338121e-32, 1.338119e-32, 1.33812e-32, 
    1.338119e-32, 1.338121e-32, 1.338119e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 
    1.33812e-32, 1.33812e-32, 1.338121e-32, 1.338121e-32, 1.338122e-32, 
    1.338122e-32, 1.338122e-32, 1.338121e-32, 1.33812e-32, 1.338119e-32, 
    1.338117e-32, 1.338117e-32, 1.338116e-32, 1.338117e-32, 1.338115e-32, 
    1.338117e-32, 1.338114e-32, 1.338119e-32, 1.338117e-32, 1.338121e-32, 
    1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338119e-32, 1.338117e-32, 
    1.33812e-32, 1.338121e-32, 1.338122e-32, 1.338123e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.338121e-32, 1.33812e-32, 1.338121e-32, 
    1.338118e-32, 1.338118e-32, 1.338115e-32, 1.338114e-32, 1.338112e-32, 
    1.338111e-32, 1.338111e-32, 1.338111e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.662544e-15, 1.667041e-15, 1.666168e-15, 1.669792e-15, 1.667782e-15, 
    1.670154e-15, 1.663457e-15, 1.667219e-15, 1.664818e-15, 1.66295e-15, 
    1.676813e-15, 1.669953e-15, 1.683933e-15, 1.679566e-15, 1.690529e-15, 
    1.683253e-15, 1.691995e-15, 1.690321e-15, 1.69536e-15, 1.693917e-15, 
    1.700354e-15, 1.696026e-15, 1.703688e-15, 1.699321e-15, 1.700004e-15, 
    1.695883e-15, 1.671336e-15, 1.675959e-15, 1.671062e-15, 1.671721e-15, 
    1.671426e-15, 1.667823e-15, 1.666006e-15, 1.662201e-15, 1.662892e-15, 
    1.665687e-15, 1.672018e-15, 1.669871e-15, 1.675283e-15, 1.675161e-15, 
    1.681176e-15, 1.678465e-15, 1.688564e-15, 1.685696e-15, 1.693978e-15, 
    1.691896e-15, 1.69388e-15, 1.693279e-15, 1.693887e-15, 1.690835e-15, 
    1.692143e-15, 1.689456e-15, 1.678973e-15, 1.682056e-15, 1.672852e-15, 
    1.667306e-15, 1.663622e-15, 1.661004e-15, 1.661374e-15, 1.66208e-15, 
    1.665704e-15, 1.669109e-15, 1.671702e-15, 1.673436e-15, 1.675143e-15, 
    1.680303e-15, 1.683035e-15, 1.689143e-15, 1.688042e-15, 1.689907e-15, 
    1.691689e-15, 1.694678e-15, 1.694187e-15, 1.695503e-15, 1.689859e-15, 
    1.69361e-15, 1.687415e-15, 1.68911e-15, 1.675602e-15, 1.670451e-15, 
    1.668255e-15, 1.666336e-15, 1.661659e-15, 1.664889e-15, 1.663616e-15, 
    1.666645e-15, 1.668568e-15, 1.667617e-15, 1.673483e-15, 1.671203e-15, 
    1.683197e-15, 1.678035e-15, 1.691482e-15, 1.688268e-15, 1.692252e-15, 
    1.69022e-15, 1.6937e-15, 1.690568e-15, 1.695993e-15, 1.697173e-15, 
    1.696366e-15, 1.699464e-15, 1.690394e-15, 1.693879e-15, 1.66759e-15, 
    1.667745e-15, 1.668468e-15, 1.66529e-15, 1.665095e-15, 1.662182e-15, 
    1.664775e-15, 1.665878e-15, 1.668679e-15, 1.670335e-15, 1.671908e-15, 
    1.675365e-15, 1.679221e-15, 1.684609e-15, 1.688476e-15, 1.691067e-15, 
    1.689479e-15, 1.690881e-15, 1.689313e-15, 1.688579e-15, 1.69673e-15, 
    1.692155e-15, 1.699019e-15, 1.698639e-15, 1.695534e-15, 1.698682e-15, 
    1.667854e-15, 1.666962e-15, 1.66386e-15, 1.666288e-15, 1.661865e-15, 
    1.66434e-15, 1.665763e-15, 1.67125e-15, 1.672456e-15, 1.673572e-15, 
    1.675777e-15, 1.678604e-15, 1.683558e-15, 1.687865e-15, 1.691793e-15, 
    1.691506e-15, 1.691607e-15, 1.692483e-15, 1.690311e-15, 1.69284e-15, 
    1.693264e-15, 1.692155e-15, 1.698589e-15, 1.696752e-15, 1.698631e-15, 
    1.697436e-15, 1.667252e-15, 1.668753e-15, 1.667942e-15, 1.669468e-15, 
    1.668393e-15, 1.673169e-15, 1.6746e-15, 1.681291e-15, 1.678548e-15, 
    1.682915e-15, 1.678992e-15, 1.679687e-15, 1.683055e-15, 1.679204e-15, 
    1.687627e-15, 1.681917e-15, 1.692518e-15, 1.68682e-15, 1.692874e-15, 
    1.691776e-15, 1.693594e-15, 1.695221e-15, 1.697268e-15, 1.70104e-15, 
    1.700167e-15, 1.70332e-15, 1.670992e-15, 1.672937e-15, 1.672767e-15, 
    1.674802e-15, 1.676307e-15, 1.679567e-15, 1.68479e-15, 1.682827e-15, 
    1.686431e-15, 1.687154e-15, 1.681679e-15, 1.685041e-15, 1.674239e-15, 
    1.675985e-15, 1.674946e-15, 1.671145e-15, 1.683279e-15, 1.677055e-15, 
    1.68854e-15, 1.685175e-15, 1.694989e-15, 1.69011e-15, 1.699686e-15, 
    1.70377e-15, 1.707614e-15, 1.712096e-15, 1.673999e-15, 1.672678e-15, 
    1.675045e-15, 1.678315e-15, 1.68135e-15, 1.68538e-15, 1.685792e-15, 
    1.686547e-15, 1.6885e-15, 1.690142e-15, 1.686784e-15, 1.690554e-15, 
    1.676388e-15, 1.683819e-15, 1.672177e-15, 1.675685e-15, 1.678123e-15, 
    1.677055e-15, 1.682603e-15, 1.683909e-15, 1.689213e-15, 1.686473e-15, 
    1.702762e-15, 1.695563e-15, 1.715508e-15, 1.709944e-15, 1.672216e-15, 
    1.673995e-15, 1.680181e-15, 1.677239e-15, 1.685649e-15, 1.687716e-15, 
    1.689397e-15, 1.691542e-15, 1.691774e-15, 1.693045e-15, 1.690962e-15, 
    1.692963e-15, 1.685388e-15, 1.688775e-15, 1.679476e-15, 1.681741e-15, 
    1.680699e-15, 1.679556e-15, 1.683083e-15, 1.686837e-15, 1.686918e-15, 
    1.688121e-15, 1.691505e-15, 1.685683e-15, 1.703687e-15, 1.692576e-15, 
    1.675935e-15, 1.679357e-15, 1.679847e-15, 1.678521e-15, 1.687509e-15, 
    1.684255e-15, 1.693014e-15, 1.690649e-15, 1.694524e-15, 1.692599e-15, 
    1.692316e-15, 1.689842e-15, 1.6883e-15, 1.684404e-15, 1.681231e-15, 
    1.678714e-15, 1.679299e-15, 1.682064e-15, 1.687067e-15, 1.691795e-15, 
    1.690759e-15, 1.69423e-15, 1.68504e-15, 1.688895e-15, 1.687405e-15, 
    1.69129e-15, 1.682775e-15, 1.690022e-15, 1.68092e-15, 1.681719e-15, 
    1.68419e-15, 1.689156e-15, 1.690256e-15, 1.691427e-15, 1.690705e-15, 
    1.687194e-15, 1.686619e-15, 1.68413e-15, 1.683442e-15, 1.681545e-15, 
    1.679973e-15, 1.681409e-15, 1.682916e-15, 1.687196e-15, 1.691048e-15, 
    1.695244e-15, 1.696271e-15, 1.701163e-15, 1.697179e-15, 1.703749e-15, 
    1.698161e-15, 1.70783e-15, 1.690444e-15, 1.698e-15, 1.684303e-15, 
    1.685781e-15, 1.688452e-15, 1.694574e-15, 1.691271e-15, 1.695134e-15, 
    1.686597e-15, 1.682158e-15, 1.681011e-15, 1.678867e-15, 1.68106e-15, 
    1.680882e-15, 1.68298e-15, 1.682306e-15, 1.687338e-15, 1.684636e-15, 
    1.692308e-15, 1.695104e-15, 1.702989e-15, 1.707815e-15, 1.712722e-15, 
    1.714886e-15, 1.715544e-15, 1.71582e-15 ;

 LITR3N_vr =
  7.663726e-06, 7.663718e-06, 7.66372e-06, 7.663713e-06, 7.663717e-06, 
    7.663712e-06, 7.663724e-06, 7.663718e-06, 7.663722e-06, 7.663725e-06, 
    7.663701e-06, 7.663712e-06, 7.663689e-06, 7.663696e-06, 7.663677e-06, 
    7.66369e-06, 7.663674e-06, 7.663677e-06, 7.663669e-06, 7.663671e-06, 
    7.66366e-06, 7.663667e-06, 7.663654e-06, 7.663662e-06, 7.663661e-06, 
    7.663668e-06, 7.663711e-06, 7.663702e-06, 7.663711e-06, 7.66371e-06, 
    7.663711e-06, 7.663717e-06, 7.66372e-06, 7.663726e-06, 7.663725e-06, 
    7.663721e-06, 7.663709e-06, 7.663713e-06, 7.663703e-06, 7.663703e-06, 
    7.663693e-06, 7.663698e-06, 7.663681e-06, 7.663685e-06, 7.663671e-06, 
    7.663674e-06, 7.663671e-06, 7.663672e-06, 7.663671e-06, 7.663676e-06, 
    7.663674e-06, 7.663679e-06, 7.663697e-06, 7.663692e-06, 7.663708e-06, 
    7.663718e-06, 7.663724e-06, 7.663729e-06, 7.663728e-06, 7.663727e-06, 
    7.663721e-06, 7.663714e-06, 7.66371e-06, 7.663707e-06, 7.663703e-06, 
    7.663695e-06, 7.66369e-06, 7.66368e-06, 7.663682e-06, 7.663678e-06, 
    7.663675e-06, 7.66367e-06, 7.663671e-06, 7.663668e-06, 7.663678e-06, 
    7.663672e-06, 7.663682e-06, 7.66368e-06, 7.663703e-06, 7.663712e-06, 
    7.663716e-06, 7.663719e-06, 7.663727e-06, 7.663722e-06, 7.663724e-06, 
    7.663719e-06, 7.663715e-06, 7.663717e-06, 7.663707e-06, 7.663711e-06, 
    7.66369e-06, 7.663699e-06, 7.663675e-06, 7.663681e-06, 7.663674e-06, 
    7.663678e-06, 7.663672e-06, 7.663677e-06, 7.663667e-06, 7.663665e-06, 
    7.663667e-06, 7.663662e-06, 7.663677e-06, 7.663671e-06, 7.663717e-06, 
    7.663717e-06, 7.663715e-06, 7.663721e-06, 7.663722e-06, 7.663726e-06, 
    7.663722e-06, 7.66372e-06, 7.663715e-06, 7.663712e-06, 7.66371e-06, 
    7.663703e-06, 7.663697e-06, 7.663687e-06, 7.663681e-06, 7.663676e-06, 
    7.663679e-06, 7.663676e-06, 7.663679e-06, 7.663681e-06, 7.663666e-06, 
    7.663674e-06, 7.663662e-06, 7.663662e-06, 7.663668e-06, 7.663662e-06, 
    7.663716e-06, 7.663718e-06, 7.663723e-06, 7.663719e-06, 7.663727e-06, 
    7.663722e-06, 7.66372e-06, 7.663711e-06, 7.663709e-06, 7.663706e-06, 
    7.663702e-06, 7.663698e-06, 7.663689e-06, 7.663682e-06, 7.663674e-06, 
    7.663675e-06, 7.663675e-06, 7.663673e-06, 7.663677e-06, 7.663672e-06, 
    7.663672e-06, 7.663674e-06, 7.663662e-06, 7.663666e-06, 7.663662e-06, 
    7.663665e-06, 7.663718e-06, 7.663715e-06, 7.663716e-06, 7.663713e-06, 
    7.663715e-06, 7.663707e-06, 7.663705e-06, 7.663693e-06, 7.663698e-06, 
    7.663691e-06, 7.663697e-06, 7.663696e-06, 7.66369e-06, 7.663697e-06, 
    7.663682e-06, 7.663692e-06, 7.663673e-06, 7.663683e-06, 7.663672e-06, 
    7.663675e-06, 7.663672e-06, 7.663669e-06, 7.663665e-06, 7.663659e-06, 
    7.66366e-06, 7.663654e-06, 7.663711e-06, 7.663708e-06, 7.663708e-06, 
    7.663704e-06, 7.663702e-06, 7.663696e-06, 7.663687e-06, 7.663691e-06, 
    7.663684e-06, 7.663682e-06, 7.663692e-06, 7.663686e-06, 7.663705e-06, 
    7.663702e-06, 7.663704e-06, 7.663711e-06, 7.66369e-06, 7.663701e-06, 
    7.663681e-06, 7.663686e-06, 7.663669e-06, 7.663678e-06, 7.663661e-06, 
    7.663653e-06, 7.663647e-06, 7.663639e-06, 7.663706e-06, 7.663708e-06, 
    7.663704e-06, 7.663698e-06, 7.663693e-06, 7.663686e-06, 7.663685e-06, 
    7.663684e-06, 7.663681e-06, 7.663678e-06, 7.663683e-06, 7.663677e-06, 
    7.663702e-06, 7.663689e-06, 7.663709e-06, 7.663702e-06, 7.663699e-06, 
    7.663701e-06, 7.663691e-06, 7.663689e-06, 7.663679e-06, 7.663684e-06, 
    7.663655e-06, 7.663668e-06, 7.663633e-06, 7.663643e-06, 7.663709e-06, 
    7.663706e-06, 7.663695e-06, 7.6637e-06, 7.663685e-06, 7.663682e-06, 
    7.663679e-06, 7.663675e-06, 7.663675e-06, 7.663672e-06, 7.663676e-06, 
    7.663672e-06, 7.663686e-06, 7.66368e-06, 7.663696e-06, 7.663692e-06, 
    7.663694e-06, 7.663696e-06, 7.66369e-06, 7.663683e-06, 7.663683e-06, 
    7.663682e-06, 7.663675e-06, 7.663685e-06, 7.663654e-06, 7.663673e-06, 
    7.663702e-06, 7.663696e-06, 7.663695e-06, 7.663698e-06, 7.663682e-06, 
    7.663688e-06, 7.663672e-06, 7.663677e-06, 7.66367e-06, 7.663673e-06, 
    7.663673e-06, 7.663678e-06, 7.663681e-06, 7.663688e-06, 7.663693e-06, 
    7.663698e-06, 7.663696e-06, 7.663692e-06, 7.663683e-06, 7.663674e-06, 
    7.663676e-06, 7.663671e-06, 7.663686e-06, 7.66368e-06, 7.663682e-06, 
    7.663675e-06, 7.663691e-06, 7.663678e-06, 7.663693e-06, 7.663692e-06, 
    7.663688e-06, 7.66368e-06, 7.663677e-06, 7.663675e-06, 7.663677e-06, 
    7.663682e-06, 7.663683e-06, 7.663688e-06, 7.66369e-06, 7.663692e-06, 
    7.663695e-06, 7.663692e-06, 7.663691e-06, 7.663682e-06, 7.663676e-06, 
    7.663669e-06, 7.663667e-06, 7.663658e-06, 7.663665e-06, 7.663654e-06, 
    7.663663e-06, 7.663647e-06, 7.663677e-06, 7.663664e-06, 7.663688e-06, 
    7.663685e-06, 7.663681e-06, 7.66367e-06, 7.663675e-06, 7.663669e-06, 
    7.663683e-06, 7.663692e-06, 7.663693e-06, 7.663697e-06, 7.663693e-06, 
    7.663693e-06, 7.66369e-06, 7.663692e-06, 7.663682e-06, 7.663687e-06, 
    7.663673e-06, 7.663669e-06, 7.663655e-06, 7.663647e-06, 7.663638e-06, 
    7.663634e-06, 7.663633e-06, 7.663632e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  6.006619e-14, 6.022866e-14, 6.019711e-14, 6.032803e-14, 6.025544e-14, 
    6.034113e-14, 6.009916e-14, 6.023509e-14, 6.014834e-14, 6.008085e-14, 
    6.058172e-14, 6.033387e-14, 6.083893e-14, 6.068116e-14, 6.107725e-14, 
    6.081437e-14, 6.113021e-14, 6.106973e-14, 6.125181e-14, 6.119968e-14, 
    6.143221e-14, 6.127587e-14, 6.155267e-14, 6.139491e-14, 6.141959e-14, 
    6.12707e-14, 6.038383e-14, 6.055087e-14, 6.037392e-14, 6.039775e-14, 
    6.038707e-14, 6.025691e-14, 6.019125e-14, 6.00538e-14, 6.007877e-14, 
    6.017974e-14, 6.040847e-14, 6.03309e-14, 6.052642e-14, 6.052201e-14, 
    6.073934e-14, 6.064139e-14, 6.100625e-14, 6.090265e-14, 6.120185e-14, 
    6.112666e-14, 6.119831e-14, 6.11766e-14, 6.119859e-14, 6.10883e-14, 
    6.113557e-14, 6.103849e-14, 6.065973e-14, 6.077113e-14, 6.043861e-14, 
    6.023823e-14, 6.010512e-14, 6.001055e-14, 6.002393e-14, 6.00494e-14, 
    6.018033e-14, 6.030337e-14, 6.039705e-14, 6.045968e-14, 6.052137e-14, 
    6.070781e-14, 6.08065e-14, 6.102716e-14, 6.098741e-14, 6.105478e-14, 
    6.111918e-14, 6.122717e-14, 6.120941e-14, 6.125695e-14, 6.105303e-14, 
    6.118858e-14, 6.096475e-14, 6.102599e-14, 6.053797e-14, 6.035184e-14, 
    6.027251e-14, 6.020316e-14, 6.00342e-14, 6.015089e-14, 6.01049e-14, 
    6.021434e-14, 6.028381e-14, 6.024946e-14, 6.046139e-14, 6.037903e-14, 
    6.081235e-14, 6.062586e-14, 6.111167e-14, 6.099557e-14, 6.113949e-14, 
    6.106607e-14, 6.119182e-14, 6.107866e-14, 6.127465e-14, 6.131728e-14, 
    6.128815e-14, 6.140007e-14, 6.107238e-14, 6.119829e-14, 6.024849e-14, 
    6.02541e-14, 6.02802e-14, 6.016538e-14, 6.015836e-14, 6.00531e-14, 
    6.014678e-14, 6.018664e-14, 6.028785e-14, 6.034766e-14, 6.040449e-14, 
    6.052939e-14, 6.066872e-14, 6.086338e-14, 6.10031e-14, 6.109668e-14, 
    6.103931e-14, 6.108995e-14, 6.103333e-14, 6.10068e-14, 6.13013e-14, 
    6.113599e-14, 6.138398e-14, 6.137027e-14, 6.125807e-14, 6.137182e-14, 
    6.025803e-14, 6.022578e-14, 6.011373e-14, 6.020143e-14, 6.004164e-14, 
    6.013108e-14, 6.018248e-14, 6.038072e-14, 6.042427e-14, 6.046461e-14, 
    6.054426e-14, 6.064641e-14, 6.082541e-14, 6.098101e-14, 6.112293e-14, 
    6.111254e-14, 6.11162e-14, 6.114786e-14, 6.106939e-14, 6.116075e-14, 
    6.117606e-14, 6.1136e-14, 6.136844e-14, 6.130207e-14, 6.136998e-14, 
    6.132678e-14, 6.023627e-14, 6.029052e-14, 6.026121e-14, 6.031632e-14, 
    6.027748e-14, 6.045006e-14, 6.050177e-14, 6.07435e-14, 6.064439e-14, 
    6.080215e-14, 6.066043e-14, 6.068555e-14, 6.080723e-14, 6.06681e-14, 
    6.09724e-14, 6.07661e-14, 6.11491e-14, 6.094327e-14, 6.116198e-14, 
    6.112232e-14, 6.1188e-14, 6.124678e-14, 6.132073e-14, 6.145701e-14, 
    6.142547e-14, 6.153939e-14, 6.037139e-14, 6.044167e-14, 6.043552e-14, 
    6.050907e-14, 6.056342e-14, 6.068122e-14, 6.086992e-14, 6.079899e-14, 
    6.09292e-14, 6.095532e-14, 6.075751e-14, 6.087896e-14, 6.048872e-14, 
    6.05518e-14, 6.051427e-14, 6.037692e-14, 6.08153e-14, 6.059046e-14, 
    6.10054e-14, 6.088381e-14, 6.123839e-14, 6.106212e-14, 6.140809e-14, 
    6.155565e-14, 6.169451e-14, 6.185644e-14, 6.048005e-14, 6.04323e-14, 
    6.051781e-14, 6.063599e-14, 6.074563e-14, 6.089122e-14, 6.090613e-14, 
    6.093338e-14, 6.100396e-14, 6.106328e-14, 6.094195e-14, 6.107814e-14, 
    6.056637e-14, 6.083481e-14, 6.041422e-14, 6.054095e-14, 6.062903e-14, 
    6.059044e-14, 6.07909e-14, 6.083809e-14, 6.102971e-14, 6.093071e-14, 
    6.151922e-14, 6.125914e-14, 6.197971e-14, 6.177871e-14, 6.041561e-14, 
    6.04799e-14, 6.07034e-14, 6.05971e-14, 6.090095e-14, 6.097563e-14, 
    6.103634e-14, 6.111385e-14, 6.112225e-14, 6.116815e-14, 6.109292e-14, 
    6.11652e-14, 6.089153e-14, 6.101389e-14, 6.06779e-14, 6.075973e-14, 
    6.07221e-14, 6.06808e-14, 6.080825e-14, 6.094386e-14, 6.094681e-14, 
    6.099025e-14, 6.111253e-14, 6.090218e-14, 6.155265e-14, 6.11512e-14, 
    6.054997e-14, 6.06736e-14, 6.069131e-14, 6.064343e-14, 6.096814e-14, 
    6.085056e-14, 6.116704e-14, 6.108159e-14, 6.122159e-14, 6.115203e-14, 
    6.11418e-14, 6.105241e-14, 6.099673e-14, 6.085595e-14, 6.074132e-14, 
    6.065038e-14, 6.067153e-14, 6.077141e-14, 6.095216e-14, 6.112298e-14, 
    6.108558e-14, 6.121095e-14, 6.087894e-14, 6.101823e-14, 6.096439e-14, 
    6.110473e-14, 6.07971e-14, 6.105895e-14, 6.073007e-14, 6.075895e-14, 
    6.084823e-14, 6.102763e-14, 6.106738e-14, 6.11097e-14, 6.108359e-14, 
    6.095675e-14, 6.093599e-14, 6.084608e-14, 6.082121e-14, 6.075267e-14, 
    6.069587e-14, 6.074775e-14, 6.080221e-14, 6.095683e-14, 6.109601e-14, 
    6.12476e-14, 6.12847e-14, 6.146144e-14, 6.131751e-14, 6.155487e-14, 
    6.1353e-14, 6.170232e-14, 6.107419e-14, 6.134715e-14, 6.085231e-14, 
    6.090571e-14, 6.100221e-14, 6.122338e-14, 6.110408e-14, 6.124362e-14, 
    6.093518e-14, 6.077483e-14, 6.073338e-14, 6.06559e-14, 6.073515e-14, 
    6.072871e-14, 6.08045e-14, 6.078015e-14, 6.096196e-14, 6.086433e-14, 
    6.114153e-14, 6.124253e-14, 6.152744e-14, 6.170177e-14, 6.187908e-14, 
    6.195725e-14, 6.198104e-14, 6.199098e-14 ;

 LITTERC =
  5.97623e-05, 5.976215e-05, 5.976218e-05, 5.976206e-05, 5.976213e-05, 
    5.976205e-05, 5.976227e-05, 5.976215e-05, 5.976223e-05, 5.976229e-05, 
    5.976183e-05, 5.976206e-05, 5.97616e-05, 5.976174e-05, 5.976138e-05, 
    5.976162e-05, 5.976133e-05, 5.976139e-05, 5.976122e-05, 5.976127e-05, 
    5.976106e-05, 5.97612e-05, 5.976095e-05, 5.976109e-05, 5.976107e-05, 
    5.97612e-05, 5.976201e-05, 5.976186e-05, 5.976202e-05, 5.9762e-05, 
    5.976201e-05, 5.976213e-05, 5.976219e-05, 5.976231e-05, 5.976229e-05, 
    5.97622e-05, 5.976199e-05, 5.976206e-05, 5.976188e-05, 5.976189e-05, 
    5.976169e-05, 5.976178e-05, 5.976145e-05, 5.976154e-05, 5.976127e-05, 
    5.976134e-05, 5.976127e-05, 5.976129e-05, 5.976127e-05, 5.976137e-05, 
    5.976133e-05, 5.976142e-05, 5.976176e-05, 5.976166e-05, 5.976196e-05, 
    5.976215e-05, 5.976227e-05, 5.976235e-05, 5.976234e-05, 5.976232e-05, 
    5.97622e-05, 5.976209e-05, 5.9762e-05, 5.976194e-05, 5.976189e-05, 
    5.976172e-05, 5.976163e-05, 5.976143e-05, 5.976146e-05, 5.97614e-05, 
    5.976134e-05, 5.976124e-05, 5.976126e-05, 5.976122e-05, 5.97614e-05, 
    5.976128e-05, 5.976148e-05, 5.976143e-05, 5.976187e-05, 5.976204e-05, 
    5.976211e-05, 5.976218e-05, 5.976233e-05, 5.976223e-05, 5.976227e-05, 
    5.976217e-05, 5.97621e-05, 5.976214e-05, 5.976194e-05, 5.976202e-05, 
    5.976162e-05, 5.976179e-05, 5.976135e-05, 5.976145e-05, 5.976132e-05, 
    5.976139e-05, 5.976127e-05, 5.976138e-05, 5.97612e-05, 5.976116e-05, 
    5.976119e-05, 5.976109e-05, 5.976138e-05, 5.976127e-05, 5.976214e-05, 
    5.976213e-05, 5.976211e-05, 5.976221e-05, 5.976222e-05, 5.976231e-05, 
    5.976223e-05, 5.976219e-05, 5.97621e-05, 5.976205e-05, 5.976199e-05, 
    5.976188e-05, 5.976175e-05, 5.976158e-05, 5.976145e-05, 5.976136e-05, 
    5.976141e-05, 5.976137e-05, 5.976142e-05, 5.976145e-05, 5.976118e-05, 
    5.976133e-05, 5.97611e-05, 5.976111e-05, 5.976122e-05, 5.976111e-05, 
    5.976213e-05, 5.976216e-05, 5.976226e-05, 5.976218e-05, 5.976233e-05, 
    5.976225e-05, 5.97622e-05, 5.976202e-05, 5.976198e-05, 5.976194e-05, 
    5.976187e-05, 5.976177e-05, 5.976161e-05, 5.976147e-05, 5.976134e-05, 
    5.976135e-05, 5.976134e-05, 5.976131e-05, 5.976139e-05, 5.97613e-05, 
    5.976129e-05, 5.976133e-05, 5.976111e-05, 5.976117e-05, 5.976111e-05, 
    5.976115e-05, 5.976215e-05, 5.97621e-05, 5.976213e-05, 5.976207e-05, 
    5.976211e-05, 5.976195e-05, 5.97619e-05, 5.976169e-05, 5.976178e-05, 
    5.976163e-05, 5.976176e-05, 5.976174e-05, 5.976163e-05, 5.976175e-05, 
    5.976147e-05, 5.976166e-05, 5.976131e-05, 5.97615e-05, 5.97613e-05, 
    5.976134e-05, 5.976128e-05, 5.976122e-05, 5.976116e-05, 5.976103e-05, 
    5.976106e-05, 5.976096e-05, 5.976202e-05, 5.976196e-05, 5.976197e-05, 
    5.97619e-05, 5.976185e-05, 5.976174e-05, 5.976157e-05, 5.976163e-05, 
    5.976151e-05, 5.976149e-05, 5.976167e-05, 5.976156e-05, 5.976192e-05, 
    5.976186e-05, 5.976189e-05, 5.976202e-05, 5.976162e-05, 5.976182e-05, 
    5.976145e-05, 5.976156e-05, 5.976123e-05, 5.976139e-05, 5.976108e-05, 
    5.976094e-05, 5.976082e-05, 5.976067e-05, 5.976193e-05, 5.976197e-05, 
    5.976189e-05, 5.976178e-05, 5.976168e-05, 5.976155e-05, 5.976154e-05, 
    5.976151e-05, 5.976145e-05, 5.976139e-05, 5.97615e-05, 5.976138e-05, 
    5.976185e-05, 5.97616e-05, 5.976198e-05, 5.976187e-05, 5.976179e-05, 
    5.976182e-05, 5.976164e-05, 5.97616e-05, 5.976142e-05, 5.976151e-05, 
    5.976098e-05, 5.976121e-05, 5.976055e-05, 5.976074e-05, 5.976198e-05, 
    5.976193e-05, 5.976172e-05, 5.976182e-05, 5.976154e-05, 5.976147e-05, 
    5.976142e-05, 5.976135e-05, 5.976134e-05, 5.97613e-05, 5.976137e-05, 
    5.97613e-05, 5.976155e-05, 5.976144e-05, 5.976174e-05, 5.976167e-05, 
    5.97617e-05, 5.976174e-05, 5.976163e-05, 5.97615e-05, 5.97615e-05, 
    5.976146e-05, 5.976135e-05, 5.976154e-05, 5.976095e-05, 5.976131e-05, 
    5.976186e-05, 5.976175e-05, 5.976173e-05, 5.976178e-05, 5.976148e-05, 
    5.976159e-05, 5.97613e-05, 5.976138e-05, 5.976125e-05, 5.976131e-05, 
    5.976132e-05, 5.97614e-05, 5.976145e-05, 5.976158e-05, 5.976169e-05, 
    5.976177e-05, 5.976175e-05, 5.976166e-05, 5.976149e-05, 5.976134e-05, 
    5.976137e-05, 5.976126e-05, 5.976156e-05, 5.976143e-05, 5.976148e-05, 
    5.976135e-05, 5.976163e-05, 5.97614e-05, 5.97617e-05, 5.976167e-05, 
    5.976159e-05, 5.976142e-05, 5.976139e-05, 5.976135e-05, 5.976137e-05, 
    5.976149e-05, 5.976151e-05, 5.976159e-05, 5.976161e-05, 5.976167e-05, 
    5.976173e-05, 5.976168e-05, 5.976163e-05, 5.976149e-05, 5.976136e-05, 
    5.976122e-05, 5.976119e-05, 5.976103e-05, 5.976116e-05, 5.976094e-05, 
    5.976113e-05, 5.976081e-05, 5.976138e-05, 5.976113e-05, 5.976158e-05, 
    5.976154e-05, 5.976145e-05, 5.976125e-05, 5.976135e-05, 5.976123e-05, 
    5.976151e-05, 5.976166e-05, 5.976169e-05, 5.976177e-05, 5.976169e-05, 
    5.97617e-05, 5.976163e-05, 5.976165e-05, 5.976149e-05, 5.976157e-05, 
    5.976132e-05, 5.976123e-05, 5.976097e-05, 5.976081e-05, 5.976065e-05, 
    5.976058e-05, 5.976055e-05, 5.976054e-05 ;

 LITTERC_HR =
  9.690869e-13, 9.717061e-13, 9.711974e-13, 9.733079e-13, 9.721376e-13, 
    9.735191e-13, 9.696185e-13, 9.718098e-13, 9.704114e-13, 9.693234e-13, 
    9.773974e-13, 9.734021e-13, 9.815437e-13, 9.790004e-13, 9.853853e-13, 
    9.811477e-13, 9.86239e-13, 9.852641e-13, 9.881991e-13, 9.873587e-13, 
    9.911072e-13, 9.885869e-13, 9.93049e-13, 9.90506e-13, 9.909036e-13, 
    9.885037e-13, 9.742074e-13, 9.769001e-13, 9.740476e-13, 9.744318e-13, 
    9.742596e-13, 9.721616e-13, 9.711031e-13, 9.688872e-13, 9.692898e-13, 
    9.709175e-13, 9.746046e-13, 9.733541e-13, 9.765059e-13, 9.764349e-13, 
    9.799384e-13, 9.783593e-13, 9.842408e-13, 9.825708e-13, 9.873939e-13, 
    9.861817e-13, 9.873367e-13, 9.869868e-13, 9.873413e-13, 9.855635e-13, 
    9.863253e-13, 9.847605e-13, 9.78655e-13, 9.804507e-13, 9.750905e-13, 
    9.718604e-13, 9.697145e-13, 9.6819e-13, 9.684057e-13, 9.688164e-13, 
    9.70927e-13, 9.729104e-13, 9.744206e-13, 9.754301e-13, 9.764246e-13, 
    9.7943e-13, 9.810209e-13, 9.845779e-13, 9.83937e-13, 9.85023e-13, 
    9.860612e-13, 9.87802e-13, 9.875156e-13, 9.88282e-13, 9.84995e-13, 
    9.871798e-13, 9.835717e-13, 9.845591e-13, 9.766921e-13, 9.736917e-13, 
    9.724129e-13, 9.712951e-13, 9.685714e-13, 9.704525e-13, 9.69711e-13, 
    9.714752e-13, 9.725951e-13, 9.720413e-13, 9.754578e-13, 9.741301e-13, 
    9.811151e-13, 9.78109e-13, 9.859402e-13, 9.840686e-13, 9.863886e-13, 
    9.852052e-13, 9.872322e-13, 9.85408e-13, 9.885674e-13, 9.892546e-13, 
    9.887849e-13, 9.90589e-13, 9.853068e-13, 9.873365e-13, 9.720257e-13, 
    9.721161e-13, 9.725369e-13, 9.70686e-13, 9.705728e-13, 9.68876e-13, 
    9.703861e-13, 9.710287e-13, 9.726602e-13, 9.736242e-13, 9.745404e-13, 
    9.765538e-13, 9.787998e-13, 9.819377e-13, 9.841899e-13, 9.856984e-13, 
    9.847737e-13, 9.855901e-13, 9.846774e-13, 9.842496e-13, 9.88997e-13, 
    9.863322e-13, 9.903297e-13, 9.901088e-13, 9.883002e-13, 9.901336e-13, 
    9.721795e-13, 9.716597e-13, 9.698534e-13, 9.712671e-13, 9.686912e-13, 
    9.70133e-13, 9.709616e-13, 9.741572e-13, 9.748594e-13, 9.755095e-13, 
    9.767935e-13, 9.784401e-13, 9.813257e-13, 9.838339e-13, 9.861217e-13, 
    9.859542e-13, 9.860131e-13, 9.865236e-13, 9.852585e-13, 9.867312e-13, 
    9.869781e-13, 9.863323e-13, 9.900791e-13, 9.890094e-13, 9.90104e-13, 
    9.894077e-13, 9.718287e-13, 9.727034e-13, 9.722308e-13, 9.731192e-13, 
    9.72493e-13, 9.752751e-13, 9.761085e-13, 9.800055e-13, 9.784076e-13, 
    9.809508e-13, 9.786663e-13, 9.790711e-13, 9.810325e-13, 9.7879e-13, 
    9.836951e-13, 9.803696e-13, 9.865434e-13, 9.832255e-13, 9.867512e-13, 
    9.861118e-13, 9.871705e-13, 9.88118e-13, 9.893101e-13, 9.915069e-13, 
    9.909985e-13, 9.928348e-13, 9.740068e-13, 9.751398e-13, 9.750406e-13, 
    9.762262e-13, 9.771025e-13, 9.790014e-13, 9.820431e-13, 9.808999e-13, 
    9.829987e-13, 9.834197e-13, 9.802312e-13, 9.821889e-13, 9.758982e-13, 
    9.769152e-13, 9.763101e-13, 9.740959e-13, 9.811626e-13, 9.775383e-13, 
    9.842271e-13, 9.82267e-13, 9.879829e-13, 9.851415e-13, 9.907185e-13, 
    9.930969e-13, 9.953354e-13, 9.979456e-13, 9.757585e-13, 9.749889e-13, 
    9.763673e-13, 9.782722e-13, 9.800396e-13, 9.823865e-13, 9.826268e-13, 
    9.830661e-13, 9.842039e-13, 9.8516e-13, 9.832044e-13, 9.853997e-13, 
    9.771499e-13, 9.814773e-13, 9.746973e-13, 9.767403e-13, 9.781602e-13, 
    9.775379e-13, 9.807693e-13, 9.815302e-13, 9.84619e-13, 9.83023e-13, 
    9.925097e-13, 9.883174e-13, 9.999327e-13, 9.966926e-13, 9.747198e-13, 
    9.757562e-13, 9.793588e-13, 9.776454e-13, 9.825434e-13, 9.837473e-13, 
    9.847259e-13, 9.859754e-13, 9.861106e-13, 9.868507e-13, 9.856378e-13, 
    9.86803e-13, 9.823915e-13, 9.84364e-13, 9.789479e-13, 9.80267e-13, 
    9.796605e-13, 9.789946e-13, 9.81049e-13, 9.832351e-13, 9.832826e-13, 
    9.839829e-13, 9.859539e-13, 9.825632e-13, 9.930485e-13, 9.865775e-13, 
    9.768857e-13, 9.788785e-13, 9.79164e-13, 9.783922e-13, 9.836265e-13, 
    9.817312e-13, 9.868328e-13, 9.854553e-13, 9.87712e-13, 9.865908e-13, 
    9.864258e-13, 9.84985e-13, 9.840873e-13, 9.818179e-13, 9.799701e-13, 
    9.785043e-13, 9.788453e-13, 9.804552e-13, 9.833689e-13, 9.861225e-13, 
    9.855195e-13, 9.875406e-13, 9.821886e-13, 9.844338e-13, 9.83566e-13, 
    9.858284e-13, 9.808694e-13, 9.850903e-13, 9.797888e-13, 9.802544e-13, 
    9.816936e-13, 9.845855e-13, 9.852261e-13, 9.859084e-13, 9.854876e-13, 
    9.834429e-13, 9.831082e-13, 9.816588e-13, 9.81258e-13, 9.801531e-13, 
    9.792375e-13, 9.800739e-13, 9.809516e-13, 9.834441e-13, 9.856877e-13, 
    9.881313e-13, 9.887294e-13, 9.915783e-13, 9.892584e-13, 9.930844e-13, 
    9.898302e-13, 9.954612e-13, 9.853359e-13, 9.897361e-13, 9.817593e-13, 
    9.826202e-13, 9.841756e-13, 9.877409e-13, 9.858178e-13, 9.880671e-13, 
    9.830951e-13, 9.805104e-13, 9.798422e-13, 9.785933e-13, 9.798707e-13, 
    9.797668e-13, 9.809886e-13, 9.805961e-13, 9.835268e-13, 9.819531e-13, 
    9.864214e-13, 9.880496e-13, 9.926422e-13, 9.954523e-13, 9.983104e-13, 
    9.995705e-13, 9.99954e-13, 1.000114e-12 ;

 LITTERC_LOSS =
  1.79474e-12, 1.79959e-12, 1.798648e-12, 1.802557e-12, 1.80039e-12, 
    1.802948e-12, 1.795724e-12, 1.799782e-12, 1.797192e-12, 1.795177e-12, 
    1.810131e-12, 1.802731e-12, 1.81781e-12, 1.813099e-12, 1.824925e-12, 
    1.817076e-12, 1.826506e-12, 1.8247e-12, 1.830136e-12, 1.828579e-12, 
    1.835521e-12, 1.830854e-12, 1.839118e-12, 1.834408e-12, 1.835145e-12, 
    1.8307e-12, 1.804223e-12, 1.80921e-12, 1.803927e-12, 1.804638e-12, 
    1.804319e-12, 1.800434e-12, 1.798473e-12, 1.79437e-12, 1.795115e-12, 
    1.79813e-12, 1.804958e-12, 1.802643e-12, 1.80848e-12, 1.808348e-12, 
    1.814837e-12, 1.811912e-12, 1.822805e-12, 1.819712e-12, 1.828644e-12, 
    1.826399e-12, 1.828539e-12, 1.82789e-12, 1.828547e-12, 1.825255e-12, 
    1.826666e-12, 1.823767e-12, 1.81246e-12, 1.815786e-12, 1.805858e-12, 
    1.799876e-12, 1.795902e-12, 1.793079e-12, 1.793478e-12, 1.794239e-12, 
    1.798147e-12, 1.801821e-12, 1.804618e-12, 1.806487e-12, 1.808329e-12, 
    1.813895e-12, 1.816842e-12, 1.823429e-12, 1.822242e-12, 1.824254e-12, 
    1.826176e-12, 1.8294e-12, 1.82887e-12, 1.830289e-12, 1.824202e-12, 
    1.828248e-12, 1.821566e-12, 1.823394e-12, 1.808825e-12, 1.803268e-12, 
    1.800899e-12, 1.798829e-12, 1.793785e-12, 1.797269e-12, 1.795895e-12, 
    1.799163e-12, 1.801237e-12, 1.800211e-12, 1.806539e-12, 1.80408e-12, 
    1.817016e-12, 1.811449e-12, 1.825952e-12, 1.822486e-12, 1.826783e-12, 
    1.824591e-12, 1.828345e-12, 1.824967e-12, 1.830818e-12, 1.83209e-12, 
    1.831221e-12, 1.834562e-12, 1.824779e-12, 1.828538e-12, 1.800182e-12, 
    1.80035e-12, 1.801129e-12, 1.797701e-12, 1.797492e-12, 1.794349e-12, 
    1.797146e-12, 1.798336e-12, 1.801357e-12, 1.803143e-12, 1.80484e-12, 
    1.808568e-12, 1.812728e-12, 1.81854e-12, 1.822711e-12, 1.825504e-12, 
    1.823792e-12, 1.825304e-12, 1.823613e-12, 1.822821e-12, 1.831613e-12, 
    1.826678e-12, 1.834081e-12, 1.833673e-12, 1.830323e-12, 1.833719e-12, 
    1.800467e-12, 1.799504e-12, 1.796159e-12, 1.798777e-12, 1.794007e-12, 
    1.796677e-12, 1.798211e-12, 1.80413e-12, 1.80543e-12, 1.806634e-12, 
    1.809012e-12, 1.812062e-12, 1.817406e-12, 1.822051e-12, 1.826288e-12, 
    1.825978e-12, 1.826087e-12, 1.827033e-12, 1.82469e-12, 1.827417e-12, 
    1.827874e-12, 1.826678e-12, 1.833618e-12, 1.831636e-12, 1.833664e-12, 
    1.832374e-12, 1.799818e-12, 1.801437e-12, 1.800562e-12, 1.802207e-12, 
    1.801048e-12, 1.8062e-12, 1.807744e-12, 1.814961e-12, 1.812002e-12, 
    1.816712e-12, 1.812481e-12, 1.81323e-12, 1.816863e-12, 1.81271e-12, 
    1.821794e-12, 1.815635e-12, 1.827069e-12, 1.820925e-12, 1.827454e-12, 
    1.82627e-12, 1.828231e-12, 1.829986e-12, 1.832193e-12, 1.836262e-12, 
    1.83532e-12, 1.838721e-12, 1.803851e-12, 1.80595e-12, 1.805766e-12, 
    1.807962e-12, 1.809585e-12, 1.813101e-12, 1.818735e-12, 1.816617e-12, 
    1.820505e-12, 1.821284e-12, 1.815379e-12, 1.819005e-12, 1.807354e-12, 
    1.809238e-12, 1.808117e-12, 1.804016e-12, 1.817104e-12, 1.810392e-12, 
    1.82278e-12, 1.819149e-12, 1.829735e-12, 1.824473e-12, 1.834802e-12, 
    1.839207e-12, 1.843352e-12, 1.848187e-12, 1.807095e-12, 1.80567e-12, 
    1.808223e-12, 1.811751e-12, 1.815024e-12, 1.819371e-12, 1.819816e-12, 
    1.820629e-12, 1.822737e-12, 1.824507e-12, 1.820885e-12, 1.824951e-12, 
    1.809672e-12, 1.817687e-12, 1.80513e-12, 1.808914e-12, 1.811543e-12, 
    1.810391e-12, 1.816376e-12, 1.817785e-12, 1.823505e-12, 1.82055e-12, 
    1.838119e-12, 1.830355e-12, 1.851867e-12, 1.845866e-12, 1.805172e-12, 
    1.807091e-12, 1.813763e-12, 1.81059e-12, 1.819661e-12, 1.821891e-12, 
    1.823703e-12, 1.826017e-12, 1.826268e-12, 1.827638e-12, 1.825392e-12, 
    1.82755e-12, 1.81938e-12, 1.823033e-12, 1.813002e-12, 1.815445e-12, 
    1.814322e-12, 1.813089e-12, 1.816894e-12, 1.820942e-12, 1.82103e-12, 
    1.822327e-12, 1.825978e-12, 1.819698e-12, 1.839117e-12, 1.827132e-12, 
    1.809183e-12, 1.812874e-12, 1.813403e-12, 1.811973e-12, 1.821667e-12, 
    1.818157e-12, 1.827605e-12, 1.825054e-12, 1.829234e-12, 1.827157e-12, 
    1.826851e-12, 1.824183e-12, 1.822521e-12, 1.818318e-12, 1.814896e-12, 
    1.812181e-12, 1.812812e-12, 1.815794e-12, 1.82119e-12, 1.82629e-12, 
    1.825173e-12, 1.828916e-12, 1.819004e-12, 1.823162e-12, 1.821555e-12, 
    1.825745e-12, 1.816561e-12, 1.824378e-12, 1.81456e-12, 1.815422e-12, 
    1.818087e-12, 1.823443e-12, 1.82463e-12, 1.825893e-12, 1.825114e-12, 
    1.821327e-12, 1.820707e-12, 1.818023e-12, 1.817281e-12, 1.815234e-12, 
    1.813539e-12, 1.815088e-12, 1.816713e-12, 1.82133e-12, 1.825484e-12, 
    1.83001e-12, 1.831118e-12, 1.836394e-12, 1.832097e-12, 1.839183e-12, 
    1.833157e-12, 1.843585e-12, 1.824833e-12, 1.832982e-12, 1.818209e-12, 
    1.819803e-12, 1.822684e-12, 1.829287e-12, 1.825725e-12, 1.829891e-12, 
    1.820683e-12, 1.815896e-12, 1.814658e-12, 1.812346e-12, 1.814711e-12, 
    1.814519e-12, 1.816782e-12, 1.816055e-12, 1.821483e-12, 1.818568e-12, 
    1.826843e-12, 1.829859e-12, 1.838364e-12, 1.843569e-12, 1.848862e-12, 
    1.851196e-12, 1.851906e-12, 1.852203e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  1.701311e-18, 1.701567e-18, 1.701518e-18, 1.701722e-18, 1.701611e-18, 
    1.701743e-18, 1.701365e-18, 1.701575e-18, 1.701442e-18, 1.701337e-18, 
    1.702113e-18, 1.701732e-18, 1.702531e-18, 1.702283e-18, 1.702912e-18, 
    1.702489e-18, 1.702998e-18, 1.702905e-18, 1.703199e-18, 1.703115e-18, 
    1.70348e-18, 1.703238e-18, 1.703679e-18, 1.703425e-18, 1.703463e-18, 
    1.703229e-18, 1.701813e-18, 1.702064e-18, 1.701797e-18, 1.701833e-18, 
    1.701818e-18, 1.701612e-18, 1.701504e-18, 1.701295e-18, 1.701334e-18, 
    1.701489e-18, 1.70185e-18, 1.701731e-18, 1.702041e-18, 1.702034e-18, 
    1.702377e-18, 1.702222e-18, 1.702803e-18, 1.702639e-18, 1.703119e-18, 
    1.702997e-18, 1.703112e-18, 1.703078e-18, 1.703112e-18, 1.702934e-18, 
    1.70301e-18, 1.702855e-18, 1.70225e-18, 1.702426e-18, 1.701899e-18, 
    1.701575e-18, 1.701373e-18, 1.701226e-18, 1.701247e-18, 1.701286e-18, 
    1.70149e-18, 1.701687e-18, 1.701836e-18, 1.701935e-18, 1.702033e-18, 
    1.702317e-18, 1.702479e-18, 1.702834e-18, 1.702774e-18, 1.702879e-18, 
    1.702985e-18, 1.703158e-18, 1.70313e-18, 1.703205e-18, 1.702879e-18, 
    1.703094e-18, 1.702739e-18, 1.702835e-18, 1.702042e-18, 1.701764e-18, 
    1.70163e-18, 1.701527e-18, 1.701263e-18, 1.701444e-18, 1.701372e-18, 
    1.701547e-18, 1.701656e-18, 1.701603e-18, 1.701937e-18, 1.701807e-18, 
    1.702488e-18, 1.702194e-18, 1.702973e-18, 1.702787e-18, 1.703018e-18, 
    1.702901e-18, 1.7031e-18, 1.702921e-18, 1.703235e-18, 1.7033e-18, 
    1.703255e-18, 1.703437e-18, 1.70291e-18, 1.70311e-18, 1.701601e-18, 
    1.701609e-18, 1.701651e-18, 1.701467e-18, 1.701456e-18, 1.701293e-18, 
    1.70144e-18, 1.701501e-18, 1.701664e-18, 1.701757e-18, 1.701846e-18, 
    1.702044e-18, 1.702262e-18, 1.702572e-18, 1.702798e-18, 1.70295e-18, 
    1.702858e-18, 1.702939e-18, 1.702848e-18, 1.702806e-18, 1.703274e-18, 
    1.70301e-18, 1.70341e-18, 1.703389e-18, 1.703206e-18, 1.703391e-18, 
    1.701615e-18, 1.701566e-18, 1.701387e-18, 1.701527e-18, 1.701275e-18, 
    1.701414e-18, 1.701493e-18, 1.701806e-18, 1.701879e-18, 1.701941e-18, 
    1.702068e-18, 1.70223e-18, 1.702512e-18, 1.702761e-18, 1.702992e-18, 
    1.702975e-18, 1.702981e-18, 1.703031e-18, 1.702905e-18, 1.703052e-18, 
    1.703075e-18, 1.703012e-18, 1.703386e-18, 1.703279e-18, 1.703388e-18, 
    1.703319e-18, 1.701582e-18, 1.701667e-18, 1.701621e-18, 1.701706e-18, 
    1.701645e-18, 1.701914e-18, 1.701995e-18, 1.702379e-18, 1.702226e-18, 
    1.702474e-18, 1.702252e-18, 1.70229e-18, 1.702475e-18, 1.702265e-18, 
    1.702744e-18, 1.702413e-18, 1.703033e-18, 1.702694e-18, 1.703054e-18, 
    1.702991e-18, 1.703097e-18, 1.703189e-18, 1.703309e-18, 1.703525e-18, 
    1.703476e-18, 1.70366e-18, 1.701795e-18, 1.701903e-18, 1.701897e-18, 
    1.702012e-18, 1.702097e-18, 1.702286e-18, 1.702585e-18, 1.702473e-18, 
    1.702681e-18, 1.702722e-18, 1.702408e-18, 1.702598e-18, 1.701978e-18, 
    1.702075e-18, 1.702019e-18, 1.701801e-18, 1.702494e-18, 1.702136e-18, 
    1.702802e-18, 1.702608e-18, 1.703176e-18, 1.702889e-18, 1.703448e-18, 
    1.703679e-18, 1.703913e-18, 1.704169e-18, 1.701966e-18, 1.701892e-18, 
    1.702027e-18, 1.702209e-18, 1.702387e-18, 1.702619e-18, 1.702644e-18, 
    1.702687e-18, 1.702801e-18, 1.702896e-18, 1.702697e-18, 1.70292e-18, 
    1.70209e-18, 1.702527e-18, 1.701861e-18, 1.702057e-18, 1.7022e-18, 
    1.70214e-18, 1.702461e-18, 1.702536e-18, 1.702839e-18, 1.702684e-18, 
    1.703619e-18, 1.703204e-18, 1.704375e-18, 1.704044e-18, 1.701865e-18, 
    1.701967e-18, 1.702318e-18, 1.702151e-18, 1.702636e-18, 1.702754e-18, 
    1.702853e-18, 1.702975e-18, 1.70299e-18, 1.703063e-18, 1.702944e-18, 
    1.703059e-18, 1.702619e-18, 1.702816e-18, 1.702281e-18, 1.702409e-18, 
    1.702352e-18, 1.702286e-18, 1.702489e-18, 1.702699e-18, 1.702709e-18, 
    1.702776e-18, 1.702956e-18, 1.702638e-18, 1.703663e-18, 1.70302e-18, 
    1.702078e-18, 1.702267e-18, 1.702301e-18, 1.702226e-18, 1.702742e-18, 
    1.702554e-18, 1.703062e-18, 1.702926e-18, 1.70315e-18, 1.703038e-18, 
    1.703021e-18, 1.702878e-18, 1.702788e-18, 1.702562e-18, 1.70238e-18, 
    1.702238e-18, 1.702271e-18, 1.702427e-18, 1.702714e-18, 1.702989e-18, 
    1.702928e-18, 1.703133e-18, 1.702601e-18, 1.702821e-18, 1.702734e-18, 
    1.702962e-18, 1.702469e-18, 1.702872e-18, 1.702364e-18, 1.70241e-18, 
    1.702551e-18, 1.702832e-18, 1.702903e-18, 1.702968e-18, 1.702929e-18, 
    1.702722e-18, 1.70269e-18, 1.702549e-18, 1.702507e-18, 1.7024e-18, 
    1.70231e-18, 1.702391e-18, 1.702476e-18, 1.702724e-18, 1.702946e-18, 
    1.70319e-18, 1.703252e-18, 1.703524e-18, 1.703294e-18, 1.703666e-18, 
    1.703339e-18, 1.703911e-18, 1.702904e-18, 1.70334e-18, 1.702559e-18, 
    1.702644e-18, 1.702793e-18, 1.703146e-18, 1.702961e-18, 1.70318e-18, 
    1.70269e-18, 1.70243e-18, 1.702369e-18, 1.702245e-18, 1.702372e-18, 
    1.702362e-18, 1.702483e-18, 1.702444e-18, 1.702733e-18, 1.702578e-18, 
    1.703019e-18, 1.70318e-18, 1.703639e-18, 1.703919e-18, 1.704213e-18, 
    1.70434e-18, 1.704379e-18, 1.704395e-18 ;

 MEG_acetic_acid =
  2.551966e-19, 2.55235e-19, 2.552277e-19, 2.552583e-19, 2.552416e-19, 
    2.552615e-19, 2.552048e-19, 2.552363e-19, 2.552163e-19, 2.552005e-19, 
    2.553169e-19, 2.552598e-19, 2.553796e-19, 2.553425e-19, 2.554368e-19, 
    2.553734e-19, 2.554498e-19, 2.554357e-19, 2.554798e-19, 2.554672e-19, 
    2.555221e-19, 2.554857e-19, 2.555519e-19, 2.555137e-19, 2.555194e-19, 
    2.554843e-19, 2.55272e-19, 2.553095e-19, 2.552696e-19, 2.55275e-19, 
    2.552727e-19, 2.552417e-19, 2.552256e-19, 2.551942e-19, 2.552001e-19, 
    2.552234e-19, 2.552774e-19, 2.552596e-19, 2.553061e-19, 2.553051e-19, 
    2.553565e-19, 2.553333e-19, 2.554204e-19, 2.553958e-19, 2.554678e-19, 
    2.554495e-19, 2.554668e-19, 2.554617e-19, 2.554668e-19, 2.554401e-19, 
    2.554515e-19, 2.554283e-19, 2.553375e-19, 2.553639e-19, 2.552848e-19, 
    2.552363e-19, 2.55206e-19, 2.55184e-19, 2.551871e-19, 2.551929e-19, 
    2.552235e-19, 2.55253e-19, 2.552754e-19, 2.552902e-19, 2.553049e-19, 
    2.553476e-19, 2.553718e-19, 2.55425e-19, 2.554161e-19, 2.554318e-19, 
    2.554477e-19, 2.554737e-19, 2.554695e-19, 2.554808e-19, 2.554318e-19, 
    2.554641e-19, 2.554108e-19, 2.554253e-19, 2.553063e-19, 2.552645e-19, 
    2.552445e-19, 2.552291e-19, 2.551894e-19, 2.552167e-19, 2.552058e-19, 
    2.552321e-19, 2.552484e-19, 2.552404e-19, 2.552906e-19, 2.55271e-19, 
    2.553733e-19, 2.553292e-19, 2.554459e-19, 2.55418e-19, 2.554527e-19, 
    2.554351e-19, 2.55465e-19, 2.554381e-19, 2.554852e-19, 2.55495e-19, 
    2.554883e-19, 2.555155e-19, 2.554366e-19, 2.554665e-19, 2.552401e-19, 
    2.552414e-19, 2.552476e-19, 2.5522e-19, 2.552185e-19, 2.551939e-19, 
    2.55216e-19, 2.552252e-19, 2.552496e-19, 2.552635e-19, 2.552769e-19, 
    2.553066e-19, 2.553393e-19, 2.553858e-19, 2.554198e-19, 2.554424e-19, 
    2.554287e-19, 2.554408e-19, 2.554272e-19, 2.554209e-19, 2.554911e-19, 
    2.554515e-19, 2.555115e-19, 2.555083e-19, 2.554809e-19, 2.555087e-19, 
    2.552423e-19, 2.552348e-19, 2.552081e-19, 2.55229e-19, 2.551913e-19, 
    2.552121e-19, 2.552239e-19, 2.552708e-19, 2.552818e-19, 2.552911e-19, 
    2.553102e-19, 2.553344e-19, 2.553768e-19, 2.554142e-19, 2.554488e-19, 
    2.554463e-19, 2.554472e-19, 2.554546e-19, 2.554358e-19, 2.554577e-19, 
    2.554612e-19, 2.554518e-19, 2.555078e-19, 2.554918e-19, 2.555082e-19, 
    2.554978e-19, 2.552373e-19, 2.5525e-19, 2.552431e-19, 2.55256e-19, 
    2.552467e-19, 2.552871e-19, 2.552992e-19, 2.553568e-19, 2.553338e-19, 
    2.553712e-19, 2.553378e-19, 2.553436e-19, 2.553713e-19, 2.553398e-19, 
    2.554116e-19, 2.553619e-19, 2.554549e-19, 2.554041e-19, 2.55458e-19, 
    2.554487e-19, 2.554645e-19, 2.554784e-19, 2.554963e-19, 2.555288e-19, 
    2.555214e-19, 2.55549e-19, 2.552692e-19, 2.552854e-19, 2.552845e-19, 
    2.553019e-19, 2.553146e-19, 2.553428e-19, 2.553877e-19, 2.55371e-19, 
    2.554022e-19, 2.554083e-19, 2.553611e-19, 2.553896e-19, 2.552967e-19, 
    2.553112e-19, 2.553029e-19, 2.552702e-19, 2.553742e-19, 2.553204e-19, 
    2.554202e-19, 2.553911e-19, 2.554763e-19, 2.554334e-19, 2.555172e-19, 
    2.555519e-19, 2.555869e-19, 2.556253e-19, 2.552948e-19, 2.552838e-19, 
    2.553041e-19, 2.553313e-19, 2.55358e-19, 2.553928e-19, 2.553966e-19, 
    2.55403e-19, 2.554202e-19, 2.554344e-19, 2.554046e-19, 2.55438e-19, 
    2.553136e-19, 2.55379e-19, 2.552791e-19, 2.553085e-19, 2.553299e-19, 
    2.55321e-19, 2.553692e-19, 2.553804e-19, 2.554258e-19, 2.554026e-19, 
    2.555429e-19, 2.554806e-19, 2.556562e-19, 2.556066e-19, 2.552798e-19, 
    2.55295e-19, 2.553476e-19, 2.553227e-19, 2.553954e-19, 2.554131e-19, 
    2.55428e-19, 2.554462e-19, 2.554485e-19, 2.554594e-19, 2.554415e-19, 
    2.554589e-19, 2.553929e-19, 2.554224e-19, 2.553422e-19, 2.553614e-19, 
    2.553527e-19, 2.553429e-19, 2.553733e-19, 2.554049e-19, 2.554064e-19, 
    2.554164e-19, 2.554433e-19, 2.553957e-19, 2.555495e-19, 2.55453e-19, 
    2.553117e-19, 2.553401e-19, 2.553451e-19, 2.553339e-19, 2.554113e-19, 
    2.553831e-19, 2.554592e-19, 2.554388e-19, 2.554725e-19, 2.554557e-19, 
    2.554532e-19, 2.554318e-19, 2.554183e-19, 2.553843e-19, 2.553569e-19, 
    2.553357e-19, 2.553407e-19, 2.55364e-19, 2.55407e-19, 2.554484e-19, 
    2.554392e-19, 2.5547e-19, 2.553901e-19, 2.554231e-19, 2.554101e-19, 
    2.554443e-19, 2.553704e-19, 2.554309e-19, 2.553546e-19, 2.553615e-19, 
    2.553826e-19, 2.554248e-19, 2.554354e-19, 2.554452e-19, 2.554393e-19, 
    2.554083e-19, 2.554036e-19, 2.553823e-19, 2.55376e-19, 2.5536e-19, 
    2.553465e-19, 2.553587e-19, 2.553713e-19, 2.554086e-19, 2.554419e-19, 
    2.554785e-19, 2.554877e-19, 2.555286e-19, 2.554941e-19, 2.555499e-19, 
    2.555008e-19, 2.555866e-19, 2.554355e-19, 2.55501e-19, 2.553838e-19, 
    2.553966e-19, 2.554189e-19, 2.554719e-19, 2.554441e-19, 2.55477e-19, 
    2.554034e-19, 2.553645e-19, 2.553554e-19, 2.553368e-19, 2.553558e-19, 
    2.553543e-19, 2.553724e-19, 2.553666e-19, 2.554099e-19, 2.553867e-19, 
    2.554529e-19, 2.554769e-19, 2.555458e-19, 2.555878e-19, 2.556319e-19, 
    2.55651e-19, 2.556569e-19, 2.556593e-19 ;

 MEG_acetone =
  8.512738e-17, 8.513581e-17, 8.513421e-17, 8.514093e-17, 8.513726e-17, 
    8.514161e-17, 8.512916e-17, 8.513608e-17, 8.513171e-17, 8.512824e-17, 
    8.515378e-17, 8.514124e-17, 8.516754e-17, 8.51594e-17, 8.518011e-17, 
    8.516618e-17, 8.518295e-17, 8.517988e-17, 8.518956e-17, 8.518679e-17, 
    8.519884e-17, 8.519084e-17, 8.520539e-17, 8.519702e-17, 8.519826e-17, 
    8.519055e-17, 8.514392e-17, 8.515216e-17, 8.51434e-17, 8.514458e-17, 
    8.514409e-17, 8.513728e-17, 8.513374e-17, 8.512685e-17, 8.512813e-17, 
    8.513326e-17, 8.514512e-17, 8.51412e-17, 8.515141e-17, 8.515118e-17, 
    8.516247e-17, 8.515737e-17, 8.517651e-17, 8.51711e-17, 8.518691e-17, 
    8.518291e-17, 8.518669e-17, 8.518557e-17, 8.518671e-17, 8.518085e-17, 
    8.518335e-17, 8.517824e-17, 8.51583e-17, 8.516409e-17, 8.514674e-17, 
    8.513608e-17, 8.512944e-17, 8.51246e-17, 8.512528e-17, 8.512655e-17, 
    8.513328e-17, 8.513977e-17, 8.514467e-17, 8.514791e-17, 8.515115e-17, 
    8.516051e-17, 8.516584e-17, 8.517753e-17, 8.517556e-17, 8.517901e-17, 
    8.518252e-17, 8.518821e-17, 8.518729e-17, 8.518977e-17, 8.517902e-17, 
    8.518611e-17, 8.51744e-17, 8.517758e-17, 8.515145e-17, 8.514228e-17, 
    8.51379e-17, 8.513449e-17, 8.51258e-17, 8.513177e-17, 8.51294e-17, 
    8.513516e-17, 8.513874e-17, 8.5137e-17, 8.514801e-17, 8.51437e-17, 
    8.516616e-17, 8.515647e-17, 8.518211e-17, 8.517598e-17, 8.51836e-17, 
    8.517973e-17, 8.518631e-17, 8.51804e-17, 8.519074e-17, 8.519291e-17, 
    8.519142e-17, 8.519739e-17, 8.518006e-17, 8.518664e-17, 8.513692e-17, 
    8.51372e-17, 8.513858e-17, 8.513251e-17, 8.513217e-17, 8.512679e-17, 
    8.513163e-17, 8.513365e-17, 8.513899e-17, 8.514206e-17, 8.514501e-17, 
    8.515151e-17, 8.515869e-17, 8.516891e-17, 8.517637e-17, 8.518135e-17, 
    8.517833e-17, 8.518099e-17, 8.5178e-17, 8.517661e-17, 8.519205e-17, 
    8.518334e-17, 8.519653e-17, 8.519582e-17, 8.51898e-17, 8.51959e-17, 
    8.513741e-17, 8.513577e-17, 8.51299e-17, 8.513449e-17, 8.512621e-17, 
    8.513078e-17, 8.513336e-17, 8.514367e-17, 8.514607e-17, 8.514813e-17, 
    8.515231e-17, 8.515763e-17, 8.516694e-17, 8.517515e-17, 8.518274e-17, 
    8.51822e-17, 8.518238e-17, 8.518403e-17, 8.517989e-17, 8.518471e-17, 
    8.518546e-17, 8.51834e-17, 8.519572e-17, 8.51922e-17, 8.51958e-17, 
    8.519352e-17, 8.513631e-17, 8.51391e-17, 8.513758e-17, 8.51404e-17, 
    8.513837e-17, 8.514724e-17, 8.51499e-17, 8.516255e-17, 8.51575e-17, 
    8.516569e-17, 8.515837e-17, 8.515963e-17, 8.516572e-17, 8.515881e-17, 
    8.517458e-17, 8.516366e-17, 8.518409e-17, 8.517292e-17, 8.518477e-17, 
    8.518271e-17, 8.518619e-17, 8.518924e-17, 8.519318e-17, 8.520032e-17, 
    8.519869e-17, 8.520476e-17, 8.514331e-17, 8.514688e-17, 8.514666e-17, 
    8.515048e-17, 8.515327e-17, 8.515948e-17, 8.516932e-17, 8.516566e-17, 
    8.517251e-17, 8.517385e-17, 8.51635e-17, 8.516975e-17, 8.514934e-17, 
    8.515252e-17, 8.515071e-17, 8.514353e-17, 8.516635e-17, 8.515455e-17, 
    8.517647e-17, 8.517008e-17, 8.518879e-17, 8.517936e-17, 8.519776e-17, 
    8.520539e-17, 8.521308e-17, 8.522151e-17, 8.514894e-17, 8.51465e-17, 
    8.515096e-17, 8.515695e-17, 8.516281e-17, 8.517045e-17, 8.517129e-17, 
    8.517269e-17, 8.517646e-17, 8.517958e-17, 8.517303e-17, 8.518037e-17, 
    8.515304e-17, 8.516743e-17, 8.514548e-17, 8.515193e-17, 8.515664e-17, 
    8.515468e-17, 8.516526e-17, 8.516772e-17, 8.517769e-17, 8.51726e-17, 
    8.520341e-17, 8.518974e-17, 8.52283e-17, 8.52174e-17, 8.514562e-17, 
    8.514898e-17, 8.516053e-17, 8.515505e-17, 8.517102e-17, 8.517491e-17, 
    8.517818e-17, 8.518218e-17, 8.518269e-17, 8.518507e-17, 8.518115e-17, 
    8.518496e-17, 8.517047e-17, 8.517695e-17, 8.515934e-17, 8.516355e-17, 
    8.516165e-17, 8.515948e-17, 8.516616e-17, 8.517311e-17, 8.517343e-17, 
    8.517563e-17, 8.518154e-17, 8.517109e-17, 8.520486e-17, 8.518367e-17, 
    8.515263e-17, 8.515887e-17, 8.515998e-17, 8.515752e-17, 8.517452e-17, 
    8.516833e-17, 8.518504e-17, 8.518055e-17, 8.518796e-17, 8.518426e-17, 
    8.518371e-17, 8.5179e-17, 8.517603e-17, 8.516857e-17, 8.516257e-17, 
    8.51579e-17, 8.5159e-17, 8.516413e-17, 8.517358e-17, 8.518266e-17, 
    8.518064e-17, 8.518739e-17, 8.516985e-17, 8.51771e-17, 8.517424e-17, 
    8.518174e-17, 8.516552e-17, 8.51788e-17, 8.516207e-17, 8.516357e-17, 
    8.51682e-17, 8.517748e-17, 8.51798e-17, 8.518195e-17, 8.518066e-17, 
    8.517385e-17, 8.517281e-17, 8.516814e-17, 8.516676e-17, 8.516325e-17, 
    8.516028e-17, 8.516296e-17, 8.516574e-17, 8.517392e-17, 8.518123e-17, 
    8.518926e-17, 8.51913e-17, 8.520026e-17, 8.519271e-17, 8.520494e-17, 
    8.519418e-17, 8.521302e-17, 8.517984e-17, 8.519422e-17, 8.516847e-17, 
    8.517128e-17, 8.517618e-17, 8.518782e-17, 8.518171e-17, 8.518894e-17, 
    8.517278e-17, 8.516423e-17, 8.516223e-17, 8.515815e-17, 8.516232e-17, 
    8.516199e-17, 8.516597e-17, 8.51647e-17, 8.517419e-17, 8.51691e-17, 
    8.518365e-17, 8.518892e-17, 8.520406e-17, 8.521328e-17, 8.522297e-17, 
    8.522716e-17, 8.522846e-17, 8.522898e-17 ;

 MEG_carene_3 =
  3.290387e-17, 3.29072e-17, 3.290657e-17, 3.290922e-17, 3.290778e-17, 
    3.290949e-17, 3.290458e-17, 3.290731e-17, 3.290558e-17, 3.290421e-17, 
    3.291429e-17, 3.290935e-17, 3.291973e-17, 3.291652e-17, 3.292469e-17, 
    3.291919e-17, 3.292582e-17, 3.29246e-17, 3.292843e-17, 3.292733e-17, 
    3.293209e-17, 3.292893e-17, 3.293467e-17, 3.293137e-17, 3.293186e-17, 
    3.292882e-17, 3.291041e-17, 3.291366e-17, 3.29102e-17, 3.291066e-17, 
    3.291047e-17, 3.290778e-17, 3.290638e-17, 3.290366e-17, 3.290417e-17, 
    3.290619e-17, 3.291088e-17, 3.290933e-17, 3.291336e-17, 3.291327e-17, 
    3.291773e-17, 3.291572e-17, 3.292327e-17, 3.292114e-17, 3.292738e-17, 
    3.29258e-17, 3.292729e-17, 3.292685e-17, 3.29273e-17, 3.292498e-17, 
    3.292597e-17, 3.292396e-17, 3.291608e-17, 3.291837e-17, 3.291151e-17, 
    3.290731e-17, 3.290469e-17, 3.290278e-17, 3.290304e-17, 3.290355e-17, 
    3.29062e-17, 3.290876e-17, 3.29107e-17, 3.291198e-17, 3.291326e-17, 
    3.291695e-17, 3.291906e-17, 3.292367e-17, 3.29229e-17, 3.292426e-17, 
    3.292564e-17, 3.292789e-17, 3.292753e-17, 3.292851e-17, 3.292426e-17, 
    3.292706e-17, 3.292244e-17, 3.292369e-17, 3.291338e-17, 3.290976e-17, 
    3.290803e-17, 3.290668e-17, 3.290325e-17, 3.290561e-17, 3.290467e-17, 
    3.290695e-17, 3.290836e-17, 3.290767e-17, 3.291202e-17, 3.291032e-17, 
    3.291918e-17, 3.291536e-17, 3.292548e-17, 3.292306e-17, 3.292607e-17, 
    3.292454e-17, 3.292714e-17, 3.292481e-17, 3.292889e-17, 3.292975e-17, 
    3.292916e-17, 3.293152e-17, 3.292467e-17, 3.292727e-17, 3.290764e-17, 
    3.290775e-17, 3.29083e-17, 3.29059e-17, 3.290576e-17, 3.290364e-17, 
    3.290555e-17, 3.290635e-17, 3.290846e-17, 3.290967e-17, 3.291083e-17, 
    3.29134e-17, 3.291623e-17, 3.292027e-17, 3.292321e-17, 3.292518e-17, 
    3.292399e-17, 3.292504e-17, 3.292386e-17, 3.292331e-17, 3.292941e-17, 
    3.292597e-17, 3.293118e-17, 3.293089e-17, 3.292852e-17, 3.293093e-17, 
    3.290783e-17, 3.290718e-17, 3.290487e-17, 3.290668e-17, 3.290341e-17, 
    3.290521e-17, 3.290623e-17, 3.29103e-17, 3.291125e-17, 3.291206e-17, 
    3.291372e-17, 3.291582e-17, 3.291949e-17, 3.292273e-17, 3.292573e-17, 
    3.292552e-17, 3.292559e-17, 3.292624e-17, 3.29246e-17, 3.292651e-17, 
    3.292681e-17, 3.292599e-17, 3.293086e-17, 3.292946e-17, 3.293089e-17, 
    3.292999e-17, 3.29074e-17, 3.29085e-17, 3.29079e-17, 3.290901e-17, 
    3.290821e-17, 3.291172e-17, 3.291277e-17, 3.291776e-17, 3.291576e-17, 
    3.2919e-17, 3.291611e-17, 3.291661e-17, 3.291901e-17, 3.291628e-17, 
    3.292251e-17, 3.29182e-17, 3.292627e-17, 3.292185e-17, 3.292654e-17, 
    3.292572e-17, 3.292709e-17, 3.29283e-17, 3.292985e-17, 3.293267e-17, 
    3.293203e-17, 3.293443e-17, 3.291016e-17, 3.291157e-17, 3.291149e-17, 
    3.291299e-17, 3.29141e-17, 3.291655e-17, 3.292044e-17, 3.291899e-17, 
    3.292169e-17, 3.292222e-17, 3.291814e-17, 3.29206e-17, 3.291255e-17, 
    3.29138e-17, 3.291309e-17, 3.291025e-17, 3.291926e-17, 3.29146e-17, 
    3.292325e-17, 3.292073e-17, 3.292812e-17, 3.29244e-17, 3.293166e-17, 
    3.293467e-17, 3.293771e-17, 3.294104e-17, 3.291238e-17, 3.291142e-17, 
    3.291319e-17, 3.291555e-17, 3.291786e-17, 3.292088e-17, 3.292121e-17, 
    3.292177e-17, 3.292325e-17, 3.292448e-17, 3.29219e-17, 3.29248e-17, 
    3.291401e-17, 3.291968e-17, 3.291102e-17, 3.291357e-17, 3.291543e-17, 
    3.291465e-17, 3.291883e-17, 3.29198e-17, 3.292374e-17, 3.292173e-17, 
    3.293389e-17, 3.292849e-17, 3.294372e-17, 3.293942e-17, 3.291108e-17, 
    3.29124e-17, 3.291696e-17, 3.29148e-17, 3.29211e-17, 3.292264e-17, 
    3.292393e-17, 3.292551e-17, 3.292571e-17, 3.292665e-17, 3.29251e-17, 
    3.292661e-17, 3.292089e-17, 3.292345e-17, 3.291649e-17, 3.291816e-17, 
    3.29174e-17, 3.291655e-17, 3.291918e-17, 3.292193e-17, 3.292206e-17, 
    3.292292e-17, 3.292526e-17, 3.292113e-17, 3.293446e-17, 3.29261e-17, 
    3.291384e-17, 3.291631e-17, 3.291675e-17, 3.291577e-17, 3.292248e-17, 
    3.292004e-17, 3.292664e-17, 3.292487e-17, 3.292779e-17, 3.292633e-17, 
    3.292611e-17, 3.292426e-17, 3.292309e-17, 3.292014e-17, 3.291777e-17, 
    3.291592e-17, 3.291636e-17, 3.291838e-17, 3.292211e-17, 3.29257e-17, 
    3.29249e-17, 3.292757e-17, 3.292064e-17, 3.292351e-17, 3.292238e-17, 
    3.292534e-17, 3.291893e-17, 3.292418e-17, 3.291757e-17, 3.291816e-17, 
    3.291999e-17, 3.292365e-17, 3.292457e-17, 3.292542e-17, 3.292491e-17, 
    3.292222e-17, 3.292181e-17, 3.291997e-17, 3.291942e-17, 3.291804e-17, 
    3.291686e-17, 3.291792e-17, 3.291902e-17, 3.292225e-17, 3.292513e-17, 
    3.292831e-17, 3.292911e-17, 3.293265e-17, 3.292967e-17, 3.29345e-17, 
    3.293025e-17, 3.293769e-17, 3.292458e-17, 3.293026e-17, 3.29201e-17, 
    3.292121e-17, 3.292314e-17, 3.292773e-17, 3.292533e-17, 3.292818e-17, 
    3.29218e-17, 3.291842e-17, 3.291763e-17, 3.291602e-17, 3.291767e-17, 
    3.291754e-17, 3.291911e-17, 3.291861e-17, 3.292236e-17, 3.292035e-17, 
    3.292609e-17, 3.292817e-17, 3.293415e-17, 3.293779e-17, 3.294161e-17, 
    3.294327e-17, 3.294378e-17, 3.294399e-17 ;

 MEG_ethanol =
  1.701311e-18, 1.701567e-18, 1.701518e-18, 1.701722e-18, 1.701611e-18, 
    1.701743e-18, 1.701365e-18, 1.701575e-18, 1.701442e-18, 1.701337e-18, 
    1.702113e-18, 1.701732e-18, 1.702531e-18, 1.702283e-18, 1.702912e-18, 
    1.702489e-18, 1.702998e-18, 1.702905e-18, 1.703199e-18, 1.703115e-18, 
    1.70348e-18, 1.703238e-18, 1.703679e-18, 1.703425e-18, 1.703463e-18, 
    1.703229e-18, 1.701813e-18, 1.702064e-18, 1.701797e-18, 1.701833e-18, 
    1.701818e-18, 1.701612e-18, 1.701504e-18, 1.701295e-18, 1.701334e-18, 
    1.701489e-18, 1.70185e-18, 1.701731e-18, 1.702041e-18, 1.702034e-18, 
    1.702377e-18, 1.702222e-18, 1.702803e-18, 1.702639e-18, 1.703119e-18, 
    1.702997e-18, 1.703112e-18, 1.703078e-18, 1.703112e-18, 1.702934e-18, 
    1.70301e-18, 1.702855e-18, 1.70225e-18, 1.702426e-18, 1.701899e-18, 
    1.701575e-18, 1.701373e-18, 1.701226e-18, 1.701247e-18, 1.701286e-18, 
    1.70149e-18, 1.701687e-18, 1.701836e-18, 1.701935e-18, 1.702033e-18, 
    1.702317e-18, 1.702479e-18, 1.702834e-18, 1.702774e-18, 1.702879e-18, 
    1.702985e-18, 1.703158e-18, 1.70313e-18, 1.703205e-18, 1.702879e-18, 
    1.703094e-18, 1.702739e-18, 1.702835e-18, 1.702042e-18, 1.701764e-18, 
    1.70163e-18, 1.701527e-18, 1.701263e-18, 1.701444e-18, 1.701372e-18, 
    1.701547e-18, 1.701656e-18, 1.701603e-18, 1.701937e-18, 1.701807e-18, 
    1.702488e-18, 1.702194e-18, 1.702973e-18, 1.702787e-18, 1.703018e-18, 
    1.702901e-18, 1.7031e-18, 1.702921e-18, 1.703235e-18, 1.7033e-18, 
    1.703255e-18, 1.703437e-18, 1.70291e-18, 1.70311e-18, 1.701601e-18, 
    1.701609e-18, 1.701651e-18, 1.701467e-18, 1.701456e-18, 1.701293e-18, 
    1.70144e-18, 1.701501e-18, 1.701664e-18, 1.701757e-18, 1.701846e-18, 
    1.702044e-18, 1.702262e-18, 1.702572e-18, 1.702798e-18, 1.70295e-18, 
    1.702858e-18, 1.702939e-18, 1.702848e-18, 1.702806e-18, 1.703274e-18, 
    1.70301e-18, 1.70341e-18, 1.703389e-18, 1.703206e-18, 1.703391e-18, 
    1.701615e-18, 1.701566e-18, 1.701387e-18, 1.701527e-18, 1.701275e-18, 
    1.701414e-18, 1.701493e-18, 1.701806e-18, 1.701879e-18, 1.701941e-18, 
    1.702068e-18, 1.70223e-18, 1.702512e-18, 1.702761e-18, 1.702992e-18, 
    1.702975e-18, 1.702981e-18, 1.703031e-18, 1.702905e-18, 1.703052e-18, 
    1.703075e-18, 1.703012e-18, 1.703386e-18, 1.703279e-18, 1.703388e-18, 
    1.703319e-18, 1.701582e-18, 1.701667e-18, 1.701621e-18, 1.701706e-18, 
    1.701645e-18, 1.701914e-18, 1.701995e-18, 1.702379e-18, 1.702226e-18, 
    1.702474e-18, 1.702252e-18, 1.70229e-18, 1.702475e-18, 1.702265e-18, 
    1.702744e-18, 1.702413e-18, 1.703033e-18, 1.702694e-18, 1.703054e-18, 
    1.702991e-18, 1.703097e-18, 1.703189e-18, 1.703309e-18, 1.703525e-18, 
    1.703476e-18, 1.70366e-18, 1.701795e-18, 1.701903e-18, 1.701897e-18, 
    1.702012e-18, 1.702097e-18, 1.702286e-18, 1.702585e-18, 1.702473e-18, 
    1.702681e-18, 1.702722e-18, 1.702408e-18, 1.702598e-18, 1.701978e-18, 
    1.702075e-18, 1.702019e-18, 1.701801e-18, 1.702494e-18, 1.702136e-18, 
    1.702802e-18, 1.702608e-18, 1.703176e-18, 1.702889e-18, 1.703448e-18, 
    1.703679e-18, 1.703913e-18, 1.704169e-18, 1.701966e-18, 1.701892e-18, 
    1.702027e-18, 1.702209e-18, 1.702387e-18, 1.702619e-18, 1.702644e-18, 
    1.702687e-18, 1.702801e-18, 1.702896e-18, 1.702697e-18, 1.70292e-18, 
    1.70209e-18, 1.702527e-18, 1.701861e-18, 1.702057e-18, 1.7022e-18, 
    1.70214e-18, 1.702461e-18, 1.702536e-18, 1.702839e-18, 1.702684e-18, 
    1.703619e-18, 1.703204e-18, 1.704375e-18, 1.704044e-18, 1.701865e-18, 
    1.701967e-18, 1.702318e-18, 1.702151e-18, 1.702636e-18, 1.702754e-18, 
    1.702853e-18, 1.702975e-18, 1.70299e-18, 1.703063e-18, 1.702944e-18, 
    1.703059e-18, 1.702619e-18, 1.702816e-18, 1.702281e-18, 1.702409e-18, 
    1.702352e-18, 1.702286e-18, 1.702489e-18, 1.702699e-18, 1.702709e-18, 
    1.702776e-18, 1.702956e-18, 1.702638e-18, 1.703663e-18, 1.70302e-18, 
    1.702078e-18, 1.702267e-18, 1.702301e-18, 1.702226e-18, 1.702742e-18, 
    1.702554e-18, 1.703062e-18, 1.702926e-18, 1.70315e-18, 1.703038e-18, 
    1.703021e-18, 1.702878e-18, 1.702788e-18, 1.702562e-18, 1.70238e-18, 
    1.702238e-18, 1.702271e-18, 1.702427e-18, 1.702714e-18, 1.702989e-18, 
    1.702928e-18, 1.703133e-18, 1.702601e-18, 1.702821e-18, 1.702734e-18, 
    1.702962e-18, 1.702469e-18, 1.702872e-18, 1.702364e-18, 1.70241e-18, 
    1.702551e-18, 1.702832e-18, 1.702903e-18, 1.702968e-18, 1.702929e-18, 
    1.702722e-18, 1.70269e-18, 1.702549e-18, 1.702507e-18, 1.7024e-18, 
    1.70231e-18, 1.702391e-18, 1.702476e-18, 1.702724e-18, 1.702946e-18, 
    1.70319e-18, 1.703252e-18, 1.703524e-18, 1.703294e-18, 1.703666e-18, 
    1.703339e-18, 1.703911e-18, 1.702904e-18, 1.70334e-18, 1.702559e-18, 
    1.702644e-18, 1.702793e-18, 1.703146e-18, 1.702961e-18, 1.70318e-18, 
    1.70269e-18, 1.70243e-18, 1.702369e-18, 1.702245e-18, 1.702372e-18, 
    1.702362e-18, 1.702483e-18, 1.702444e-18, 1.702733e-18, 1.702578e-18, 
    1.703019e-18, 1.70318e-18, 1.703639e-18, 1.703919e-18, 1.704213e-18, 
    1.70434e-18, 1.704379e-18, 1.704395e-18 ;

 MEG_formaldehyde =
  3.402622e-19, 3.403134e-19, 3.403037e-19, 3.403445e-19, 3.403222e-19, 
    3.403486e-19, 3.40273e-19, 3.40315e-19, 3.402885e-19, 3.402674e-19, 
    3.404225e-19, 3.403464e-19, 3.405061e-19, 3.404567e-19, 3.405824e-19, 
    3.404978e-19, 3.405997e-19, 3.40581e-19, 3.406398e-19, 3.40623e-19, 
    3.406961e-19, 3.406475e-19, 3.407358e-19, 3.40685e-19, 3.406925e-19, 
    3.406458e-19, 3.403627e-19, 3.404127e-19, 3.403595e-19, 3.403667e-19, 
    3.403637e-19, 3.403223e-19, 3.403008e-19, 3.40259e-19, 3.402667e-19, 
    3.402979e-19, 3.403699e-19, 3.403461e-19, 3.404081e-19, 3.404068e-19, 
    3.404753e-19, 3.404444e-19, 3.405606e-19, 3.405277e-19, 3.406237e-19, 
    3.405994e-19, 3.406224e-19, 3.406155e-19, 3.406225e-19, 3.405869e-19, 
    3.406021e-19, 3.40571e-19, 3.404499e-19, 3.404852e-19, 3.403798e-19, 
    3.40315e-19, 3.402747e-19, 3.402453e-19, 3.402494e-19, 3.402572e-19, 
    3.40298e-19, 3.403374e-19, 3.403672e-19, 3.403869e-19, 3.404065e-19, 
    3.404634e-19, 3.404958e-19, 3.405667e-19, 3.405548e-19, 3.405757e-19, 
    3.40597e-19, 3.406316e-19, 3.40626e-19, 3.40641e-19, 3.405758e-19, 
    3.406188e-19, 3.405478e-19, 3.405671e-19, 3.404084e-19, 3.403527e-19, 
    3.403261e-19, 3.403054e-19, 3.402526e-19, 3.402888e-19, 3.402744e-19, 
    3.403094e-19, 3.403312e-19, 3.403206e-19, 3.403875e-19, 3.403613e-19, 
    3.404977e-19, 3.404389e-19, 3.405945e-19, 3.405573e-19, 3.406036e-19, 
    3.405801e-19, 3.4062e-19, 3.405841e-19, 3.406469e-19, 3.406601e-19, 
    3.40651e-19, 3.406873e-19, 3.405821e-19, 3.40622e-19, 3.403201e-19, 
    3.403218e-19, 3.403302e-19, 3.402933e-19, 3.402913e-19, 3.402586e-19, 
    3.40288e-19, 3.403002e-19, 3.403327e-19, 3.403513e-19, 3.403692e-19, 
    3.404087e-19, 3.404523e-19, 3.405144e-19, 3.405597e-19, 3.405899e-19, 
    3.405716e-19, 3.405878e-19, 3.405696e-19, 3.405612e-19, 3.406548e-19, 
    3.40602e-19, 3.406821e-19, 3.406777e-19, 3.406412e-19, 3.406782e-19, 
    3.403231e-19, 3.403131e-19, 3.402775e-19, 3.403054e-19, 3.402551e-19, 
    3.402828e-19, 3.402985e-19, 3.403611e-19, 3.403757e-19, 3.403882e-19, 
    3.404136e-19, 3.404459e-19, 3.405024e-19, 3.405523e-19, 3.405984e-19, 
    3.405951e-19, 3.405962e-19, 3.406062e-19, 3.40581e-19, 3.406103e-19, 
    3.406149e-19, 3.406024e-19, 3.406771e-19, 3.406557e-19, 3.406776e-19, 
    3.406638e-19, 3.403165e-19, 3.403334e-19, 3.403242e-19, 3.403413e-19, 
    3.40329e-19, 3.403828e-19, 3.40399e-19, 3.404758e-19, 3.404451e-19, 
    3.404949e-19, 3.404504e-19, 3.404581e-19, 3.40495e-19, 3.40453e-19, 
    3.405489e-19, 3.404825e-19, 3.406066e-19, 3.405388e-19, 3.406107e-19, 
    3.405982e-19, 3.406193e-19, 3.406378e-19, 3.406617e-19, 3.407051e-19, 
    3.406951e-19, 3.40732e-19, 3.403589e-19, 3.403806e-19, 3.403793e-19, 
    3.404025e-19, 3.404195e-19, 3.404571e-19, 3.405169e-19, 3.404946e-19, 
    3.405363e-19, 3.405444e-19, 3.404816e-19, 3.405195e-19, 3.403956e-19, 
    3.404149e-19, 3.404039e-19, 3.403603e-19, 3.404989e-19, 3.404272e-19, 
    3.405603e-19, 3.405215e-19, 3.406351e-19, 3.405778e-19, 3.406896e-19, 
    3.407358e-19, 3.407825e-19, 3.408337e-19, 3.403931e-19, 3.403783e-19, 
    3.404054e-19, 3.404417e-19, 3.404774e-19, 3.405238e-19, 3.405289e-19, 
    3.405374e-19, 3.405602e-19, 3.405792e-19, 3.405394e-19, 3.40584e-19, 
    3.404181e-19, 3.405054e-19, 3.403721e-19, 3.404113e-19, 3.404399e-19, 
    3.40428e-19, 3.404923e-19, 3.405072e-19, 3.405677e-19, 3.405368e-19, 
    3.407238e-19, 3.406408e-19, 3.408749e-19, 3.408088e-19, 3.40373e-19, 
    3.403934e-19, 3.404635e-19, 3.404302e-19, 3.405272e-19, 3.405508e-19, 
    3.405707e-19, 3.40595e-19, 3.405981e-19, 3.406125e-19, 3.405887e-19, 
    3.406119e-19, 3.405238e-19, 3.405632e-19, 3.404563e-19, 3.404819e-19, 
    3.404703e-19, 3.404571e-19, 3.404977e-19, 3.405399e-19, 3.405419e-19, 
    3.405552e-19, 3.405911e-19, 3.405276e-19, 3.407327e-19, 3.40604e-19, 
    3.404156e-19, 3.404535e-19, 3.404602e-19, 3.404453e-19, 3.405484e-19, 
    3.405109e-19, 3.406123e-19, 3.405851e-19, 3.4063e-19, 3.406076e-19, 
    3.406042e-19, 3.405757e-19, 3.405577e-19, 3.405124e-19, 3.404759e-19, 
    3.404475e-19, 3.404542e-19, 3.404854e-19, 3.405427e-19, 3.405979e-19, 
    3.405856e-19, 3.406266e-19, 3.405201e-19, 3.405641e-19, 3.405468e-19, 
    3.405923e-19, 3.404938e-19, 3.405745e-19, 3.404729e-19, 3.40482e-19, 
    3.405101e-19, 3.405664e-19, 3.405805e-19, 3.405936e-19, 3.405857e-19, 
    3.405444e-19, 3.405381e-19, 3.405097e-19, 3.405014e-19, 3.404801e-19, 
    3.40462e-19, 3.404782e-19, 3.404951e-19, 3.405448e-19, 3.405892e-19, 
    3.406379e-19, 3.406503e-19, 3.407047e-19, 3.406589e-19, 3.407331e-19, 
    3.406678e-19, 3.407822e-19, 3.405807e-19, 3.40668e-19, 3.405118e-19, 
    3.405288e-19, 3.405585e-19, 3.406292e-19, 3.405921e-19, 3.40636e-19, 
    3.405379e-19, 3.404859e-19, 3.404738e-19, 3.404491e-19, 3.404744e-19, 
    3.404724e-19, 3.404966e-19, 3.404888e-19, 3.405465e-19, 3.405155e-19, 
    3.406039e-19, 3.406359e-19, 3.407278e-19, 3.407837e-19, 3.408425e-19, 
    3.40868e-19, 3.408758e-19, 3.408791e-19 ;

 MEG_isoprene =
  2.338708e-19, 2.339128e-19, 2.339048e-19, 2.339383e-19, 2.3392e-19, 
    2.339417e-19, 2.338796e-19, 2.339141e-19, 2.338923e-19, 2.33875e-19, 
    2.340023e-19, 2.339399e-19, 2.340709e-19, 2.340304e-19, 2.341335e-19, 
    2.340641e-19, 2.341477e-19, 2.341323e-19, 2.341806e-19, 2.341668e-19, 
    2.342267e-19, 2.341869e-19, 2.342593e-19, 2.342176e-19, 2.342238e-19, 
    2.341855e-19, 2.339532e-19, 2.339943e-19, 2.339506e-19, 2.339565e-19, 
    2.339541e-19, 2.339201e-19, 2.339025e-19, 2.338681e-19, 2.338745e-19, 
    2.339001e-19, 2.339592e-19, 2.339396e-19, 2.339905e-19, 2.339894e-19, 
    2.340456e-19, 2.340203e-19, 2.341156e-19, 2.340886e-19, 2.341674e-19, 
    2.341474e-19, 2.341663e-19, 2.341607e-19, 2.341664e-19, 2.341372e-19, 
    2.341496e-19, 2.341242e-19, 2.340248e-19, 2.340537e-19, 2.339672e-19, 
    2.339141e-19, 2.33881e-19, 2.338569e-19, 2.338603e-19, 2.338666e-19, 
    2.339002e-19, 2.339325e-19, 2.339569e-19, 2.339731e-19, 2.339892e-19, 
    2.340359e-19, 2.340624e-19, 2.341207e-19, 2.341108e-19, 2.34128e-19, 
    2.341455e-19, 2.341738e-19, 2.341693e-19, 2.341816e-19, 2.341281e-19, 
    2.341634e-19, 2.341051e-19, 2.341209e-19, 2.339908e-19, 2.33945e-19, 
    2.339232e-19, 2.339062e-19, 2.338629e-19, 2.338926e-19, 2.338808e-19, 
    2.339095e-19, 2.339274e-19, 2.339187e-19, 2.339736e-19, 2.339521e-19, 
    2.34064e-19, 2.340158e-19, 2.341435e-19, 2.341129e-19, 2.341509e-19, 
    2.341316e-19, 2.341644e-19, 2.341349e-19, 2.341864e-19, 2.341972e-19, 
    2.341898e-19, 2.342195e-19, 2.341332e-19, 2.34166e-19, 2.339183e-19, 
    2.339197e-19, 2.339266e-19, 2.338963e-19, 2.338946e-19, 2.338678e-19, 
    2.338919e-19, 2.33902e-19, 2.339287e-19, 2.339439e-19, 2.339586e-19, 
    2.33991e-19, 2.340268e-19, 2.340777e-19, 2.341149e-19, 2.341397e-19, 
    2.341246e-19, 2.341379e-19, 2.34123e-19, 2.341161e-19, 2.341929e-19, 
    2.341496e-19, 2.342152e-19, 2.342117e-19, 2.341818e-19, 2.342121e-19, 
    2.339207e-19, 2.339126e-19, 2.338833e-19, 2.339062e-19, 2.338649e-19, 
    2.338877e-19, 2.339005e-19, 2.339519e-19, 2.339639e-19, 2.339741e-19, 
    2.33995e-19, 2.340215e-19, 2.340679e-19, 2.341088e-19, 2.341466e-19, 
    2.341439e-19, 2.341448e-19, 2.34153e-19, 2.341324e-19, 2.341564e-19, 
    2.341602e-19, 2.341499e-19, 2.342111e-19, 2.341936e-19, 2.342116e-19, 
    2.342002e-19, 2.339153e-19, 2.339292e-19, 2.339216e-19, 2.339357e-19, 
    2.339256e-19, 2.339698e-19, 2.33983e-19, 2.34046e-19, 2.340208e-19, 
    2.340617e-19, 2.340252e-19, 2.340315e-19, 2.340618e-19, 2.340274e-19, 
    2.34106e-19, 2.340516e-19, 2.341533e-19, 2.340977e-19, 2.341567e-19, 
    2.341464e-19, 2.341638e-19, 2.34179e-19, 2.341985e-19, 2.342341e-19, 
    2.34226e-19, 2.342562e-19, 2.339501e-19, 2.339679e-19, 2.339669e-19, 
    2.339859e-19, 2.339998e-19, 2.340307e-19, 2.340798e-19, 2.340615e-19, 
    2.340957e-19, 2.341023e-19, 2.340508e-19, 2.340819e-19, 2.339802e-19, 
    2.339961e-19, 2.33987e-19, 2.339512e-19, 2.34065e-19, 2.340062e-19, 
    2.341154e-19, 2.340836e-19, 2.341767e-19, 2.341298e-19, 2.342214e-19, 
    2.342593e-19, 2.342976e-19, 2.343396e-19, 2.339782e-19, 2.339661e-19, 
    2.339883e-19, 2.340181e-19, 2.340473e-19, 2.340854e-19, 2.340896e-19, 
    2.340966e-19, 2.341153e-19, 2.341308e-19, 2.340982e-19, 2.341348e-19, 
    2.339987e-19, 2.340703e-19, 2.33961e-19, 2.339931e-19, 2.340166e-19, 
    2.340068e-19, 2.340595e-19, 2.340718e-19, 2.341215e-19, 2.340961e-19, 
    2.342495e-19, 2.341814e-19, 2.343734e-19, 2.343191e-19, 2.339617e-19, 
    2.339784e-19, 2.34036e-19, 2.340086e-19, 2.340882e-19, 2.341076e-19, 
    2.341239e-19, 2.341438e-19, 2.341463e-19, 2.341582e-19, 2.341387e-19, 
    2.341577e-19, 2.340855e-19, 2.341178e-19, 2.3403e-19, 2.34051e-19, 
    2.340416e-19, 2.340307e-19, 2.34064e-19, 2.340986e-19, 2.341002e-19, 
    2.341112e-19, 2.341406e-19, 2.340885e-19, 2.342567e-19, 2.341512e-19, 
    2.339966e-19, 2.340277e-19, 2.340332e-19, 2.34021e-19, 2.341056e-19, 
    2.340748e-19, 2.341581e-19, 2.341357e-19, 2.341726e-19, 2.341542e-19, 
    2.341514e-19, 2.34128e-19, 2.341132e-19, 2.340761e-19, 2.340461e-19, 
    2.340229e-19, 2.340283e-19, 2.340539e-19, 2.34101e-19, 2.341462e-19, 
    2.341362e-19, 2.341698e-19, 2.340824e-19, 2.341185e-19, 2.341043e-19, 
    2.341416e-19, 2.340608e-19, 2.34127e-19, 2.340436e-19, 2.340511e-19, 
    2.340742e-19, 2.341204e-19, 2.341319e-19, 2.341427e-19, 2.341362e-19, 
    2.341023e-19, 2.340971e-19, 2.340738e-19, 2.34067e-19, 2.340495e-19, 
    2.340347e-19, 2.34048e-19, 2.340619e-19, 2.341027e-19, 2.341391e-19, 
    2.341791e-19, 2.341892e-19, 2.342338e-19, 2.341962e-19, 2.342571e-19, 
    2.342035e-19, 2.342973e-19, 2.341322e-19, 2.342037e-19, 2.340755e-19, 
    2.340895e-19, 2.341139e-19, 2.341719e-19, 2.341415e-19, 2.341774e-19, 
    2.34097e-19, 2.340544e-19, 2.340444e-19, 2.340241e-19, 2.340449e-19, 
    2.340432e-19, 2.340631e-19, 2.340568e-19, 2.34104e-19, 2.340786e-19, 
    2.341511e-19, 2.341774e-19, 2.342527e-19, 2.342986e-19, 2.343468e-19, 
    2.343677e-19, 2.343742e-19, 2.343768e-19 ;

 MEG_methanol =
  5.849211e-17, 5.84976e-17, 5.849656e-17, 5.850093e-17, 5.849854e-17, 
    5.850138e-17, 5.849327e-17, 5.849778e-17, 5.849492e-17, 5.849267e-17, 
    5.850931e-17, 5.850114e-17, 5.851828e-17, 5.851298e-17, 5.852646e-17, 
    5.851739e-17, 5.852832e-17, 5.852631e-17, 5.853262e-17, 5.853082e-17, 
    5.853866e-17, 5.853345e-17, 5.854293e-17, 5.853747e-17, 5.853828e-17, 
    5.853327e-17, 5.850289e-17, 5.850826e-17, 5.850255e-17, 5.850331e-17, 
    5.8503e-17, 5.849856e-17, 5.849625e-17, 5.849176e-17, 5.849259e-17, 
    5.849594e-17, 5.850367e-17, 5.850111e-17, 5.850777e-17, 5.850762e-17, 
    5.851497e-17, 5.851165e-17, 5.852412e-17, 5.85206e-17, 5.85309e-17, 
    5.852828e-17, 5.853075e-17, 5.853002e-17, 5.853076e-17, 5.852695e-17, 
    5.852857e-17, 5.852525e-17, 5.851226e-17, 5.851603e-17, 5.850472e-17, 
    5.849778e-17, 5.849345e-17, 5.849029e-17, 5.849074e-17, 5.849157e-17, 
    5.849596e-17, 5.850018e-17, 5.850337e-17, 5.850549e-17, 5.85076e-17, 
    5.85137e-17, 5.851717e-17, 5.852478e-17, 5.85235e-17, 5.852575e-17, 
    5.852803e-17, 5.853174e-17, 5.853114e-17, 5.853276e-17, 5.852575e-17, 
    5.853037e-17, 5.852275e-17, 5.852482e-17, 5.850779e-17, 5.850182e-17, 
    5.849896e-17, 5.849674e-17, 5.849107e-17, 5.849497e-17, 5.849342e-17, 
    5.849718e-17, 5.849951e-17, 5.849837e-17, 5.850555e-17, 5.850274e-17, 
    5.851738e-17, 5.851106e-17, 5.852777e-17, 5.852377e-17, 5.852874e-17, 
    5.852622e-17, 5.85305e-17, 5.852665e-17, 5.853338e-17, 5.85348e-17, 
    5.853383e-17, 5.853772e-17, 5.852643e-17, 5.853072e-17, 5.849833e-17, 
    5.84985e-17, 5.84994e-17, 5.849545e-17, 5.849523e-17, 5.849172e-17, 
    5.849488e-17, 5.849619e-17, 5.849968e-17, 5.850167e-17, 5.850359e-17, 
    5.850783e-17, 5.851251e-17, 5.851917e-17, 5.852403e-17, 5.852727e-17, 
    5.85253e-17, 5.852704e-17, 5.852509e-17, 5.852419e-17, 5.853424e-17, 
    5.852857e-17, 5.853716e-17, 5.853669e-17, 5.853278e-17, 5.853675e-17, 
    5.849864e-17, 5.849757e-17, 5.849375e-17, 5.849674e-17, 5.849134e-17, 
    5.849432e-17, 5.8496e-17, 5.850272e-17, 5.850429e-17, 5.850562e-17, 
    5.850836e-17, 5.851182e-17, 5.851789e-17, 5.852323e-17, 5.852818e-17, 
    5.852783e-17, 5.852795e-17, 5.852901e-17, 5.852632e-17, 5.852946e-17, 
    5.852995e-17, 5.852861e-17, 5.853663e-17, 5.853434e-17, 5.853669e-17, 
    5.85352e-17, 5.849793e-17, 5.849974e-17, 5.849876e-17, 5.85006e-17, 
    5.849927e-17, 5.850505e-17, 5.850678e-17, 5.851502e-17, 5.851173e-17, 
    5.851707e-17, 5.85123e-17, 5.851313e-17, 5.851709e-17, 5.851259e-17, 
    5.852286e-17, 5.851575e-17, 5.852906e-17, 5.852178e-17, 5.85295e-17, 
    5.852816e-17, 5.853042e-17, 5.853241e-17, 5.853497e-17, 5.853962e-17, 
    5.853857e-17, 5.854252e-17, 5.850249e-17, 5.850481e-17, 5.850468e-17, 
    5.850716e-17, 5.850898e-17, 5.851302e-17, 5.851944e-17, 5.851705e-17, 
    5.852151e-17, 5.852239e-17, 5.851564e-17, 5.851971e-17, 5.850642e-17, 
    5.850849e-17, 5.850731e-17, 5.850263e-17, 5.85175e-17, 5.850981e-17, 
    5.852409e-17, 5.851993e-17, 5.853212e-17, 5.852597e-17, 5.853796e-17, 
    5.854293e-17, 5.854794e-17, 5.855343e-17, 5.850615e-17, 5.850457e-17, 
    5.850748e-17, 5.851138e-17, 5.851519e-17, 5.852017e-17, 5.852072e-17, 
    5.852163e-17, 5.852409e-17, 5.852612e-17, 5.852186e-17, 5.852663e-17, 
    5.850883e-17, 5.85182e-17, 5.85039e-17, 5.850811e-17, 5.851118e-17, 
    5.85099e-17, 5.851679e-17, 5.85184e-17, 5.852489e-17, 5.852157e-17, 
    5.854164e-17, 5.853274e-17, 5.855785e-17, 5.855075e-17, 5.8504e-17, 
    5.850619e-17, 5.851371e-17, 5.851014e-17, 5.852054e-17, 5.852307e-17, 
    5.852521e-17, 5.852781e-17, 5.852814e-17, 5.85297e-17, 5.852714e-17, 
    5.852963e-17, 5.852018e-17, 5.85244e-17, 5.851293e-17, 5.851568e-17, 
    5.851444e-17, 5.851302e-17, 5.851738e-17, 5.85219e-17, 5.852212e-17, 
    5.852354e-17, 5.85274e-17, 5.852059e-17, 5.854258e-17, 5.852878e-17, 
    5.850856e-17, 5.851263e-17, 5.851335e-17, 5.851175e-17, 5.852282e-17, 
    5.851879e-17, 5.852967e-17, 5.852675e-17, 5.853157e-17, 5.852917e-17, 
    5.852881e-17, 5.852574e-17, 5.852381e-17, 5.851895e-17, 5.851503e-17, 
    5.8512e-17, 5.851271e-17, 5.851605e-17, 5.852221e-17, 5.852812e-17, 
    5.852681e-17, 5.853121e-17, 5.851978e-17, 5.85245e-17, 5.852264e-17, 
    5.852753e-17, 5.851696e-17, 5.852562e-17, 5.851471e-17, 5.851569e-17, 
    5.851871e-17, 5.852475e-17, 5.852626e-17, 5.852767e-17, 5.852682e-17, 
    5.852239e-17, 5.852171e-17, 5.851866e-17, 5.851777e-17, 5.851548e-17, 
    5.851355e-17, 5.851529e-17, 5.85171e-17, 5.852243e-17, 5.852719e-17, 
    5.853243e-17, 5.853375e-17, 5.853959e-17, 5.853467e-17, 5.854264e-17, 
    5.853563e-17, 5.85479e-17, 5.852628e-17, 5.853565e-17, 5.851889e-17, 
    5.852071e-17, 5.85239e-17, 5.853149e-17, 5.852751e-17, 5.853221e-17, 
    5.852169e-17, 5.851611e-17, 5.851482e-17, 5.851216e-17, 5.851488e-17, 
    5.851466e-17, 5.851725e-17, 5.851642e-17, 5.852261e-17, 5.851929e-17, 
    5.852877e-17, 5.85322e-17, 5.854207e-17, 5.854807e-17, 5.855438e-17, 
    5.855711e-17, 5.855795e-17, 5.855829e-17 ;

 MEG_pinene_a =
  4.843399e-17, 4.843907e-17, 4.843811e-17, 4.844216e-17, 4.843995e-17, 
    4.844258e-17, 4.843506e-17, 4.843924e-17, 4.84366e-17, 4.843451e-17, 
    4.844992e-17, 4.844236e-17, 4.845823e-17, 4.845332e-17, 4.846582e-17, 
    4.845741e-17, 4.846754e-17, 4.846568e-17, 4.847152e-17, 4.846985e-17, 
    4.847712e-17, 4.84723e-17, 4.848108e-17, 4.847602e-17, 4.847677e-17, 
    4.847212e-17, 4.844397e-17, 4.844895e-17, 4.844366e-17, 4.844437e-17, 
    4.844407e-17, 4.843996e-17, 4.843783e-17, 4.843367e-17, 4.843444e-17, 
    4.843754e-17, 4.84447e-17, 4.844233e-17, 4.844849e-17, 4.844836e-17, 
    4.845517e-17, 4.845209e-17, 4.846365e-17, 4.846038e-17, 4.846993e-17, 
    4.846751e-17, 4.846979e-17, 4.846911e-17, 4.84698e-17, 4.846626e-17, 
    4.846777e-17, 4.846469e-17, 4.845265e-17, 4.845615e-17, 4.844567e-17, 
    4.843924e-17, 4.843523e-17, 4.843231e-17, 4.843272e-17, 4.843349e-17, 
    4.843755e-17, 4.844146e-17, 4.844442e-17, 4.844638e-17, 4.844834e-17, 
    4.845399e-17, 4.845721e-17, 4.846426e-17, 4.846307e-17, 4.846515e-17, 
    4.846727e-17, 4.847071e-17, 4.847015e-17, 4.847165e-17, 4.846516e-17, 
    4.846944e-17, 4.846237e-17, 4.846429e-17, 4.844852e-17, 4.844298e-17, 
    4.844034e-17, 4.843828e-17, 4.843303e-17, 4.843664e-17, 4.843521e-17, 
    4.843868e-17, 4.844085e-17, 4.843979e-17, 4.844644e-17, 4.844384e-17, 
    4.84574e-17, 4.845155e-17, 4.846702e-17, 4.846332e-17, 4.846792e-17, 
    4.846559e-17, 4.846956e-17, 4.846599e-17, 4.847223e-17, 4.847354e-17, 
    4.847264e-17, 4.847625e-17, 4.846579e-17, 4.846976e-17, 4.843975e-17, 
    4.843992e-17, 4.844075e-17, 4.843708e-17, 4.843688e-17, 4.843363e-17, 
    4.843655e-17, 4.843777e-17, 4.8441e-17, 4.844285e-17, 4.844463e-17, 
    4.844855e-17, 4.845289e-17, 4.845906e-17, 4.846356e-17, 4.846657e-17, 
    4.846474e-17, 4.846635e-17, 4.846454e-17, 4.846371e-17, 4.847303e-17, 
    4.846777e-17, 4.847573e-17, 4.84753e-17, 4.847167e-17, 4.847535e-17, 
    4.844004e-17, 4.843905e-17, 4.843551e-17, 4.843828e-17, 4.843328e-17, 
    4.843604e-17, 4.84376e-17, 4.844382e-17, 4.844527e-17, 4.844651e-17, 
    4.844904e-17, 4.845225e-17, 4.845787e-17, 4.846282e-17, 4.846741e-17, 
    4.846708e-17, 4.846719e-17, 4.846818e-17, 4.846568e-17, 4.84686e-17, 
    4.846905e-17, 4.846781e-17, 4.847524e-17, 4.847311e-17, 4.847529e-17, 
    4.847392e-17, 4.843938e-17, 4.844106e-17, 4.844015e-17, 4.844185e-17, 
    4.844062e-17, 4.844598e-17, 4.844758e-17, 4.845521e-17, 4.845217e-17, 
    4.845712e-17, 4.84527e-17, 4.845346e-17, 4.845713e-17, 4.845296e-17, 
    4.846248e-17, 4.845589e-17, 4.846822e-17, 4.846148e-17, 4.846863e-17, 
    4.846739e-17, 4.846949e-17, 4.847133e-17, 4.847371e-17, 4.847802e-17, 
    4.847703e-17, 4.84807e-17, 4.84436e-17, 4.844575e-17, 4.844563e-17, 
    4.844793e-17, 4.844962e-17, 4.845337e-17, 4.845931e-17, 4.845709e-17, 
    4.846123e-17, 4.846204e-17, 4.845579e-17, 4.845957e-17, 4.844725e-17, 
    4.844917e-17, 4.844807e-17, 4.844374e-17, 4.845751e-17, 4.845039e-17, 
    4.846362e-17, 4.845976e-17, 4.847106e-17, 4.846537e-17, 4.847648e-17, 
    4.848108e-17, 4.848572e-17, 4.849081e-17, 4.8447e-17, 4.844553e-17, 
    4.844822e-17, 4.845184e-17, 4.845538e-17, 4.845999e-17, 4.84605e-17, 
    4.846134e-17, 4.846362e-17, 4.84655e-17, 4.846155e-17, 4.846598e-17, 
    4.844948e-17, 4.845816e-17, 4.844491e-17, 4.844881e-17, 4.845165e-17, 
    4.845047e-17, 4.845686e-17, 4.845834e-17, 4.846436e-17, 4.846128e-17, 
    4.847988e-17, 4.847163e-17, 4.849491e-17, 4.848833e-17, 4.8445e-17, 
    4.844703e-17, 4.8454e-17, 4.845069e-17, 4.846033e-17, 4.846268e-17, 
    4.846465e-17, 4.846707e-17, 4.846737e-17, 4.846882e-17, 4.846645e-17, 
    4.846875e-17, 4.846e-17, 4.846391e-17, 4.845328e-17, 4.845582e-17, 
    4.845468e-17, 4.845337e-17, 4.84574e-17, 4.846159e-17, 4.846179e-17, 
    4.846312e-17, 4.846668e-17, 4.846037e-17, 4.848076e-17, 4.846797e-17, 
    4.844923e-17, 4.8453e-17, 4.845367e-17, 4.845218e-17, 4.846244e-17, 
    4.845871e-17, 4.846879e-17, 4.846609e-17, 4.847055e-17, 4.846832e-17, 
    4.846799e-17, 4.846515e-17, 4.846336e-17, 4.845886e-17, 4.845523e-17, 
    4.845241e-17, 4.845307e-17, 4.845617e-17, 4.846188e-17, 4.846736e-17, 
    4.846614e-17, 4.847022e-17, 4.845963e-17, 4.8464e-17, 4.846228e-17, 
    4.846681e-17, 4.845701e-17, 4.846503e-17, 4.845493e-17, 4.845583e-17, 
    4.845863e-17, 4.846423e-17, 4.846563e-17, 4.846693e-17, 4.846615e-17, 
    4.846204e-17, 4.846141e-17, 4.845859e-17, 4.845776e-17, 4.845564e-17, 
    4.845384e-17, 4.845546e-17, 4.845714e-17, 4.846208e-17, 4.846649e-17, 
    4.847134e-17, 4.847257e-17, 4.847799e-17, 4.847342e-17, 4.848081e-17, 
    4.847431e-17, 4.848568e-17, 4.846565e-17, 4.847433e-17, 4.845879e-17, 
    4.846049e-17, 4.846345e-17, 4.847047e-17, 4.846679e-17, 4.847115e-17, 
    4.84614e-17, 4.845623e-17, 4.845503e-17, 4.845256e-17, 4.845508e-17, 
    4.845488e-17, 4.845729e-17, 4.845652e-17, 4.846225e-17, 4.845917e-17, 
    4.846795e-17, 4.847114e-17, 4.848028e-17, 4.848584e-17, 4.849169e-17, 
    4.849422e-17, 4.8495e-17, 4.849532e-17 ;

 MEG_thujene_a =
  1.221556e-18, 1.22168e-18, 1.221656e-18, 1.221755e-18, 1.221701e-18, 
    1.221765e-18, 1.221582e-18, 1.221684e-18, 1.22162e-18, 1.221569e-18, 
    1.221943e-18, 1.22176e-18, 1.222145e-18, 1.222026e-18, 1.222329e-18, 
    1.222125e-18, 1.222371e-18, 1.222326e-18, 1.222468e-18, 1.222427e-18, 
    1.222604e-18, 1.222487e-18, 1.2227e-18, 1.222577e-18, 1.222595e-18, 
    1.222482e-18, 1.221799e-18, 1.22192e-18, 1.221791e-18, 1.221808e-18, 
    1.221801e-18, 1.221701e-18, 1.22165e-18, 1.221549e-18, 1.221567e-18, 
    1.221642e-18, 1.221816e-18, 1.221759e-18, 1.221909e-18, 1.221905e-18, 
    1.222071e-18, 1.221996e-18, 1.222277e-18, 1.222197e-18, 1.222429e-18, 
    1.22237e-18, 1.222426e-18, 1.222409e-18, 1.222426e-18, 1.22234e-18, 
    1.222377e-18, 1.222302e-18, 1.222009e-18, 1.222094e-18, 1.22184e-18, 
    1.221684e-18, 1.221586e-18, 1.221515e-18, 1.221526e-18, 1.221544e-18, 
    1.221643e-18, 1.221738e-18, 1.22181e-18, 1.221857e-18, 1.221905e-18, 
    1.222042e-18, 1.22212e-18, 1.222291e-18, 1.222263e-18, 1.222313e-18, 
    1.222364e-18, 1.222448e-18, 1.222434e-18, 1.222471e-18, 1.222313e-18, 
    1.222417e-18, 1.222246e-18, 1.222292e-18, 1.221909e-18, 1.221775e-18, 
    1.22171e-18, 1.221661e-18, 1.221533e-18, 1.221621e-18, 1.221586e-18, 
    1.22167e-18, 1.221723e-18, 1.221697e-18, 1.221859e-18, 1.221795e-18, 
    1.222125e-18, 1.221983e-18, 1.222358e-18, 1.222269e-18, 1.22238e-18, 
    1.222324e-18, 1.22242e-18, 1.222333e-18, 1.222485e-18, 1.222517e-18, 
    1.222495e-18, 1.222583e-18, 1.222328e-18, 1.222425e-18, 1.221696e-18, 
    1.2217e-18, 1.22172e-18, 1.221632e-18, 1.221627e-18, 1.221548e-18, 
    1.221619e-18, 1.221648e-18, 1.221727e-18, 1.221771e-18, 1.221815e-18, 
    1.22191e-18, 1.222015e-18, 1.222165e-18, 1.222274e-18, 1.222347e-18, 
    1.222303e-18, 1.222342e-18, 1.222298e-18, 1.222278e-18, 1.222504e-18, 
    1.222376e-18, 1.22257e-18, 1.22256e-18, 1.222471e-18, 1.222561e-18, 
    1.221703e-18, 1.221679e-18, 1.221593e-18, 1.221661e-18, 1.221539e-18, 
    1.221606e-18, 1.221644e-18, 1.221795e-18, 1.22183e-18, 1.22186e-18, 
    1.221922e-18, 1.222e-18, 1.222136e-18, 1.222256e-18, 1.222368e-18, 
    1.22236e-18, 1.222363e-18, 1.222387e-18, 1.222326e-18, 1.222397e-18, 
    1.222408e-18, 1.222378e-18, 1.222558e-18, 1.222506e-18, 1.222559e-18, 
    1.222526e-18, 1.221687e-18, 1.221728e-18, 1.221706e-18, 1.221747e-18, 
    1.221717e-18, 1.221847e-18, 1.221886e-18, 1.222072e-18, 1.221998e-18, 
    1.222118e-18, 1.222011e-18, 1.222029e-18, 1.222118e-18, 1.222017e-18, 
    1.222248e-18, 1.222088e-18, 1.222388e-18, 1.222224e-18, 1.222398e-18, 
    1.222367e-18, 1.222418e-18, 1.222463e-18, 1.222521e-18, 1.222625e-18, 
    1.222602e-18, 1.222691e-18, 1.22179e-18, 1.221842e-18, 1.221839e-18, 
    1.221895e-18, 1.221936e-18, 1.222027e-18, 1.222171e-18, 1.222117e-18, 
    1.222218e-18, 1.222238e-18, 1.222086e-18, 1.222177e-18, 1.221878e-18, 
    1.221925e-18, 1.221898e-18, 1.221793e-18, 1.222128e-18, 1.221955e-18, 
    1.222276e-18, 1.222182e-18, 1.222457e-18, 1.222318e-18, 1.222588e-18, 
    1.2227e-18, 1.222813e-18, 1.222936e-18, 1.221872e-18, 1.221837e-18, 
    1.221902e-18, 1.22199e-18, 1.222076e-18, 1.222188e-18, 1.2222e-18, 
    1.22222e-18, 1.222276e-18, 1.222321e-18, 1.222225e-18, 1.222333e-18, 
    1.221933e-18, 1.222143e-18, 1.221822e-18, 1.221916e-18, 1.221985e-18, 
    1.221956e-18, 1.222112e-18, 1.222148e-18, 1.222294e-18, 1.222219e-18, 
    1.222671e-18, 1.22247e-18, 1.223036e-18, 1.222876e-18, 1.221824e-18, 
    1.221873e-18, 1.222042e-18, 1.221962e-18, 1.222196e-18, 1.222253e-18, 
    1.222301e-18, 1.22236e-18, 1.222367e-18, 1.222402e-18, 1.222345e-18, 
    1.2224e-18, 1.222188e-18, 1.222283e-18, 1.222025e-18, 1.222086e-18, 
    1.222059e-18, 1.222027e-18, 1.222125e-18, 1.222227e-18, 1.222231e-18, 
    1.222264e-18, 1.22235e-18, 1.222197e-18, 1.222692e-18, 1.222381e-18, 
    1.221927e-18, 1.222018e-18, 1.222034e-18, 1.221998e-18, 1.222247e-18, 
    1.222156e-18, 1.222402e-18, 1.222336e-18, 1.222444e-18, 1.22239e-18, 
    1.222382e-18, 1.222313e-18, 1.222269e-18, 1.22216e-18, 1.222072e-18, 
    1.222004e-18, 1.22202e-18, 1.222095e-18, 1.222233e-18, 1.222367e-18, 
    1.222337e-18, 1.222436e-18, 1.222179e-18, 1.222285e-18, 1.222243e-18, 
    1.222353e-18, 1.222115e-18, 1.22231e-18, 1.222065e-18, 1.222087e-18, 
    1.222155e-18, 1.222291e-18, 1.222325e-18, 1.222356e-18, 1.222337e-18, 
    1.222237e-18, 1.222222e-18, 1.222154e-18, 1.222134e-18, 1.222082e-18, 
    1.222038e-18, 1.222078e-18, 1.222119e-18, 1.222238e-18, 1.222346e-18, 
    1.222463e-18, 1.222493e-18, 1.222625e-18, 1.222514e-18, 1.222693e-18, 
    1.222535e-18, 1.222812e-18, 1.222325e-18, 1.222536e-18, 1.222159e-18, 
    1.2222e-18, 1.222272e-18, 1.222442e-18, 1.222353e-18, 1.222459e-18, 
    1.222222e-18, 1.222096e-18, 1.222067e-18, 1.222007e-18, 1.222068e-18, 
    1.222064e-18, 1.222122e-18, 1.222103e-18, 1.222242e-18, 1.222168e-18, 
    1.222381e-18, 1.222458e-18, 1.22268e-18, 1.222815e-18, 1.222957e-18, 
    1.223019e-18, 1.223038e-18, 1.223046e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  2.280031e-25, 2.389912e-25, -1.510863e-25, 3.433782e-25, -1.043869e-25, 
    -3.40631e-25, -2.966786e-25, -2.527262e-25, 1.098811e-25, -4.230417e-25, 
    -6.098394e-25, 7.142273e-26, 2.774496e-25, -5.6314e-25, 5.136937e-25, 
    -1.428452e-25, 2.747107e-27, 2.527264e-25, 1.620745e-25, -5.60393e-25, 
    -6.345626e-25, -2.087738e-25, 1.346043e-25, -3.653542e-25, 8.241083e-26, 
    6.592867e-26, -5.768751e-25, -2.170149e-25, 4.230419e-25, 1.977859e-25, 
    -3.323899e-25, -3.159078e-25, -1.455922e-25, -3.845826e-26, 
    -2.554732e-25, -5.823692e-25, 8.515785e-26, 2.197628e-26, -7.691661e-26, 
    -1.373504e-26, -2.637143e-25, -1.318571e-25, 1.730626e-25, 2.747107e-27, 
    2.582204e-25, 3.928246e-25, -3.021719e-26, 2.362442e-25, 2.060269e-25, 
    -1.565803e-25, 3.873306e-25, -7.142256e-26, -1.977857e-25, -6.345626e-25, 
    -1.071339e-25, -1.895446e-25, 3.076668e-25, 1.977859e-25, 5.52152e-25, 
    3.26896e-25, -3.516191e-25, -1.15375e-25, -2.417381e-25, 2.829436e-25, 
    7.691677e-26, 1.538335e-25, 1.730626e-25, -4.56006e-25, 8.515785e-26, 
    -3.049197e-25, -4.669934e-26, -5.411638e-25, -8.240992e-27, -3.46125e-25, 
    -5.219339e-26, 4.010657e-25, -1.20869e-25, -2.527262e-25, -8.515768e-26, 
    -4.724882e-25, 1.840507e-25, -2.472314e-26, 6.592867e-26, -2.747016e-26, 
    -1.538333e-25, 2.527264e-25, -2.527262e-25, -2.911845e-25, -1.538333e-25, 
    -2.746942e-27, 7.059854e-25, -8.790471e-26, -1.400982e-25, 8.241083e-26, 
    7.416975e-26, -2.554732e-25, -1.648207e-26, 5.76876e-26, -3.131607e-25, 
    3.351371e-25, -2.746942e-27, -8.790471e-26, 1.922918e-25, 1.455924e-25, 
    1.785567e-25, 3.296431e-25, 1.346043e-25, -3.873304e-25, 5.76876e-26, 
    1.0164e-25, -3.653542e-25, -6.043446e-26, 2.225091e-25, -1.346041e-25, 
    -3.186548e-25, -1.373504e-26, 2.08774e-25, 7.96638e-26, -1.400982e-25, 
    1.895448e-25, 3.626074e-25, -5.411638e-25, 1.263632e-25, -2.499792e-25, 
    -1.620744e-25, -4.669934e-26, 8.515785e-26, -2.36244e-25, -1.593274e-25, 
    -4.202947e-25, -4.367769e-25, -1.291101e-25, -3.296421e-26, 
    -7.691661e-26, -4.697411e-25, -1.291101e-25, -8.240992e-27, 
    -2.499792e-25, 3.296438e-26, 3.955716e-25, -2.197619e-25, 1.483394e-25, 
    1.648223e-26, 1.538335e-25, -1.043869e-25, -2.032798e-25, -1.730625e-25, 
    1.373521e-26, -1.318571e-25, -8.240992e-27, 3.873306e-25, -1.867976e-25, 
    -1.648207e-26, -1.291101e-25, -9.889281e-26, -1.510863e-25, 
    -5.768744e-26, -3.214018e-25, -2.582203e-25, 3.21402e-25, -6.318148e-26, 
    3.708484e-25, -3.900774e-25, 3.406311e-25, -2.197612e-26, -1.977857e-25, 
    -4.120529e-26, -3.076667e-25, -1.538333e-25, -3.626072e-25, 8.79048e-25, 
    -6.318148e-26, 7.96638e-26, -7.966364e-26, -1.648214e-25, -4.093066e-25, 
    1.785567e-25, 8.790487e-26, -1.455922e-25, -5.521519e-25, 1.895448e-25, 
    -2.087738e-25, -4.395239e-25, 1.236162e-25, 2.225091e-25, -2.609673e-25, 
    -1.071339e-25, -1.043869e-25, 1.236162e-25, 3.296431e-25, -1.043869e-25, 
    -9.889281e-26, 5.961045e-25, 2.692085e-25, 6.043463e-26, 3.21402e-25, 
    -1.098809e-25, -7.416958e-26, 2.225091e-25, 2.197628e-26, 6.812622e-25, 
    8.241157e-27, -3.790893e-25, -4.065596e-25, 2.362442e-25, -4.669934e-26, 
    7.96638e-26, -3.214018e-25, 3.845843e-26, -4.175477e-25, 1.208692e-25, 
    -6.675269e-25, 1.263632e-25, 2.334972e-25, 4.038127e-25, 1.922918e-25, 
    2.14268e-25, -2.499792e-25, -3.296421e-26, 3.18655e-25, -7.719139e-25, 
    1.648223e-26, 2.362442e-25, 3.845843e-26, 9.614595e-26, -1.318571e-25, 
    1.785567e-25, -9.339876e-26, -2.225089e-25, 3.296438e-26, 1.867978e-25, 
    -3.681012e-25, 5.494132e-27, -2.28003e-25, 2.637145e-25, 2.197621e-25, 
    4.120545e-26, 1.373513e-25, -1.977857e-25, -3.626072e-25, -1.15375e-25, 
    -6.043446e-26, -6.867554e-26, 1.648216e-25, -1.593274e-25, -1.922909e-26, 
    -6.592851e-26, -9.339876e-26, 3.461252e-25, 3.296431e-25, -1.20869e-25, 
    8.257549e-32, -4.752352e-25, -1.400982e-25, 4.3403e-25, 3.21402e-25, 
    -1.648207e-26, -2.774494e-25, 5.109467e-25, -4.175477e-25, -1.510863e-25, 
    5.219355e-26, -1.895446e-25, 1.153751e-25, 3.296438e-26, 1.098811e-25, 
    -7.416958e-26, -4.669934e-26, -2.33497e-25, 5.219348e-25, 2.417383e-25, 
    -3.571124e-26, 2.444853e-25, -2.36244e-25, 2.032799e-25, -3.955715e-25, 
    -1.318571e-25, -3.351369e-25, -6.043446e-26, 2.472331e-26, 2.389912e-25, 
    -3.571124e-26, 3.873306e-25, 1.538335e-25, -1.950387e-25, -3.021727e-25, 
    -2.911845e-25, -2.115208e-25, -2.087738e-25, -4.148007e-25, 
    -9.065174e-26, -6.043446e-26, -3.37884e-25, -2.747016e-26, 1.730626e-25, 
    -4.312828e-25, -1.455922e-25, -2.087738e-25, -6.318148e-26, 
    -1.400982e-25, -1.703155e-25, 1.510864e-25, -8.240992e-27, 9.889298e-26, 
    7.96638e-26, -1.400982e-25, 6.318165e-26, 4.065598e-25, 5.027056e-25, 
    -7.416958e-26, -2.142679e-25, 8.257342e-32, 1.373521e-26, -1.895446e-25, 
    8.515785e-26, -1.867976e-25, -3.241488e-25, -2.197612e-26, -1.098809e-25, 
    -1.346041e-25, 2.032799e-25, 3.57114e-26, 1.758097e-25, 6.86757e-26, 
    1.181221e-25, -1.867976e-25, -4.862233e-25, -3.214018e-25, 4.999586e-25, 
    1.181221e-25, -3.845826e-26, 3.845843e-26, -1.455922e-25, -1.098802e-26, 
    1.510864e-25, -1.098809e-25, -2.609673e-25, 3.296438e-26 ;

 M_LITR2C_TO_LEACHING =
  2.472328e-26, -1.043869e-25, -2.087738e-25, -2.362441e-25, -6.318152e-26, 
    7.966377e-26, 2.197625e-26, 2.747078e-27, 5.351469e-32, -2.142679e-25, 
    -1.291101e-25, 1.373513e-25, -1.263631e-25, 1.346043e-25, -4.724882e-25, 
    -3.076667e-25, 7.966377e-26, 1.04387e-25, 7.691675e-26, -3.571127e-26, 
    8.790485e-26, -2.74702e-26, -3.35137e-25, -1.758095e-25, -6.043449e-26, 
    -1.813036e-25, 4.94465e-26, -1.18122e-25, -1.785566e-25, 8.790485e-26, 
    -3.845829e-26, -1.428452e-25, -2.939316e-25, 6.592865e-26, -9.065177e-26, 
    8.24108e-26, 5.494055e-26, -1.098809e-25, -2.499792e-25, 5.768757e-26, 
    4.395245e-26, -1.593274e-25, -8.790474e-26, 2.74703e-26, -6.043449e-26, 
    -1.15375e-25, -3.461251e-25, -4.340298e-25, 8.515782e-26, 1.565805e-25, 
    -5.219342e-26, -1.18122e-25, -1.263631e-25, -3.049197e-25, -2.664613e-25, 
    5.494103e-27, -1.263631e-25, 4.669947e-26, -2.087738e-25, -1.263631e-25, 
    -5.494044e-26, -3.845829e-26, -2.444852e-25, -7.416961e-26, 
    -1.867976e-25, 6.592865e-26, 4.477651e-25, 4.395245e-26, -1.813036e-25, 
    3.021728e-25, 1.785567e-25, 1.126281e-25, 3.571138e-26, 1.648215e-25, 
    -3.571127e-26, -2.032798e-25, 4.395245e-26, -1.510863e-25, -4.395234e-26, 
    -1.785566e-25, 1.648215e-25, 2.444853e-25, -2.74702e-26, 1.538334e-25, 
    1.098815e-26, 9.065187e-26, -1.071339e-25, -1.785566e-25, -2.966786e-25, 
    -2.609673e-25, 2.472328e-26, 9.339889e-26, -1.291101e-25, 1.098815e-26, 
    1.922923e-26, 2.389912e-25, -1.977857e-25, -5.493996e-27, -1.373512e-25, 
    -3.296424e-26, -6.592854e-26, 6.592865e-26, -1.593274e-25, 3.021728e-25, 
    1.428453e-25, 1.483394e-25, -7.966367e-26, 1.098815e-26, 1.483394e-25, 
    1.09881e-25, 7.691675e-26, 7.691675e-26, -2.554732e-25, -1.12628e-25, 
    1.922923e-26, 3.461252e-25, -1.593274e-25, -2.362441e-25, -2.197614e-26, 
    -1.648209e-26, -9.614581e-26, -2.142679e-25, -3.021722e-26, 
    -1.620744e-25, -7.416961e-26, 2.747025e-25, -2.087738e-25, -3.900775e-25, 
    9.889295e-26, 4.395245e-26, 1.291102e-25, -1.373512e-25, 1.64822e-26, 
    7.691675e-26, 3.021733e-26, -1.538333e-25, 1.64822e-26, -9.065177e-26, 
    1.126281e-25, -3.845829e-26, 8.790485e-26, -1.620744e-25, -2.444852e-25, 
    1.483394e-25, 9.889295e-26, 7.691675e-26, -1.483393e-25, 1.208691e-25, 
    -8.515771e-26, -2.032798e-25, -3.845829e-26, 4.94465e-26, -6.043449e-26, 
    -5.493996e-27, -1.785566e-25, 1.318572e-25, -2.664613e-25, 1.785567e-25, 
    -2.28003e-25, -8.241069e-26, -1.538333e-25, -2.032798e-25, -7.966367e-26, 
    5.351449e-32, -2.74702e-26, -2.747024e-25, -6.867557e-26, -1.20869e-25, 
    1.0164e-25, 2.417382e-25, -1.977857e-25, -4.120532e-26, -3.900775e-25, 
    -1.867976e-25, 1.593275e-25, 5.494103e-27, 2.14268e-25, -2.74702e-26, 
    -2.197614e-26, -2.334971e-25, 2.087739e-25, 3.296435e-26, -1.620744e-25, 
    -5.493996e-27, 6.867567e-26, -1.373512e-25, -8.241021e-27, 1.098815e-26, 
    3.84584e-26, 7.416973e-26, 4.395245e-26, 3.296435e-26, -7.142259e-26, 
    3.296435e-26, -5.494044e-26, 1.098815e-26, 2.74703e-26, -2.362441e-25, 
    6.04346e-26, 9.339889e-26, -2.692084e-25, -6.318152e-26, -2.005328e-25, 
    2.060269e-25, -1.15375e-25, -6.592854e-26, -6.592854e-26, 9.065187e-26, 
    -1.20869e-25, -8.241069e-26, 1.318572e-25, -9.889284e-26, 5.494055e-26, 
    -1.15375e-25, -1.428452e-25, -1.236161e-25, -5.493996e-27, -4.175477e-25, 
    -1.758095e-25, 2.966787e-25, -5.494044e-26, -2.911846e-25, 1.64822e-26, 
    1.565805e-25, -1.098805e-26, -2.444852e-25, -1.20869e-25, -2.417381e-25, 
    -1.428452e-25, 1.126281e-25, -2.28003e-25, 1.126281e-25, 8.24108e-26, 
    6.867567e-26, 8.24108e-26, -7.966367e-26, -3.571127e-26, 9.065187e-26, 
    -6.867557e-26, 6.04346e-26, 2.527263e-25, -3.186548e-25, -2.115208e-25, 
    2.11521e-25, -1.373507e-26, 4.395245e-26, -4.669937e-26, 8.790485e-26, 
    -2.911846e-25, 1.208691e-25, 2.417382e-25, -1.730625e-25, 3.104139e-25, 
    -5.219342e-26, -8.241069e-26, 4.120543e-26, -1.098805e-26, -1.922912e-26, 
    -2.197619e-25, 6.318163e-26, 6.318163e-26, -2.389911e-25, -3.323899e-25, 
    -7.691664e-26, -1.15375e-25, -7.142259e-26, -6.867557e-26, 2.554734e-25, 
    6.04346e-26, -1.565804e-25, -3.021722e-26, -3.43378e-25, 2.637144e-25, 
    -1.373512e-25, 2.252561e-25, -4.395234e-26, 4.94465e-26, 5.494103e-27, 
    -2.692084e-25, -2.005328e-25, 5.219352e-26, -2.334971e-25, 1.208691e-25, 
    2.747078e-27, 1.510864e-25, -6.043449e-26, 3.296435e-26, 7.14227e-26, 
    -9.339879e-26, 4.395245e-26, 1.09881e-25, -1.895447e-25, -1.373512e-25, 
    1.895448e-25, -7.691664e-26, 2.197625e-26, -3.735953e-25, -1.15375e-25, 
    4.669947e-26, -4.120532e-26, -1.098809e-25, -3.571127e-26, 5.768757e-26, 
    -4.944639e-26, -2.884375e-25, 5.351432e-32, -7.966367e-26, -6.867557e-26, 
    -1.043869e-25, -1.236161e-25, 1.758096e-25, 1.373518e-26, 6.592865e-26, 
    1.510864e-25, -6.592854e-26, 3.021733e-26, -3.021722e-26, 1.07134e-25, 
    -6.592854e-26, 2.197625e-26, 2.664615e-25, 2.499793e-25, 1.318572e-25, 
    -1.648214e-25, -1.730625e-25, 1.098815e-26, 1.0164e-25, 7.14227e-26, 
    2.582204e-25, -9.339879e-26, 2.11521e-25, 1.428453e-25, -1.15375e-25, 
    -1.648209e-26, 7.14227e-26, 2.417382e-25, 8.241128e-27, -1.400982e-25 ;

 M_LITR3C_TO_LEACHING =
  8.241101e-27, -7.416964e-26, -4.944642e-26, 4.12054e-26, -1.18122e-25, 
    -3.57113e-26, -1.37351e-26, 9.614589e-26, -7.142262e-26, -1.771831e-25, 
    -4.669939e-26, 2.197622e-26, 1.002664e-25, 6.180808e-26, 9.889292e-26, 
    -1.497128e-25, 9.065185e-26, -1.414718e-25, 4.669945e-26, 1.373539e-27, 
    7.829024e-26, -3.845832e-26, -1.140015e-25, 1.098813e-26, 1.236161e-25, 
    -1.057604e-25, -9.751935e-26, -3.159076e-26, -1.15375e-25, 6.730214e-26, 
    8.241101e-27, 3.296432e-26, 1.153751e-25, -4.120511e-27, -4.395237e-26, 
    -8.241071e-26, 1.181221e-25, -5.906101e-26, -4.120511e-27, 1.373513e-25, 
    -1.318572e-25, -1.703155e-25, 2.747028e-26, -2.334968e-26, -4.807291e-26, 
    -6.180803e-26, 3.159081e-26, -1.37351e-26, -1.469658e-25, -3.708481e-26, 
    -1.373512e-25, -1.098807e-26, 5.906106e-26, -1.249896e-25, 1.373515e-26, 
    -9.889287e-26, -5.494023e-27, -1.098807e-26, -7.691667e-26, 1.167486e-25, 
    -2.197617e-26, -5.219344e-26, 5.494076e-27, 3.983189e-26, -7.691667e-26, 
    -2.746998e-27, -3.708481e-26, -6.867559e-26, -1.37351e-26, -6.592857e-26, 
    1.60701e-25, 3.159081e-26, -1.09881e-25, -3.708481e-26, -1.098807e-26, 
    1.469658e-25, -9.20253e-26, -2.197617e-26, 3.433784e-26, -9.20253e-26, 
    -1.057604e-25, -2.747022e-26, 1.483394e-25, -1.758096e-25, -9.614584e-26, 
    -2.334968e-26, 2.472325e-26, -7.416964e-26, 8.241101e-27, -1.785563e-26, 
    -8.927828e-26, 2.747052e-27, 6.867565e-26, -4.944642e-26, 6.455511e-26, 
    7.416969e-26, -4.395237e-26, 6.867589e-27, 1.840507e-25, -6.867535e-27, 
    6.592862e-26, -1.813036e-25, 5.494052e-26, -2.334968e-26, 3.159081e-26, 
    -9.065179e-26, 1.098813e-26, -1.648212e-26, 6.867565e-26, -1.208691e-25, 
    4.257891e-26, -9.477233e-26, -6.867559e-26, 2.747028e-26, -1.552069e-25, 
    1.922918e-25, -2.334968e-26, -6.592857e-26, -1.057604e-25, -1.236161e-25, 
    1.648217e-26, 2.472325e-26, -4.669939e-26, 1.208691e-25, -5.494023e-27, 
    7.691672e-26, -6.592857e-26, 3.296432e-26, -1.263631e-25, 7.004916e-26, 
    1.373515e-26, -9.751935e-26, 4.669945e-26, -1.098807e-26, 7.554321e-26, 
    -7.142262e-26, 1.675685e-25, -1.620744e-25, 3.571135e-26, 1.92292e-26, 
    8.378428e-26, 4.120564e-27, 1.510866e-26, -1.208691e-25, -1.579539e-25, 
    2.334974e-26, 9.339887e-26, -6.592857e-26, 1.181221e-25, 2.675717e-32, 
    1.236164e-26, -2.747022e-26, 2.197622e-26, -1.455923e-25, -1.922917e-25, 
    5.906106e-26, 6.043457e-26, 4.12054e-26, -3.021725e-26, 2.884379e-26, 
    3.433784e-26, -5.219344e-26, 3.845837e-26, 3.296432e-26, -8.241047e-27, 
    8.653131e-26, -5.219344e-26, -7.966369e-26, -1.236161e-25, 1.510866e-26, 
    1.442188e-25, 2.197622e-26, -3.159076e-26, 1.181221e-25, 6.180808e-26, 
    2.060271e-26, 3.845837e-26, 3.571135e-26, -5.906101e-26, -2.197617e-26, 
    -3.57113e-26, -1.37351e-26, 3.983189e-26, -1.74436e-25, -1.922915e-26, 
    9.889292e-26, -4.669939e-26, -3.845832e-26, -5.631398e-26, -1.291101e-25, 
    2.156415e-25, -1.071339e-25, -3.296427e-26, 3.571135e-26, 2.747028e-26, 
    -1.318572e-25, -3.845832e-26, -1.112545e-25, -1.648212e-26, 
    -6.318154e-26, 1.373539e-27, 2.884379e-26, 9.614589e-26, -8.241047e-27, 
    9.065185e-26, -3.845832e-26, 3.571135e-26, -5.494023e-27, -5.768749e-26, 
    1.12628e-25, -4.944642e-26, 2.675725e-32, -2.747022e-26, -7.691667e-26, 
    2.884379e-26, -5.494023e-27, 2.197622e-26, -5.768749e-26, 2.747052e-27, 
    2.472325e-26, 4.944647e-26, -1.483393e-25, -7.554316e-26, -1.304836e-25, 
    -1.09881e-25, 1.510864e-25, 1.098813e-26, 2.747052e-27, -1.854241e-25, 
    -4.257886e-26, -1.620744e-25, -4.395237e-26, -3.159076e-26, 
    -9.889287e-26, -1.346042e-25, 8.241101e-27, 9.889292e-26, -9.889287e-26, 
    -6.318154e-26, -7.554316e-26, -1.304836e-25, -5.906101e-26, 8.241101e-27, 
    8.790482e-26, -1.291101e-25, 7.829024e-26, 6.31816e-26, 6.867565e-26, 
    6.867589e-27, 7.279618e-26, -8.790477e-26, -1.098807e-26, -3.021725e-26, 
    3.571135e-26, 1.098813e-26, -1.071339e-25, -3.983183e-26, -1.071339e-25, 
    -5.081993e-26, -6.867559e-26, 2.884379e-26, 1.098813e-26, -2.47232e-26, 
    -8.241071e-26, 3.845837e-26, -1.37351e-26, 6.043457e-26, -5.494047e-26, 
    -1.565804e-25, -6.592857e-26, 6.31816e-26, -8.241047e-27, -4.120535e-26, 
    7.279618e-26, 5.21935e-26, 1.469658e-25, -8.241071e-26, 2.675723e-32, 
    -1.510863e-25, 5.768755e-26, -1.400982e-25, -1.428453e-25, 8.241101e-27, 
    5.494076e-27, 1.222426e-25, -7.691667e-26, 4.669945e-26, 5.081998e-26, 
    3.02173e-26, -7.142262e-26, 1.785569e-26, 3.983189e-26, 4.395242e-26, 
    -1.37351e-26, 3.571135e-26, -9.889287e-26, -6.730208e-26, -1.524598e-25, 
    6.592862e-26, -1.098807e-26, -7.416964e-26, -4.120511e-27, -2.197617e-26, 
    -8.10372e-26, 8.790482e-26, -7.966369e-26, -7.279613e-26, 1.016399e-25, 
    -3.845832e-26, -8.10372e-26, 1.016399e-25, 5.768755e-26, -1.950387e-25, 
    6.867589e-27, -4.120535e-26, -8.241047e-27, 3.433784e-26, -4.944642e-26, 
    -3.708481e-26, 1.373515e-26, 5.494076e-27, 8.241101e-27, -4.395237e-26, 
    2.747052e-27, -7.279613e-26, 5.768755e-26, 5.494076e-27, -2.197617e-26, 
    1.373515e-26, -2.197617e-26, 3.983189e-26, -9.889287e-26, -1.675685e-25, 
    -3.296427e-26, 2.115209e-25, 9.889292e-26, -2.747022e-26, 3.571135e-26 ;

 M_SOIL1C_TO_LEACHING =
  4.135503e-20, 1.727991e-20, 1.959381e-20, 4.637576e-20, 1.660758e-21, 
    -8.47881e-21, -3.013344e-20, -1.915246e-20, 9.781932e-21, -4.377807e-21, 
    1.725902e-20, 6.141336e-20, 1.93388e-22, -2.85202e-20, -4.45669e-21, 
    1.156538e-20, 2.05545e-22, -3.357004e-20, 1.763081e-20, -3.005537e-22, 
    -2.769356e-21, -1.972017e-20, -2.096135e-21, -1.514279e-20, 1.877417e-20, 
    1.597088e-20, 1.565283e-20, -9.934879e-21, -6.52657e-21, -1.524259e-20, 
    -7.22434e-21, 2.24231e-20, 2.422973e-20, 2.798865e-20, 4.160639e-20, 
    1.948583e-21, -1.846882e-20, 3.62441e-20, -3.204498e-20, 1.181391e-20, 
    -4.435773e-21, 5.607391e-21, -3.214377e-21, 5.801913e-21, -8.770005e-21, 
    -2.63409e-20, -3.039628e-21, 3.388815e-21, -7.001241e-21, -6.418548e-21, 
    2.220654e-20, 2.453536e-20, 3.742904e-20, -1.075706e-20, -6.917876e-21, 
    1.306952e-20, -3.138086e-20, 7.096824e-21, -1.348201e-20, -3.874513e-20, 
    3.507494e-23, 4.627033e-20, 1.958984e-20, -2.770932e-20, -4.481112e-20, 
    -6.200117e-20, 1.06321e-20, -4.168865e-21, 2.210094e-21, 3.415133e-20, 
    4.495343e-22, -5.618169e-21, 1.04325e-20, -1.849055e-22, 2.347516e-21, 
    -1.718947e-20, 2.441381e-21, 3.628822e-20, -2.327921e-20, -1.078336e-20, 
    -1.326121e-20, 9.075662e-21, 9.514435e-21, 1.833651e-20, -4.051814e-20, 
    -3.222859e-21, -1.003356e-20, 2.49341e-21, -8.100534e-21, -1.030807e-20, 
    -2.405106e-20, -8.054446e-21, 1.316168e-20, -3.001528e-20, 8.220948e-21, 
    -7.158956e-22, 1.191962e-20, 2.636747e-20, -4.126746e-21, 1.843207e-20, 
    -2.551559e-20, 1.995429e-20, 2.208946e-20, 1.332624e-20, 1.539183e-21, 
    1.724347e-20, -2.087684e-20, 1.859634e-20, -6.939601e-21, -3.058355e-20, 
    -2.486676e-20, 2.618213e-22, -1.215262e-20, -7.431591e-21, -5.038914e-20, 
    3.365654e-20, -3.17176e-20, -1.874789e-20, -6.983175e-21, 5.581959e-21, 
    3.053181e-20, -5.368504e-21, 6.774249e-22, -8.57296e-21, 2.128228e-20, 
    3.99671e-20, -2.453593e-20, 2.987058e-21, -2.054718e-20, -4.089729e-20, 
    -4.905652e-21, 1.506305e-20, 1.259875e-20, -2.216807e-20, -1.187327e-20, 
    4.28591e-21, 1.410771e-20, 9.758735e-21, 4.56383e-21, -3.741746e-20, 
    -1.001661e-20, 1.234515e-20, 2.658289e-20, -2.528036e-20, -1.295193e-21, 
    3.644938e-20, 3.097065e-20, 1.022328e-20, 1.597712e-20, 1.426094e-20, 
    -5.659153e-21, 1.554934e-20, -1.29567e-20, -1.618435e-20, -7.09963e-21, 
    -1.108871e-20, -1.968824e-20, 3.490564e-20, 7.162144e-21, -1.157754e-20, 
    2.037557e-20, 2.278016e-20, -1.882534e-20, 2.09396e-20, -1.337655e-20, 
    -2.232584e-20, -6.041389e-21, -4.227502e-20, -2.255033e-20, 
    -4.366222e-21, -1.273333e-20, 2.851048e-21, -1.000925e-20, 1.869303e-20, 
    -3.520366e-20, 4.061257e-20, -9.237388e-21, 2.068597e-20, 5.296675e-21, 
    -9.388085e-21, 8.680126e-21, -1.165785e-20, 1.759519e-20, -1.574273e-20, 
    8.949564e-21, 5.361744e-21, -1.594205e-20, -2.447542e-20, 1.197647e-20, 
    -1.439354e-20, -1.356683e-20, -2.460776e-20, 4.288734e-21, 1.679565e-22, 
    -1.95678e-20, -9.474344e-22, -1.675492e-20, -1.152554e-20, 2.519414e-20, 
    -4.677497e-20, 2.046772e-20, -3.995042e-20, 1.175058e-20, -2.537905e-20, 
    -1.020205e-20, -1.831645e-20, 3.338684e-20, 4.145738e-20, 1.665623e-20, 
    1.844268e-21, -7.693102e-21, 3.17451e-21, -2.927124e-21, -2.617577e-20, 
    4.004878e-21, 2.471915e-21, -3.244987e-20, 2.841558e-20, 3.350916e-21, 
    -5.019611e-21, 3.527209e-20, 3.794387e-20, 1.651142e-21, -2.600077e-20, 
    -2.568751e-20, 2.487468e-21, -5.248064e-21, 2.700248e-20, 7.000696e-21, 
    2.743703e-20, 1.76878e-21, -6.844956e-22, 3.930043e-20, -2.457949e-20, 
    3.019282e-21, 3.485818e-20, -2.506378e-20, 3.776804e-20, -2.880406e-20, 
    -5.414861e-20, -3.391639e-21, 8.349299e-21, -4.797368e-21, -3.451153e-20, 
    2.902288e-20, -2.085621e-20, 9.332943e-21, 3.725062e-20, -2.189297e-20, 
    -2.553344e-21, -2.421674e-20, -8.226623e-21, -3.973199e-21, 1.47625e-20, 
    -1.866363e-20, 1.243816e-20, -3.195819e-20, -2.323931e-20, 2.492554e-21, 
    -1.398937e-21, -4.288751e-21, -1.764014e-20, 3.69559e-21, -2.383111e-20, 
    2.678253e-20, -8.852385e-22, 1.590811e-20, -1.493891e-20, -2.020478e-20, 
    -5.56128e-22, -3.663711e-20, 1.392251e-20, 8.297008e-21, -1.740518e-20, 
    1.374078e-21, 3.830634e-20, 1.533758e-20, -3.331672e-20, 1.267002e-20, 
    -2.18418e-20, -1.309495e-20, 2.507736e-20, -1.094163e-21, 2.642346e-20, 
    5.452475e-21, -2.014371e-20, -3.878216e-21, -2.368607e-20, -2.431502e-21, 
    1.123034e-21, 2.57189e-20, 1.570882e-20, 1.750837e-20, -1.635003e-20, 
    3.787176e-21, 6.093134e-21, -3.332377e-20, 5.660976e-20, -1.797608e-21, 
    -3.36899e-20, 1.249104e-20, 1.297168e-20, 1.16943e-20, 1.259793e-20, 
    8.178829e-21, -1.098466e-20, -2.081351e-20, -3.227909e-20, -2.69909e-20, 
    2.289809e-20, 2.918714e-20, -3.51474e-20, 1.460107e-20, -2.673785e-21, 
    1.929043e-20, 2.463716e-20, -7.778761e-21, -7.283046e-22, -6.003873e-20, 
    2.720123e-20, 1.95029e-21, 9.033153e-22, -1.197987e-20, 4.77555e-22, 
    8.511345e-21, 4.175113e-20, -1.660053e-20, -2.703131e-20, 4.892378e-21, 
    2.530453e-21, 3.857805e-20, 4.773905e-21, 4.346447e-20, -1.064395e-20, 
    3.603319e-20, 1.172315e-20, 1.366127e-20, -1.192108e-20 ;

 M_SOIL2C_TO_LEACHING =
  -1.759351e-20, 4.237282e-21, 4.365054e-20, -1.951435e-20, -5.106027e-22, 
    -1.299707e-21, -2.739394e-21, 1.639978e-20, -1.203244e-20, -6.194053e-21, 
    -4.314476e-21, 4.927977e-22, 1.922653e-20, -1.123373e-20, -1.011102e-20, 
    -3.139244e-20, -4.644023e-20, 4.461793e-21, -3.47674e-20, -9.649595e-21, 
    -2.309967e-20, 1.652848e-21, 2.338183e-21, -2.04302e-21, -2.309033e-20, 
    8.154515e-21, -1.582672e-20, 5.47282e-21, -1.82217e-20, 9.403066e-21, 
    3.626163e-20, -3.574763e-20, -9.38526e-21, 5.038561e-21, -1.602716e-20, 
    2.309033e-20, -7.70155e-22, 3.861197e-20, -2.308215e-20, 1.602122e-20, 
    -6.330937e-20, -2.718486e-20, -2.312654e-20, 4.689373e-21, -1.587336e-20, 
    1.260612e-20, 2.074849e-20, -1.928452e-20, -1.013081e-20, -2.492384e-20, 
    2.06498e-20, -2.096336e-20, -8.467769e-22, 1.136804e-20, -3.165593e-20, 
    -9.598994e-21, 1.010734e-20, 4.236181e-21, 1.332624e-20, 3.164321e-21, 
    7.761519e-21, -3.140685e-20, 1.103355e-20, -1.321456e-20, -1.508991e-20, 
    -5.506733e-21, 3.105531e-21, 7.807607e-21, -3.812738e-20, -2.803728e-20, 
    -4.251717e-21, 6.582846e-21, 1.984884e-20, -3.689495e-20, 1.01116e-20, 
    -4.539893e-20, 1.539272e-20, -1.424107e-21, -3.680362e-20, 3.838628e-21, 
    1.887766e-20, 1.00734e-20, 2.051664e-20, -9.839586e-21, 2.777717e-20, 
    -7.686603e-21, 8.973788e-22, 5.762123e-22, -8.21983e-21, -3.143907e-22, 
    -1.807161e-20, -2.050052e-20, -1.775262e-21, -3.672671e-21, 
    -2.258566e-20, -1.457308e-20, -7.608854e-21, 3.76683e-21, 1.388236e-20, 
    -3.768716e-20, -2.834603e-20, -6.511374e-20, 6.741993e-21, 1.669667e-20, 
    1.278523e-21, 6.044776e-22, -3.264155e-20, 1.519762e-20, 1.226372e-20, 
    2.199475e-20, -1.361348e-21, 4.085574e-20, 1.142292e-20, 1.237992e-20, 
    6.328079e-21, 1.984544e-20, -3.343122e-20, 1.251451e-20, -1.656237e-20, 
    -3.630207e-20, 8.775108e-21, 1.657362e-21, -7.49435e-21, 1.819966e-20, 
    2.750604e-20, 3.942427e-20, 3.52602e-20, 2.431485e-21, 3.094035e-20, 
    1.495646e-20, 2.722151e-21, -3.688225e-21, -1.919996e-20, 4.884571e-20, 
    -3.163532e-20, 8.900652e-21, 2.479153e-20, -6.962519e-21, -4.901732e-20, 
    -3.02881e-20, -3.538659e-20, 4.459808e-21, -3.349568e-20, 3.373799e-20, 
    -3.474181e-21, -3.940248e-20, -2.38294e-20, 3.322228e-20, 1.035755e-20, 
    1.955422e-20, 1.21631e-21, -7.756154e-21, 9.205147e-21, -4.218147e-20, 
    7.807345e-21, -1.012853e-20, 1.885531e-20, -1.064481e-20, -1.332624e-20, 
    -1.62395e-20, 1.328834e-20, 7.653807e-21, -1.430647e-20, 2.242027e-20, 
    -1.840124e-20, -4.05733e-20, -1.724232e-20, -2.814558e-20, 3.853357e-21, 
    4.405483e-20, 4.283768e-20, 2.550232e-20, -2.728061e-21, 2.923013e-20, 
    8.862752e-21, 1.674616e-20, 2.921449e-21, 5.951448e-22, -1.114976e-20, 
    -3.204613e-20, 2.586419e-21, 1.912193e-20, 3.301743e-21, 6.343632e-21, 
    -8.941947e-21, -1.469803e-20, -2.86556e-20, 9.07509e-21, -1.05375e-21, 
    6.242141e-21, -2.853827e-20, 1.075592e-20, 3.06706e-21, 1.516822e-20, 
    -1.069147e-20, 3.299464e-21, -3.360593e-20, 3.673606e-20, 2.848427e-20, 
    -8.533942e-21, -2.109908e-20, -3.651754e-21, -8.137272e-21, 
    -1.072426e-20, -2.296085e-20, -3.022591e-20, 1.220039e-20, 4.52143e-20, 
    -7.291066e-21, -7.656145e-22, 2.640903e-20, -1.143959e-20, -2.342028e-20, 
    -7.434416e-21, -1.49149e-20, 3.207806e-20, -2.61464e-20, 1.703735e-20, 
    9.48449e-21, 1.404975e-20, -7.822309e-21, -4.863155e-22, 4.941845e-21, 
    3.70971e-20, 4.10689e-20, 4.293351e-20, 4.803616e-21, 4.32793e-20, 
    -1.001744e-20, 1.015258e-20, -6.804751e-21, -1.19759e-20, 1.762601e-20, 
    5.958285e-21, 1.719909e-20, 3.166583e-21, -4.819882e-20, -2.588683e-20, 
    4.556009e-20, -2.825951e-20, 2.331993e-20, -2.306773e-20, -2.275134e-20, 
    2.067327e-20, -2.269734e-20, 1.157772e-21, 1.828985e-20, -4.24547e-21, 
    5.472541e-21, 6.078153e-21, 7.661162e-21, -6.462095e-21, 3.376428e-20, 
    -3.414557e-21, -6.62721e-21, 1.237457e-20, 3.263393e-20, 3.366559e-20, 
    1.006976e-20, -1.766221e-20, -1.802126e-20, 1.737492e-20, 1.725108e-20, 
    6.992792e-21, -3.265936e-20, -1.830201e-20, -8.906872e-21, 5.130719e-21, 
    -2.276248e-21, -8.262243e-21, -4.324093e-21, 3.049254e-21, -3.445353e-21, 
    -3.98065e-20, -2.436689e-20, -2.368379e-20, 3.313578e-20, 4.10409e-20, 
    3.339023e-20, -8.288247e-21, 2.039451e-20, -1.013448e-20, 1.603083e-20, 
    3.50029e-20, -1.045313e-20, -5.432587e-20, 2.708194e-20, -2.922502e-20, 
    -2.182371e-20, 2.897338e-20, -3.493702e-21, 2.422947e-20, -1.266409e-20, 
    2.226533e-20, 9.97304e-21, -2.223508e-20, -1.176556e-20, -6.164947e-21, 
    -1.394512e-20, 9.130232e-21, -9.581751e-21, -8.354973e-21, 1.892997e-20, 
    5.546339e-21, -2.660638e-20, 1.285999e-20, -8.216728e-21, -5.322209e-20, 
    1.570862e-21, 3.28619e-21, 1.939814e-20, -3.488361e-20, 2.298093e-20, 
    1.313624e-20, -1.694291e-20, 1.112773e-20, 3.864732e-20, -5.9363e-20, 
    2.864061e-20, 3.894194e-20, 4.581662e-21, 8.503981e-21, -5.507635e-22, 
    -9.12797e-21, -1.424622e-20, -2.454272e-20, -1.356092e-20, 2.981143e-20, 
    -1.984884e-20, 7.783865e-21, 4.340882e-20, -1.6406e-20, 2.60918e-20, 
    -7.2198e-21, 1.096656e-20, -2.172305e-20, 9.002029e-22, -2.785405e-20 ;

 M_SOIL3C_TO_LEACHING =
  2.261537e-20, 1.98576e-20, -6.485968e-22, -2.363235e-20, -1.402204e-20, 
    -3.729048e-20, -1.287751e-20, -2.541267e-20, 1.623863e-20, -6.661991e-21, 
    -2.533849e-21, -4.598332e-21, -3.922579e-20, -2.368405e-20, 2.246748e-20, 
    2.128736e-20, -1.720728e-20, -8.719421e-21, -1.380545e-20, 2.026071e-21, 
    -1.064029e-20, 2.664596e-20, -1.364459e-20, -2.069677e-20, -1.820477e-20, 
    -3.503544e-20, -2.225797e-20, -1.758019e-21, -5.260482e-21, 2.96268e-20, 
    6.659158e-21, 4.085189e-21, 2.301373e-20, 1.909932e-20, 1.435536e-20, 
    -3.710983e-20, -1.276274e-20, 1.430478e-20, 3.30207e-20, -4.050686e-21, 
    8.895287e-21, -3.265539e-20, 8.396841e-21, 3.636822e-20, -1.349305e-20, 
    -3.776944e-20, 1.987524e-22, -5.634529e-21, 7.912232e-21, 4.176189e-20, 
    1.796555e-20, 8.960014e-21, 1.377805e-20, 3.048389e-21, -9.958076e-21, 
    -6.180779e-21, 1.378455e-20, -3.914919e-20, -3.190702e-20, -4.960222e-21, 
    2.235834e-20, 1.430043e-21, -2.860105e-20, -8.669374e-21, 4.575941e-20, 
    3.370689e-20, 2.359642e-20, -2.366963e-20, 3.918787e-22, -2.456678e-20, 
    5.937335e-21, -2.814048e-20, 1.025464e-20, -1.529319e-20, 2.940399e-21, 
    2.615288e-20, 1.776032e-20, -3.365148e-20, 1.095441e-20, 3.261894e-20, 
    -8.600669e-21, 7.122539e-21, 2.848258e-20, -1.621997e-20, 2.245957e-20, 
    -1.488581e-21, 3.763255e-22, -5.797383e-21, 8.794058e-21, 1.579475e-20, 
    -3.575045e-20, 3.07328e-21, -3.6105e-20, -3.409109e-20, -1.836391e-20, 
    1.112205e-20, 1.96071e-20, -8.152825e-21, 1.312663e-20, 4.108051e-20, 
    1.787419e-21, -1.549221e-20, 3.030252e-20, 1.153145e-20, 1.282665e-20, 
    -1.566639e-20, 1.742444e-20, -8.523754e-21, -3.949457e-21, 2.948335e-21, 
    -4.521998e-20, 2.288733e-20, 1.120376e-20, -2.058759e-20, -1.371357e-20, 
    2.934178e-21, -2.549016e-20, -2.709326e-20, -4.510149e-20, 4.179298e-20, 
    5.145714e-22, -1.719284e-20, 2.267499e-20, -5.401274e-21, 2.030291e-21, 
    -3.589098e-20, 1.908603e-20, -7.467211e-21, -1.789403e-20, -2.23075e-21, 
    1.318402e-20, 2.052048e-21, 3.597862e-20, -1.717731e-20, -1.372687e-20, 
    -4.044775e-20, 1.278226e-20, 1.388493e-20, -2.409319e-20, 1.450747e-20, 
    -8.905754e-21, -7.575469e-21, -2.581249e-20, 3.879923e-21, 2.315027e-20, 
    -4.4646e-21, 4.125269e-20, 2.579976e-20, -4.76401e-21, 5.682852e-22, 
    1.210635e-21, 4.319223e-20, -4.522109e-20, 1.136607e-20, 8.995634e-21, 
    -2.716873e-20, -2.835773e-21, 3.851078e-21, 4.062276e-20, 1.540176e-20, 
    -1.404578e-20, -2.642695e-21, 3.118211e-20, -3.111709e-20, -1.784229e-20, 
    1.417923e-20, 1.375767e-21, 1.892429e-20, -1.369577e-20, 1.251705e-20, 
    -1.035359e-20, 1.566273e-20, 1.894213e-20, -2.819674e-21, 3.010995e-22, 
    -1.034542e-20, -3.426951e-20, -1.742809e-20, -3.475864e-20, 
    -1.686066e-20, 1.38509e-21, -2.711107e-20, 1.314304e-20, -2.647124e-20, 
    -7.891593e-21, -1.646911e-21, -2.486448e-20, -1.541732e-20, 
    -1.026318e-21, 1.741508e-20, -3.448328e-20, 9.164987e-21, 3.247106e-20, 
    1.354337e-20, -6.964225e-21, 4.66738e-20, -2.889256e-20, 2.057263e-20, 
    -3.677757e-21, 4.823944e-21, 6.900895e-21, 3.741349e-20, -9.560261e-21, 
    1.87869e-20, 4.990447e-22, -2.969182e-20, -9.043983e-21, -4.150234e-20, 
    1.629349e-20, 3.618647e-21, -8.170918e-21, -1.758019e-21, -4.63507e-21, 
    7.807607e-21, 3.944371e-21, 1.009076e-21, 8.060928e-21, 1.122297e-20, 
    -3.287585e-21, -1.961048e-20, -1.396804e-20, -3.403683e-20, 4.538477e-20, 
    3.821106e-21, -1.937216e-20, 3.033782e-22, -5.238747e-20, -5.779383e-20, 
    -7.009152e-21, -9.388085e-21, 5.452448e-21, -3.9301e-20, -1.986662e-20, 
    1.396067e-20, -2.905878e-20, -2.112571e-21, 4.894346e-21, 3.64102e-21, 
    -2.13405e-20, 3.855628e-20, -4.611188e-22, 1.930034e-20, -2.074339e-20, 
    -2.369058e-20, 3.539201e-21, -2.311323e-21, 4.424059e-20, 6.966766e-21, 
    6.325817e-21, -2.033005e-20, 2.570138e-20, 1.525644e-20, -1.54405e-20, 
    -9.078797e-21, 2.170638e-20, -1.125496e-20, -1.353121e-20, -1.550045e-20, 
    -7.598665e-21, -1.218855e-20, 2.060825e-21, 2.059609e-20, 1.000189e-20, 
    2.348167e-20, 4.20237e-20, -1.132988e-20, 2.261309e-20, 2.185961e-20, 
    -2.38673e-20, -2.084122e-20, -1.928792e-20, 1.14127e-20, -1.467628e-20, 
    1.25411e-20, -7.275513e-21, 2.824311e-20, 5.458116e-20, -6.659713e-21, 
    2.937234e-20, -2.938692e-21, -1.320297e-20, -8.712039e-21, 2.173918e-20, 
    2.087345e-20, -2.447542e-20, -1.85951e-21, -2.823831e-20, -2.527896e-20, 
    -5.159044e-20, -2.249801e-20, -1.320637e-20, 1.384589e-20, -3.81678e-20, 
    -4.479581e-21, 2.108606e-20, 2.274625e-20, 2.987898e-20, -2.542004e-20, 
    -1.253429e-20, -3.321945e-20, -3.016908e-20, -2.147312e-20, 8.738304e-23, 
    1.108589e-20, 8.134448e-21, 2.761118e-20, -2.979474e-20, -7.901193e-21, 
    1.410771e-20, 1.429628e-20, -2.820378e-20, 2.74441e-20, 3.791308e-20, 
    1.217948e-20, -5.720777e-21, -1.556404e-20, 1.364742e-20, 3.478149e-21, 
    1.701755e-20, 1.264541e-20, 1.354219e-22, 5.210534e-22, -1.457477e-20, 
    -2.003007e-20, -1.235788e-20, 1.029715e-21, -2.07072e-20, -6.713989e-21, 
    -3.297772e-20, 4.589572e-21, -3.983226e-20, 1.656322e-20, -4.505864e-21, 
    6.174955e-20, -2.694284e-20, 1.416424e-22, 2.019009e-20, 3.498963e-20 ;

 NBP =
  -6.215762e-08, -6.243169e-08, -6.237841e-08, -6.259947e-08, -6.247685e-08, 
    -6.26216e-08, -6.221319e-08, -6.244257e-08, -6.229614e-08, -6.21823e-08, 
    -6.302847e-08, -6.260934e-08, -6.346394e-08, -6.319659e-08, 
    -6.386823e-08, -6.342233e-08, -6.395815e-08, -6.385538e-08, 
    -6.416472e-08, -6.40761e-08, -6.447177e-08, -6.420563e-08, -6.46769e-08, 
    -6.440823e-08, -6.445025e-08, -6.419685e-08, -6.269369e-08, 
    -6.297628e-08, -6.267695e-08, -6.271725e-08, -6.269916e-08, 
    -6.247938e-08, -6.236861e-08, -6.213668e-08, -6.217878e-08, 
    -6.234914e-08, -6.273537e-08, -6.260426e-08, -6.29347e-08, -6.292724e-08, 
    -6.329513e-08, -6.312926e-08, -6.374764e-08, -6.357188e-08, -6.40798e-08, 
    -6.395206e-08, -6.40738e-08, -6.403688e-08, -6.407428e-08, -6.388693e-08, 
    -6.39672e-08, -6.380235e-08, -6.316031e-08, -6.334899e-08, -6.278628e-08, 
    -6.244793e-08, -6.222324e-08, -6.20638e-08, -6.208634e-08, -6.212931e-08, 
    -6.235014e-08, -6.255778e-08, -6.271602e-08, -6.282187e-08, 
    -6.292617e-08, -6.324185e-08, -6.340898e-08, -6.378317e-08, 
    -6.371565e-08, -6.383004e-08, -6.393935e-08, -6.412285e-08, 
    -6.409265e-08, -6.417349e-08, -6.382704e-08, -6.405729e-08, 
    -6.367719e-08, -6.378114e-08, -6.295448e-08, -6.263964e-08, 
    -6.250578e-08, -6.238865e-08, -6.210367e-08, -6.230047e-08, 
    -6.222289e-08, -6.240747e-08, -6.252476e-08, -6.246675e-08, 
    -6.282476e-08, -6.268557e-08, -6.341888e-08, -6.310301e-08, -6.39266e-08, 
    -6.372951e-08, -6.397384e-08, -6.384917e-08, -6.406279e-08, 
    -6.387053e-08, -6.420358e-08, -6.427612e-08, -6.422655e-08, 
    -6.441695e-08, -6.385987e-08, -6.40738e-08, -6.246512e-08, -6.247458e-08, 
    -6.251866e-08, -6.232491e-08, -6.231306e-08, -6.213552e-08, 
    -6.229349e-08, -6.236077e-08, -6.253156e-08, -6.263257e-08, -6.27286e-08, 
    -6.293975e-08, -6.317556e-08, -6.350534e-08, -6.374228e-08, 
    -6.390112e-08, -6.380372e-08, -6.388971e-08, -6.379359e-08, 
    -6.374854e-08, -6.424895e-08, -6.396795e-08, -6.438957e-08, 
    -6.436624e-08, -6.417542e-08, -6.436887e-08, -6.248122e-08, 
    -6.242679e-08, -6.223777e-08, -6.238569e-08, -6.211619e-08, 
    -6.226703e-08, -6.235377e-08, -6.268847e-08, -6.276202e-08, 
    -6.283021e-08, -6.296489e-08, -6.313774e-08, -6.344097e-08, 
    -6.370482e-08, -6.394571e-08, -6.392806e-08, -6.393427e-08, 
    -6.398808e-08, -6.385479e-08, -6.400997e-08, -6.403601e-08, 
    -6.396792e-08, -6.436311e-08, -6.425022e-08, -6.436574e-08, 
    -6.429224e-08, -6.244449e-08, -6.253608e-08, -6.248658e-08, 
    -6.257967e-08, -6.251409e-08, -6.280568e-08, -6.289311e-08, 
    -6.330224e-08, -6.313434e-08, -6.340156e-08, -6.316149e-08, 
    -6.320403e-08, -6.341026e-08, -6.317446e-08, -6.369027e-08, 
    -6.334054e-08, -6.399017e-08, -6.36409e-08, -6.401206e-08, -6.394467e-08, 
    -6.405626e-08, -6.415619e-08, -6.428195e-08, -6.451393e-08, 
    -6.446022e-08, -6.465423e-08, -6.267265e-08, -6.279146e-08, 
    -6.278102e-08, -6.290536e-08, -6.299733e-08, -6.319667e-08, -6.35164e-08, 
    -6.339616e-08, -6.361689e-08, -6.366121e-08, -6.332587e-08, 
    -6.353175e-08, -6.2871e-08, -6.297773e-08, -6.291419e-08, -6.268202e-08, 
    -6.342385e-08, -6.304312e-08, -6.37462e-08, -6.353994e-08, -6.414194e-08, 
    -6.384253e-08, -6.443064e-08, -6.468203e-08, -6.491868e-08, -6.51952e-08, 
    -6.285632e-08, -6.277559e-08, -6.292016e-08, -6.312016e-08, 
    -6.330577e-08, -6.355251e-08, -6.357777e-08, -6.362399e-08, 
    -6.374373e-08, -6.384442e-08, -6.363859e-08, -6.386966e-08, 
    -6.300247e-08, -6.345691e-08, -6.274506e-08, -6.295939e-08, 
    -6.310837e-08, -6.304303e-08, -6.338242e-08, -6.346242e-08, 
    -6.378748e-08, -6.361945e-08, -6.461998e-08, -6.417729e-08, 
    -6.540579e-08, -6.506244e-08, -6.274738e-08, -6.285605e-08, 
    -6.323427e-08, -6.305431e-08, -6.356899e-08, -6.369568e-08, 
    -6.379868e-08, -6.393034e-08, -6.394456e-08, -6.402257e-08, 
    -6.389474e-08, -6.401752e-08, -6.355304e-08, -6.37606e-08, -6.319105e-08, 
    -6.332966e-08, -6.326589e-08, -6.319594e-08, -6.341183e-08, 
    -6.364183e-08, -6.364677e-08, -6.372051e-08, -6.392831e-08, 
    -6.357108e-08, -6.467708e-08, -6.399399e-08, -6.297455e-08, 
    -6.318386e-08, -6.321378e-08, -6.313269e-08, -6.368298e-08, 
    -6.348358e-08, -6.402067e-08, -6.387551e-08, -6.411335e-08, 
    -6.399516e-08, -6.397777e-08, -6.382598e-08, -6.373148e-08, 
    -6.349272e-08, -6.329847e-08, -6.314445e-08, -6.318027e-08, 
    -6.334945e-08, -6.365591e-08, -6.394584e-08, -6.388233e-08, 
    -6.409527e-08, -6.353167e-08, -6.376798e-08, -6.367664e-08, 
    -6.391483e-08, -6.339297e-08, -6.383731e-08, -6.327939e-08, 
    -6.332831e-08, -6.347963e-08, -6.378401e-08, -6.385137e-08, 
    -6.392327e-08, -6.387891e-08, -6.366369e-08, -6.362843e-08, 
    -6.347595e-08, -6.343384e-08, -6.331766e-08, -6.322146e-08, 
    -6.330935e-08, -6.340164e-08, -6.366378e-08, -6.390003e-08, 
    -6.415761e-08, -6.422066e-08, -6.452161e-08, -6.427662e-08, 
    -6.468089e-08, -6.433715e-08, -6.493221e-08, -6.386308e-08, 
    -6.432707e-08, -6.348652e-08, -6.357706e-08, -6.374083e-08, -6.41165e-08, 
    -6.39137e-08, -6.415087e-08, -6.362706e-08, -6.335529e-08, -6.328499e-08, 
    -6.315381e-08, -6.328799e-08, -6.327708e-08, -6.340547e-08, 
    -6.336422e-08, -6.367249e-08, -6.35069e-08, -6.397733e-08, -6.414901e-08, 
    -6.463389e-08, -6.493114e-08, -6.523376e-08, -6.536735e-08, 
    -6.540802e-08, -6.542501e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.215762e-08, 6.243169e-08, 6.237841e-08, 6.259947e-08, 6.247685e-08, 
    6.26216e-08, 6.221319e-08, 6.244257e-08, 6.229614e-08, 6.21823e-08, 
    6.302847e-08, 6.260934e-08, 6.346394e-08, 6.319659e-08, 6.386823e-08, 
    6.342233e-08, 6.395815e-08, 6.385538e-08, 6.416472e-08, 6.40761e-08, 
    6.447177e-08, 6.420563e-08, 6.46769e-08, 6.440823e-08, 6.445025e-08, 
    6.419685e-08, 6.269369e-08, 6.297628e-08, 6.267695e-08, 6.271725e-08, 
    6.269916e-08, 6.247938e-08, 6.236861e-08, 6.213668e-08, 6.217878e-08, 
    6.234914e-08, 6.273537e-08, 6.260426e-08, 6.29347e-08, 6.292724e-08, 
    6.329513e-08, 6.312926e-08, 6.374764e-08, 6.357188e-08, 6.40798e-08, 
    6.395206e-08, 6.40738e-08, 6.403688e-08, 6.407428e-08, 6.388693e-08, 
    6.39672e-08, 6.380235e-08, 6.316031e-08, 6.334899e-08, 6.278628e-08, 
    6.244793e-08, 6.222324e-08, 6.20638e-08, 6.208634e-08, 6.212931e-08, 
    6.235014e-08, 6.255778e-08, 6.271602e-08, 6.282187e-08, 6.292617e-08, 
    6.324185e-08, 6.340898e-08, 6.378317e-08, 6.371565e-08, 6.383004e-08, 
    6.393935e-08, 6.412285e-08, 6.409265e-08, 6.417349e-08, 6.382704e-08, 
    6.405729e-08, 6.367719e-08, 6.378114e-08, 6.295448e-08, 6.263964e-08, 
    6.250578e-08, 6.238865e-08, 6.210367e-08, 6.230047e-08, 6.222289e-08, 
    6.240747e-08, 6.252476e-08, 6.246675e-08, 6.282476e-08, 6.268557e-08, 
    6.341888e-08, 6.310301e-08, 6.39266e-08, 6.372951e-08, 6.397384e-08, 
    6.384917e-08, 6.406279e-08, 6.387053e-08, 6.420358e-08, 6.427612e-08, 
    6.422655e-08, 6.441695e-08, 6.385987e-08, 6.40738e-08, 6.246512e-08, 
    6.247458e-08, 6.251866e-08, 6.232491e-08, 6.231306e-08, 6.213552e-08, 
    6.229349e-08, 6.236077e-08, 6.253156e-08, 6.263257e-08, 6.27286e-08, 
    6.293975e-08, 6.317556e-08, 6.350534e-08, 6.374228e-08, 6.390112e-08, 
    6.380372e-08, 6.388971e-08, 6.379359e-08, 6.374854e-08, 6.424895e-08, 
    6.396795e-08, 6.438957e-08, 6.436624e-08, 6.417542e-08, 6.436887e-08, 
    6.248122e-08, 6.242679e-08, 6.223777e-08, 6.238569e-08, 6.211619e-08, 
    6.226703e-08, 6.235377e-08, 6.268847e-08, 6.276202e-08, 6.283021e-08, 
    6.296489e-08, 6.313774e-08, 6.344097e-08, 6.370482e-08, 6.394571e-08, 
    6.392806e-08, 6.393427e-08, 6.398808e-08, 6.385479e-08, 6.400997e-08, 
    6.403601e-08, 6.396792e-08, 6.436311e-08, 6.425022e-08, 6.436574e-08, 
    6.429224e-08, 6.244449e-08, 6.253608e-08, 6.248658e-08, 6.257967e-08, 
    6.251409e-08, 6.280568e-08, 6.289311e-08, 6.330224e-08, 6.313434e-08, 
    6.340156e-08, 6.316149e-08, 6.320403e-08, 6.341026e-08, 6.317446e-08, 
    6.369027e-08, 6.334054e-08, 6.399017e-08, 6.36409e-08, 6.401206e-08, 
    6.394467e-08, 6.405626e-08, 6.415619e-08, 6.428195e-08, 6.451393e-08, 
    6.446022e-08, 6.465423e-08, 6.267265e-08, 6.279146e-08, 6.278102e-08, 
    6.290536e-08, 6.299733e-08, 6.319667e-08, 6.35164e-08, 6.339616e-08, 
    6.361689e-08, 6.366121e-08, 6.332587e-08, 6.353175e-08, 6.2871e-08, 
    6.297773e-08, 6.291419e-08, 6.268202e-08, 6.342385e-08, 6.304312e-08, 
    6.37462e-08, 6.353994e-08, 6.414194e-08, 6.384253e-08, 6.443064e-08, 
    6.468203e-08, 6.491868e-08, 6.51952e-08, 6.285632e-08, 6.277559e-08, 
    6.292016e-08, 6.312016e-08, 6.330577e-08, 6.355251e-08, 6.357777e-08, 
    6.362399e-08, 6.374373e-08, 6.384442e-08, 6.363859e-08, 6.386966e-08, 
    6.300247e-08, 6.345691e-08, 6.274506e-08, 6.295939e-08, 6.310837e-08, 
    6.304303e-08, 6.338242e-08, 6.346242e-08, 6.378748e-08, 6.361945e-08, 
    6.461998e-08, 6.417729e-08, 6.540579e-08, 6.506244e-08, 6.274738e-08, 
    6.285605e-08, 6.323427e-08, 6.305431e-08, 6.356899e-08, 6.369568e-08, 
    6.379868e-08, 6.393034e-08, 6.394456e-08, 6.402257e-08, 6.389474e-08, 
    6.401752e-08, 6.355304e-08, 6.37606e-08, 6.319105e-08, 6.332966e-08, 
    6.326589e-08, 6.319594e-08, 6.341183e-08, 6.364183e-08, 6.364677e-08, 
    6.372051e-08, 6.392831e-08, 6.357108e-08, 6.467708e-08, 6.399399e-08, 
    6.297455e-08, 6.318386e-08, 6.321378e-08, 6.313269e-08, 6.368298e-08, 
    6.348358e-08, 6.402067e-08, 6.387551e-08, 6.411335e-08, 6.399516e-08, 
    6.397777e-08, 6.382598e-08, 6.373148e-08, 6.349272e-08, 6.329847e-08, 
    6.314445e-08, 6.318027e-08, 6.334945e-08, 6.365591e-08, 6.394584e-08, 
    6.388233e-08, 6.409527e-08, 6.353167e-08, 6.376798e-08, 6.367664e-08, 
    6.391483e-08, 6.339297e-08, 6.383731e-08, 6.327939e-08, 6.332831e-08, 
    6.347963e-08, 6.378401e-08, 6.385137e-08, 6.392327e-08, 6.387891e-08, 
    6.366369e-08, 6.362843e-08, 6.347595e-08, 6.343384e-08, 6.331766e-08, 
    6.322146e-08, 6.330935e-08, 6.340164e-08, 6.366378e-08, 6.390003e-08, 
    6.415761e-08, 6.422066e-08, 6.452161e-08, 6.427662e-08, 6.468089e-08, 
    6.433715e-08, 6.493221e-08, 6.386308e-08, 6.432707e-08, 6.348652e-08, 
    6.357706e-08, 6.374083e-08, 6.41165e-08, 6.39137e-08, 6.415087e-08, 
    6.362706e-08, 6.335529e-08, 6.328499e-08, 6.315381e-08, 6.328799e-08, 
    6.327708e-08, 6.340547e-08, 6.336422e-08, 6.367249e-08, 6.35069e-08, 
    6.397733e-08, 6.414901e-08, 6.463389e-08, 6.493114e-08, 6.523376e-08, 
    6.536735e-08, 6.540802e-08, 6.542501e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.215762e-08, -6.243169e-08, -6.237841e-08, -6.259947e-08, -6.247685e-08, 
    -6.26216e-08, -6.221319e-08, -6.244257e-08, -6.229614e-08, -6.21823e-08, 
    -6.302847e-08, -6.260934e-08, -6.346394e-08, -6.319659e-08, 
    -6.386823e-08, -6.342233e-08, -6.395815e-08, -6.385538e-08, 
    -6.416472e-08, -6.40761e-08, -6.447177e-08, -6.420563e-08, -6.46769e-08, 
    -6.440823e-08, -6.445025e-08, -6.419685e-08, -6.269369e-08, 
    -6.297628e-08, -6.267695e-08, -6.271725e-08, -6.269916e-08, 
    -6.247938e-08, -6.236861e-08, -6.213668e-08, -6.217878e-08, 
    -6.234914e-08, -6.273537e-08, -6.260426e-08, -6.29347e-08, -6.292724e-08, 
    -6.329513e-08, -6.312926e-08, -6.374764e-08, -6.357188e-08, -6.40798e-08, 
    -6.395206e-08, -6.40738e-08, -6.403688e-08, -6.407428e-08, -6.388693e-08, 
    -6.39672e-08, -6.380235e-08, -6.316031e-08, -6.334899e-08, -6.278628e-08, 
    -6.244793e-08, -6.222324e-08, -6.20638e-08, -6.208634e-08, -6.212931e-08, 
    -6.235014e-08, -6.255778e-08, -6.271602e-08, -6.282187e-08, 
    -6.292617e-08, -6.324185e-08, -6.340898e-08, -6.378317e-08, 
    -6.371565e-08, -6.383004e-08, -6.393935e-08, -6.412285e-08, 
    -6.409265e-08, -6.417349e-08, -6.382704e-08, -6.405729e-08, 
    -6.367719e-08, -6.378114e-08, -6.295448e-08, -6.263964e-08, 
    -6.250578e-08, -6.238865e-08, -6.210367e-08, -6.230047e-08, 
    -6.222289e-08, -6.240747e-08, -6.252476e-08, -6.246675e-08, 
    -6.282476e-08, -6.268557e-08, -6.341888e-08, -6.310301e-08, -6.39266e-08, 
    -6.372951e-08, -6.397384e-08, -6.384917e-08, -6.406279e-08, 
    -6.387053e-08, -6.420358e-08, -6.427612e-08, -6.422655e-08, 
    -6.441695e-08, -6.385987e-08, -6.40738e-08, -6.246512e-08, -6.247458e-08, 
    -6.251866e-08, -6.232491e-08, -6.231306e-08, -6.213552e-08, 
    -6.229349e-08, -6.236077e-08, -6.253156e-08, -6.263257e-08, -6.27286e-08, 
    -6.293975e-08, -6.317556e-08, -6.350534e-08, -6.374228e-08, 
    -6.390112e-08, -6.380372e-08, -6.388971e-08, -6.379359e-08, 
    -6.374854e-08, -6.424895e-08, -6.396795e-08, -6.438957e-08, 
    -6.436624e-08, -6.417542e-08, -6.436887e-08, -6.248122e-08, 
    -6.242679e-08, -6.223777e-08, -6.238569e-08, -6.211619e-08, 
    -6.226703e-08, -6.235377e-08, -6.268847e-08, -6.276202e-08, 
    -6.283021e-08, -6.296489e-08, -6.313774e-08, -6.344097e-08, 
    -6.370482e-08, -6.394571e-08, -6.392806e-08, -6.393427e-08, 
    -6.398808e-08, -6.385479e-08, -6.400997e-08, -6.403601e-08, 
    -6.396792e-08, -6.436311e-08, -6.425022e-08, -6.436574e-08, 
    -6.429224e-08, -6.244449e-08, -6.253608e-08, -6.248658e-08, 
    -6.257967e-08, -6.251409e-08, -6.280568e-08, -6.289311e-08, 
    -6.330224e-08, -6.313434e-08, -6.340156e-08, -6.316149e-08, 
    -6.320403e-08, -6.341026e-08, -6.317446e-08, -6.369027e-08, 
    -6.334054e-08, -6.399017e-08, -6.36409e-08, -6.401206e-08, -6.394467e-08, 
    -6.405626e-08, -6.415619e-08, -6.428195e-08, -6.451393e-08, 
    -6.446022e-08, -6.465423e-08, -6.267265e-08, -6.279146e-08, 
    -6.278102e-08, -6.290536e-08, -6.299733e-08, -6.319667e-08, -6.35164e-08, 
    -6.339616e-08, -6.361689e-08, -6.366121e-08, -6.332587e-08, 
    -6.353175e-08, -6.2871e-08, -6.297773e-08, -6.291419e-08, -6.268202e-08, 
    -6.342385e-08, -6.304312e-08, -6.37462e-08, -6.353994e-08, -6.414194e-08, 
    -6.384253e-08, -6.443064e-08, -6.468203e-08, -6.491868e-08, -6.51952e-08, 
    -6.285632e-08, -6.277559e-08, -6.292016e-08, -6.312016e-08, 
    -6.330577e-08, -6.355251e-08, -6.357777e-08, -6.362399e-08, 
    -6.374373e-08, -6.384442e-08, -6.363859e-08, -6.386966e-08, 
    -6.300247e-08, -6.345691e-08, -6.274506e-08, -6.295939e-08, 
    -6.310837e-08, -6.304303e-08, -6.338242e-08, -6.346242e-08, 
    -6.378748e-08, -6.361945e-08, -6.461998e-08, -6.417729e-08, 
    -6.540579e-08, -6.506244e-08, -6.274738e-08, -6.285605e-08, 
    -6.323427e-08, -6.305431e-08, -6.356899e-08, -6.369568e-08, 
    -6.379868e-08, -6.393034e-08, -6.394456e-08, -6.402257e-08, 
    -6.389474e-08, -6.401752e-08, -6.355304e-08, -6.37606e-08, -6.319105e-08, 
    -6.332966e-08, -6.326589e-08, -6.319594e-08, -6.341183e-08, 
    -6.364183e-08, -6.364677e-08, -6.372051e-08, -6.392831e-08, 
    -6.357108e-08, -6.467708e-08, -6.399399e-08, -6.297455e-08, 
    -6.318386e-08, -6.321378e-08, -6.313269e-08, -6.368298e-08, 
    -6.348358e-08, -6.402067e-08, -6.387551e-08, -6.411335e-08, 
    -6.399516e-08, -6.397777e-08, -6.382598e-08, -6.373148e-08, 
    -6.349272e-08, -6.329847e-08, -6.314445e-08, -6.318027e-08, 
    -6.334945e-08, -6.365591e-08, -6.394584e-08, -6.388233e-08, 
    -6.409527e-08, -6.353167e-08, -6.376798e-08, -6.367664e-08, 
    -6.391483e-08, -6.339297e-08, -6.383731e-08, -6.327939e-08, 
    -6.332831e-08, -6.347963e-08, -6.378401e-08, -6.385137e-08, 
    -6.392327e-08, -6.387891e-08, -6.366369e-08, -6.362843e-08, 
    -6.347595e-08, -6.343384e-08, -6.331766e-08, -6.322146e-08, 
    -6.330935e-08, -6.340164e-08, -6.366378e-08, -6.390003e-08, 
    -6.415761e-08, -6.422066e-08, -6.452161e-08, -6.427662e-08, 
    -6.468089e-08, -6.433715e-08, -6.493221e-08, -6.386308e-08, 
    -6.432707e-08, -6.348652e-08, -6.357706e-08, -6.374083e-08, -6.41165e-08, 
    -6.39137e-08, -6.415087e-08, -6.362706e-08, -6.335529e-08, -6.328499e-08, 
    -6.315381e-08, -6.328799e-08, -6.327708e-08, -6.340547e-08, 
    -6.336422e-08, -6.367249e-08, -6.35069e-08, -6.397733e-08, -6.414901e-08, 
    -6.463389e-08, -6.493114e-08, -6.523376e-08, -6.536735e-08, 
    -6.540802e-08, -6.542501e-08 ;

 NET_NMIN =
  8.756534e-09, 8.795142e-09, 8.787637e-09, 8.818777e-09, 8.801504e-09, 
    8.821893e-09, 8.764363e-09, 8.796674e-09, 8.776047e-09, 8.76001e-09, 
    8.879208e-09, 8.820166e-09, 8.940552e-09, 8.902892e-09, 8.997502e-09, 
    8.93469e-09, 9.010169e-09, 8.995692e-09, 9.039268e-09, 9.026785e-09, 
    9.082521e-09, 9.04503e-09, 9.111416e-09, 9.073569e-09, 9.079488e-09, 
    9.043793e-09, 8.83205e-09, 8.871857e-09, 8.829691e-09, 8.835367e-09, 
    8.832821e-09, 8.80186e-09, 8.786256e-09, 8.753585e-09, 8.759517e-09, 
    8.783513e-09, 8.83792e-09, 8.819452e-09, 8.865999e-09, 8.864949e-09, 
    8.916772e-09, 8.893406e-09, 8.980515e-09, 8.955756e-09, 9.027305e-09, 
    9.009311e-09, 9.02646e-09, 9.02126e-09, 9.026527e-09, 9.000137e-09, 
    9.011443e-09, 8.988222e-09, 8.897781e-09, 8.924359e-09, 8.845092e-09, 
    8.79743e-09, 8.765779e-09, 8.743318e-09, 8.746493e-09, 8.752546e-09, 
    8.783654e-09, 8.812903e-09, 8.835195e-09, 8.850106e-09, 8.864798e-09, 
    8.909266e-09, 8.932809e-09, 8.985521e-09, 8.976009e-09, 8.992123e-09, 
    9.007521e-09, 9.03337e-09, 9.029115e-09, 9.040503e-09, 8.9917e-09, 
    9.024133e-09, 8.970591e-09, 8.985235e-09, 8.868785e-09, 8.824435e-09, 
    8.805578e-09, 8.78908e-09, 8.748935e-09, 8.776657e-09, 8.765729e-09, 
    8.79173e-09, 8.808251e-09, 8.800081e-09, 8.850513e-09, 8.830906e-09, 
    8.934204e-09, 8.889709e-09, 9.005725e-09, 8.977961e-09, 9.012379e-09, 
    8.994817e-09, 9.024909e-09, 8.997826e-09, 9.044742e-09, 9.05496e-09, 
    9.047977e-09, 9.074798e-09, 8.996325e-09, 9.026459e-09, 8.799852e-09, 
    8.801184e-09, 8.807393e-09, 8.780099e-09, 8.77843e-09, 8.753422e-09, 
    8.775675e-09, 8.785151e-09, 8.809209e-09, 8.823439e-09, 8.836967e-09, 
    8.86671e-09, 8.899929e-09, 8.946384e-09, 8.979761e-09, 9.002135e-09, 
    8.988416e-09, 9.000528e-09, 8.986988e-09, 8.980642e-09, 9.051132e-09, 
    9.011549e-09, 9.070941e-09, 9.067655e-09, 9.040774e-09, 9.068025e-09, 
    8.80212e-09, 8.794451e-09, 8.767825e-09, 8.788662e-09, 8.750698e-09, 
    8.771948e-09, 8.784165e-09, 8.831313e-09, 8.841675e-09, 8.85128e-09, 
    8.870253e-09, 8.894601e-09, 8.937316e-09, 8.974484e-09, 9.008417e-09, 
    9.00593e-09, 9.006806e-09, 9.014386e-09, 8.99561e-09, 9.017469e-09, 
    9.021136e-09, 9.011544e-09, 9.067215e-09, 9.051311e-09, 9.067585e-09, 
    9.057231e-09, 8.796944e-09, 8.809848e-09, 8.802875e-09, 8.815987e-09, 
    8.806749e-09, 8.847825e-09, 8.860141e-09, 8.917773e-09, 8.894122e-09, 
    8.931766e-09, 8.897946e-09, 8.903938e-09, 8.93299e-09, 8.899774e-09, 
    8.972433e-09, 8.92317e-09, 9.01468e-09, 8.96548e-09, 9.017763e-09, 
    9.00827e-09, 9.023989e-09, 9.038065e-09, 9.05578e-09, 9.088459e-09, 
    9.080892e-09, 9.108223e-09, 8.829086e-09, 8.845823e-09, 8.84435e-09, 
    8.861867e-09, 8.874822e-09, 8.902902e-09, 8.94794e-09, 8.931004e-09, 
    8.962098e-09, 8.96834e-09, 8.921102e-09, 8.950104e-09, 8.857025e-09, 
    8.872061e-09, 8.86311e-09, 8.830406e-09, 8.934905e-09, 8.881273e-09, 
    8.980312e-09, 8.951257e-09, 9.036058e-09, 8.993883e-09, 9.076726e-09, 
    9.112139e-09, 9.145475e-09, 9.184426e-09, 8.854959e-09, 8.843586e-09, 
    8.86395e-09, 8.892124e-09, 8.918271e-09, 8.953029e-09, 8.956586e-09, 
    8.963097e-09, 8.979965e-09, 8.994148e-09, 8.965155e-09, 8.997703e-09, 
    8.875547e-09, 8.939561e-09, 8.839286e-09, 8.869478e-09, 8.890464e-09, 
    8.881259e-09, 8.929069e-09, 8.940337e-09, 8.986128e-09, 8.962457e-09, 
    9.103397e-09, 9.041037e-09, 9.21409e-09, 9.165726e-09, 8.839613e-09, 
    8.85492e-09, 8.908198e-09, 8.882848e-09, 8.955349e-09, 8.973196e-09, 
    8.987706e-09, 9.006251e-09, 9.008255e-09, 9.019243e-09, 9.001236e-09, 
    9.018532e-09, 8.953102e-09, 8.982341e-09, 8.902109e-09, 8.921636e-09, 
    8.912654e-09, 8.902799e-09, 8.933212e-09, 8.96561e-09, 8.966305e-09, 
    8.976694e-09, 9.005966e-09, 8.955643e-09, 9.111441e-09, 9.015218e-09, 
    8.871613e-09, 8.901098e-09, 8.905311e-09, 8.893889e-09, 8.971407e-09, 
    8.943318e-09, 9.018975e-09, 8.998528e-09, 9.032031e-09, 9.015382e-09, 
    9.012933e-09, 8.991551e-09, 8.978238e-09, 8.944606e-09, 8.917243e-09, 
    8.895547e-09, 8.900591e-09, 8.924425e-09, 8.967593e-09, 9.008435e-09, 
    8.999488e-09, 9.029485e-09, 8.950092e-09, 8.983381e-09, 8.970514e-09, 
    9.004065e-09, 8.930554e-09, 8.993147e-09, 8.914554e-09, 8.921446e-09, 
    8.942761e-09, 8.985638e-09, 8.995127e-09, 9.005256e-09, 8.999007e-09, 
    8.96869e-09, 8.963724e-09, 8.942243e-09, 8.936311e-09, 8.919946e-09, 
    8.906395e-09, 8.918775e-09, 8.931776e-09, 8.968703e-09, 9.001981e-09, 
    9.038266e-09, 9.047147e-09, 9.089541e-09, 9.05503e-09, 9.111977e-09, 
    9.063557e-09, 9.14738e-09, 8.996777e-09, 9.062137e-09, 8.943732e-09, 
    8.956487e-09, 8.979557e-09, 9.032474e-09, 9.003908e-09, 9.037318e-09, 
    8.963529e-09, 8.925246e-09, 8.915344e-09, 8.896865e-09, 8.915766e-09, 
    8.914229e-09, 8.932316e-09, 8.926504e-09, 8.969929e-09, 8.946603e-09, 
    9.012871e-09, 9.037055e-09, 9.105358e-09, 9.147229e-09, 9.189857e-09, 
    9.208676e-09, 9.214404e-09, 9.216799e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14 ;

 O_SCALAR =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5 ;

 PCH4 =
  0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627 ;

 PCO2 =
  28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  5.065059e-14, 5.07875e-14, 5.076091e-14, 5.087123e-14, 5.081006e-14, 
    5.088227e-14, 5.067837e-14, 5.079292e-14, 5.071982e-14, 5.066294e-14, 
    5.1085e-14, 5.087615e-14, 5.130174e-14, 5.116879e-14, 5.150255e-14, 
    5.128103e-14, 5.154717e-14, 5.149621e-14, 5.164964e-14, 5.160571e-14, 
    5.180164e-14, 5.166991e-14, 5.190315e-14, 5.177022e-14, 5.179101e-14, 
    5.166555e-14, 5.091825e-14, 5.1059e-14, 5.09099e-14, 5.092998e-14, 
    5.092098e-14, 5.081131e-14, 5.075598e-14, 5.064015e-14, 5.066119e-14, 
    5.074628e-14, 5.093901e-14, 5.087365e-14, 5.10384e-14, 5.103468e-14, 
    5.121782e-14, 5.113528e-14, 5.144272e-14, 5.135543e-14, 5.160754e-14, 
    5.154418e-14, 5.160456e-14, 5.158626e-14, 5.16048e-14, 5.151186e-14, 
    5.155169e-14, 5.146989e-14, 5.115073e-14, 5.124461e-14, 5.096441e-14, 
    5.079556e-14, 5.06834e-14, 5.060371e-14, 5.061498e-14, 5.063645e-14, 
    5.074677e-14, 5.085045e-14, 5.092939e-14, 5.098216e-14, 5.103415e-14, 
    5.119125e-14, 5.127441e-14, 5.146034e-14, 5.142685e-14, 5.148361e-14, 
    5.153788e-14, 5.162887e-14, 5.161391e-14, 5.165397e-14, 5.148214e-14, 
    5.159635e-14, 5.140775e-14, 5.145936e-14, 5.104813e-14, 5.089129e-14, 
    5.082445e-14, 5.076601e-14, 5.062364e-14, 5.072197e-14, 5.068321e-14, 
    5.077543e-14, 5.083397e-14, 5.080502e-14, 5.098361e-14, 5.091421e-14, 
    5.127934e-14, 5.11222e-14, 5.153155e-14, 5.143372e-14, 5.155499e-14, 
    5.149313e-14, 5.159909e-14, 5.150374e-14, 5.166889e-14, 5.170481e-14, 
    5.168026e-14, 5.177457e-14, 5.149844e-14, 5.160454e-14, 5.080421e-14, 
    5.080893e-14, 5.083093e-14, 5.073417e-14, 5.072826e-14, 5.063956e-14, 
    5.07185e-14, 5.075209e-14, 5.083737e-14, 5.088776e-14, 5.093566e-14, 
    5.10409e-14, 5.115831e-14, 5.132234e-14, 5.144007e-14, 5.151892e-14, 
    5.147058e-14, 5.151325e-14, 5.146554e-14, 5.144318e-14, 5.169134e-14, 
    5.155205e-14, 5.176101e-14, 5.174946e-14, 5.165492e-14, 5.175076e-14, 
    5.081224e-14, 5.078507e-14, 5.069065e-14, 5.076455e-14, 5.06299e-14, 
    5.070527e-14, 5.074858e-14, 5.091562e-14, 5.095233e-14, 5.098631e-14, 
    5.105343e-14, 5.113951e-14, 5.129034e-14, 5.142145e-14, 5.154104e-14, 
    5.153229e-14, 5.153537e-14, 5.156205e-14, 5.149592e-14, 5.157291e-14, 
    5.158581e-14, 5.155205e-14, 5.174791e-14, 5.169199e-14, 5.174921e-14, 
    5.171281e-14, 5.079391e-14, 5.083963e-14, 5.081492e-14, 5.086136e-14, 
    5.082864e-14, 5.097406e-14, 5.101763e-14, 5.122133e-14, 5.11378e-14, 
    5.127075e-14, 5.115133e-14, 5.117249e-14, 5.127502e-14, 5.115779e-14, 
    5.14142e-14, 5.124037e-14, 5.156309e-14, 5.138965e-14, 5.157395e-14, 
    5.154053e-14, 5.159587e-14, 5.16454e-14, 5.170771e-14, 5.182254e-14, 
    5.179597e-14, 5.189196e-14, 5.090776e-14, 5.096699e-14, 5.09618e-14, 
    5.102377e-14, 5.106958e-14, 5.116884e-14, 5.132784e-14, 5.126809e-14, 
    5.13778e-14, 5.13998e-14, 5.123313e-14, 5.133547e-14, 5.100663e-14, 
    5.105979e-14, 5.102816e-14, 5.091242e-14, 5.128182e-14, 5.109236e-14, 
    5.1442e-14, 5.133955e-14, 5.163833e-14, 5.14898e-14, 5.178133e-14, 
    5.190566e-14, 5.202267e-14, 5.215911e-14, 5.099933e-14, 5.09591e-14, 
    5.103115e-14, 5.113072e-14, 5.122311e-14, 5.13458e-14, 5.135836e-14, 
    5.138131e-14, 5.14408e-14, 5.149077e-14, 5.138855e-14, 5.15033e-14, 
    5.107206e-14, 5.129826e-14, 5.094386e-14, 5.105065e-14, 5.112487e-14, 
    5.109234e-14, 5.126126e-14, 5.130103e-14, 5.146249e-14, 5.137907e-14, 
    5.187496e-14, 5.165582e-14, 5.226298e-14, 5.209362e-14, 5.094503e-14, 
    5.09992e-14, 5.118753e-14, 5.109796e-14, 5.135399e-14, 5.141692e-14, 
    5.146808e-14, 5.15334e-14, 5.154046e-14, 5.157915e-14, 5.151575e-14, 
    5.157666e-14, 5.134606e-14, 5.144916e-14, 5.116605e-14, 5.1235e-14, 
    5.120329e-14, 5.116848e-14, 5.127588e-14, 5.139015e-14, 5.139263e-14, 
    5.142924e-14, 5.153227e-14, 5.135503e-14, 5.190313e-14, 5.156487e-14, 
    5.105825e-14, 5.116242e-14, 5.117735e-14, 5.1137e-14, 5.141061e-14, 
    5.131154e-14, 5.157821e-14, 5.150621e-14, 5.162417e-14, 5.156557e-14, 
    5.155694e-14, 5.148162e-14, 5.14347e-14, 5.131607e-14, 5.121948e-14, 
    5.114286e-14, 5.116068e-14, 5.124484e-14, 5.139715e-14, 5.154109e-14, 
    5.150956e-14, 5.161521e-14, 5.133544e-14, 5.145281e-14, 5.140745e-14, 
    5.152571e-14, 5.126649e-14, 5.148713e-14, 5.121001e-14, 5.123434e-14, 
    5.130957e-14, 5.146074e-14, 5.149423e-14, 5.152989e-14, 5.150789e-14, 
    5.140102e-14, 5.138352e-14, 5.130775e-14, 5.12868e-14, 5.122905e-14, 
    5.118119e-14, 5.12249e-14, 5.127079e-14, 5.140108e-14, 5.151836e-14, 
    5.16461e-14, 5.167735e-14, 5.182628e-14, 5.170501e-14, 5.1905e-14, 
    5.17349e-14, 5.202925e-14, 5.149997e-14, 5.172998e-14, 5.131301e-14, 
    5.135801e-14, 5.143931e-14, 5.162568e-14, 5.152515e-14, 5.164273e-14, 
    5.138283e-14, 5.124772e-14, 5.121279e-14, 5.114751e-14, 5.121429e-14, 
    5.120886e-14, 5.127272e-14, 5.125221e-14, 5.14054e-14, 5.132314e-14, 
    5.155671e-14, 5.164182e-14, 5.188189e-14, 5.202878e-14, 5.217819e-14, 
    5.224405e-14, 5.22641e-14, 5.227248e-14 ;

 POT_F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POT_F_NIT =
  3.862229e-11, 3.895483e-11, 3.889006e-11, 3.915913e-11, 3.900975e-11, 
    3.91861e-11, 3.868957e-11, 3.896803e-11, 3.879014e-11, 3.865213e-11, 
    3.9684e-11, 3.917112e-11, 4.022054e-11, 3.989069e-11, 4.072198e-11, 
    4.016909e-11, 4.083394e-11, 4.070598e-11, 4.109177e-11, 4.098104e-11, 
    4.147654e-11, 4.114291e-11, 4.173464e-11, 4.139675e-11, 4.14495e-11, 
    4.11319e-11, 3.92741e-11, 3.961999e-11, 3.925365e-11, 3.930286e-11, 
    3.928077e-11, 3.901281e-11, 3.887813e-11, 3.85969e-11, 3.864787e-11, 
    3.885446e-11, 3.932497e-11, 3.916492e-11, 3.956894e-11, 3.95598e-11, 
    4.001207e-11, 3.980781e-11, 4.057205e-11, 4.035406e-11, 4.098566e-11, 
    4.082632e-11, 4.097815e-11, 4.093208e-11, 4.097874e-11, 4.07452e-11, 
    4.084516e-11, 4.063998e-11, 3.984608e-11, 4.007857e-11, 3.938724e-11, 
    3.897455e-11, 3.870174e-11, 3.850875e-11, 3.853599e-11, 3.858797e-11, 
    3.885567e-11, 3.910825e-11, 3.930132e-11, 3.943073e-11, 3.955847e-11, 
    3.99464e-11, 4.015257e-11, 4.061618e-11, 4.053232e-11, 4.067444e-11, 
    4.081048e-11, 4.10394e-11, 4.100168e-11, 4.110269e-11, 4.067068e-11, 
    4.095752e-11, 4.048455e-11, 4.061362e-11, 3.959322e-11, 3.920809e-11, 
    3.904494e-11, 3.890246e-11, 3.855695e-11, 3.879537e-11, 3.870129e-11, 
    3.892531e-11, 3.906801e-11, 3.89974e-11, 3.943427e-11, 3.926411e-11, 
    4.01648e-11, 3.977553e-11, 4.079461e-11, 4.054952e-11, 4.085346e-11, 
    4.069822e-11, 4.096439e-11, 4.072479e-11, 4.114031e-11, 4.123111e-11, 
    4.116903e-11, 4.140766e-11, 4.071149e-11, 4.09781e-11, 3.899545e-11, 
    3.900696e-11, 3.906061e-11, 3.882503e-11, 3.881064e-11, 3.859547e-11, 
    3.878689e-11, 3.886856e-11, 3.907629e-11, 3.919942e-11, 3.931666e-11, 
    3.95751e-11, 3.986476e-11, 4.027168e-11, 4.056537e-11, 4.076285e-11, 
    4.06417e-11, 4.074864e-11, 4.062909e-11, 4.057311e-11, 4.119707e-11, 
    4.084608e-11, 4.137328e-11, 4.134403e-11, 4.110505e-11, 4.13473e-11, 
    3.901503e-11, 3.89488e-11, 3.871931e-11, 3.889884e-11, 3.857207e-11, 
    3.875479e-11, 3.886005e-11, 3.926764e-11, 3.93575e-11, 3.944091e-11, 
    3.960593e-11, 3.981822e-11, 4.019208e-11, 4.051885e-11, 4.081839e-11, 
    4.07964e-11, 4.080413e-11, 4.087118e-11, 4.070518e-11, 4.089846e-11, 
    4.093093e-11, 4.084603e-11, 4.134009e-11, 4.119863e-11, 4.134338e-11, 
    4.125124e-11, 3.897032e-11, 3.908181e-11, 3.902153e-11, 3.913491e-11, 
    3.9055e-11, 3.94109e-11, 3.951793e-11, 4.002081e-11, 3.981403e-11, 
    4.014339e-11, 3.984742e-11, 3.989977e-11, 4.015412e-11, 3.986337e-11, 
    4.050077e-11, 4.006803e-11, 4.087378e-11, 4.043953e-11, 4.090106e-11, 
    4.081705e-11, 4.095619e-11, 4.108101e-11, 4.123835e-11, 4.152944e-11, 
    4.146193e-11, 4.170599e-11, 3.924834e-11, 3.939352e-11, 3.938073e-11, 
    3.953295e-11, 3.964572e-11, 3.989074e-11, 4.028535e-11, 4.013671e-11, 
    4.04098e-11, 4.046474e-11, 4.004993e-11, 4.030433e-11, 3.949081e-11, 
    3.962163e-11, 3.954371e-11, 3.925971e-11, 4.017088e-11, 3.970188e-11, 
    4.057018e-11, 4.031442e-11, 4.106318e-11, 4.06899e-11, 4.142479e-11, 
    4.174102e-11, 4.203983e-11, 4.239039e-11, 3.947288e-11, 3.937409e-11, 
    3.955107e-11, 3.97966e-11, 4.002515e-11, 4.033005e-11, 4.036131e-11, 
    4.041858e-11, 4.056714e-11, 4.069228e-11, 4.043668e-11, 4.072366e-11, 
    3.965198e-11, 4.021173e-11, 3.93367e-11, 3.959912e-11, 3.978204e-11, 
    3.970175e-11, 4.011969e-11, 4.021851e-11, 4.062144e-11, 4.041289e-11, 
    4.166283e-11, 4.110735e-11, 4.265837e-11, 4.222189e-11, 3.93396e-11, 
    3.947253e-11, 3.993702e-11, 3.971566e-11, 4.035044e-11, 4.05075e-11, 
    4.063541e-11, 4.079922e-11, 4.081693e-11, 4.091417e-11, 4.075487e-11, 
    4.090787e-11, 4.033065e-11, 4.058806e-11, 3.988374e-11, 4.005456e-11, 
    3.997593e-11, 3.988975e-11, 4.015599e-11, 4.044064e-11, 4.044674e-11, 
    4.053824e-11, 4.079663e-11, 4.035294e-11, 4.173475e-11, 4.087846e-11, 
    3.961775e-11, 3.987494e-11, 3.991176e-11, 3.981198e-11, 4.049172e-11, 
    4.024472e-11, 4.09118e-11, 4.073094e-11, 4.102748e-11, 4.087998e-11, 
    4.085829e-11, 4.066932e-11, 4.055187e-11, 4.025599e-11, 4.001608e-11, 
    3.982639e-11, 3.987045e-11, 4.007897e-11, 4.045808e-11, 4.081846e-11, 
    4.073937e-11, 4.100485e-11, 4.030414e-11, 4.059717e-11, 4.048377e-11, 
    4.07798e-11, 4.013274e-11, 4.068344e-11, 3.99926e-11, 4.005292e-11, 
    4.023982e-11, 4.061715e-11, 4.07009e-11, 4.07904e-11, 4.073515e-11, 
    4.046776e-11, 4.042404e-11, 4.023524e-11, 4.018318e-11, 4.003974e-11, 
    3.992117e-11, 4.002948e-11, 4.014339e-11, 4.046784e-11, 4.07614e-11, 
    4.108272e-11, 4.116157e-11, 4.153903e-11, 4.123162e-11, 4.173952e-11, 
    4.130746e-11, 4.205689e-11, 4.071549e-11, 4.129491e-11, 4.024834e-11, 
    4.036041e-11, 4.056351e-11, 4.10314e-11, 4.077846e-11, 4.107436e-11, 
    4.042233e-11, 4.008617e-11, 3.999945e-11, 3.98379e-11, 4.000314e-11, 
    3.998969e-11, 4.014812e-11, 4.009716e-11, 4.047863e-11, 4.027349e-11, 
    4.085768e-11, 4.107197e-11, 4.168032e-11, 4.205554e-11, 4.243934e-11, 
    4.260935e-11, 4.266116e-11, 4.268283e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.0005835941, 0.0005835972, 0.0005835966, 0.000583599, 0.0005835977, 
    0.0005835993, 0.0005835948, 0.0005835973, 0.0005835957, 0.0005835944, 
    0.0005836036, 0.0005835991, 0.0005836086, 0.0005836057, 0.0005836102, 
    0.0005836081, 0.0005836113, 0.0005836101, 0.0005836136, 0.0005836127, 
    0.0005835862, 0.0005836141, 0.0005835884, 0.0005835856, 0.0005835861, 
    0.000583614, 0.0005836001, 0.000583603, 0.0005835999, 0.0005836003, 
    0.0005836001, 0.0005835977, 0.0005835964, 0.0005835939, 0.0005835944, 
    0.0005835962, 0.0005836005, 0.0005835991, 0.0005836028, 0.0005836027, 
    0.0005836068, 0.0005836049, 0.0005836118, 0.0005836099, 0.0005836127, 
    0.0005836113, 0.0005836126, 0.0005836122, 0.0005836126, 0.0005836105, 
    0.0005836114, 0.0005836125, 0.0005836053, 0.0005836074, 0.0005836011, 
    0.0005835973, 0.0005835948, 0.0005835932, 0.0005835934, 0.0005835939, 
    0.0005835962, 0.0005835986, 0.0005836004, 0.0005836015, 0.0005836027, 
    0.0005836061, 0.000583608, 0.0005836122, 0.0005836115, 0.0005836127, 
    0.0005836111, 0.0005836132, 0.0005836128, 0.0005836137, 0.0005836127, 
    0.0005836124, 0.0005836111, 0.0005836122, 0.0005836028, 0.0005835995, 
    0.0005835979, 0.0005835967, 0.0005835936, 0.0005835957, 0.0005835948, 
    0.0005835969, 0.0005835982, 0.0005835976, 0.0005836015, 0.0005836, 
    0.0005836081, 0.0005836046, 0.000583611, 0.0005836117, 0.0005836115, 
    0.000583613, 0.0005836125, 0.0005836103, 0.000583614, 0.0005835842, 
    0.0005836143, 0.0005835858, 0.0005836102, 0.0005836126, 0.0005835976, 
    0.0005835976, 0.0005835982, 0.0005835959, 0.0005835958, 0.0005835939, 
    0.0005835957, 0.0005835964, 0.0005835983, 0.0005835994, 0.0005836005, 
    0.0005836028, 0.0005836054, 0.0005836091, 0.0005836118, 0.0005836107, 
    0.0005836125, 0.0005836106, 0.0005836124, 0.0005836118, 0.000583584, 
    0.0005836114, 0.0005835855, 0.0005835852, 0.0005836138, 0.0005835852, 
    0.0005835977, 0.0005835972, 0.000583595, 0.0005835967, 0.0005835937, 
    0.0005835954, 0.0005835963, 0.0005836, 0.0005836008, 0.0005836016, 
    0.0005836031, 0.000583605, 0.0005836084, 0.0005836113, 0.0005836112, 
    0.000583611, 0.0005836111, 0.0005836117, 0.0005836101, 0.0005836119, 
    0.0005836122, 0.0005836114, 0.0005835852, 0.000583584, 0.0005835852, 
    0.0005835844, 0.0005835973, 0.0005835983, 0.0005835978, 0.0005835988, 
    0.0005835981, 0.0005836013, 0.0005836022, 0.0005836068, 0.000583605, 
    0.0005836079, 0.0005836053, 0.0005836057, 0.0005836079, 0.0005836054, 
    0.0005836111, 0.0005836072, 0.0005836117, 0.0005836106, 0.0005836119, 
    0.0005836112, 0.0005836124, 0.0005836135, 0.0005835843, 0.0005835867, 
    0.0005835862, 0.0005835883, 0.0005835998, 0.0005836011, 0.0005836011, 
    0.0005836025, 0.0005836035, 0.0005836057, 0.0005836092, 0.0005836079, 
    0.0005836104, 0.0005836108, 0.0005836071, 0.0005836094, 0.0005836021, 
    0.0005836032, 0.0005836025, 0.0005836, 0.0005836082, 0.0005836039, 
    0.0005836118, 0.0005836095, 0.0005836133, 0.0005836129, 0.0005835859, 
    0.0005835885, 0.0005835911, 0.000583594, 0.0005836019, 0.000583601, 
    0.0005836026, 0.0005836048, 0.0005836069, 0.0005836096, 0.0005836099, 
    0.0005836104, 0.0005836118, 0.0005836129, 0.0005836106, 0.0005836103, 
    0.0005836034, 0.0005836086, 0.0005836007, 0.000583603, 0.0005836047, 
    0.000583604, 0.0005836078, 0.0005836086, 0.0005836122, 0.0005836104, 
    0.0005835878, 0.0005836137, 0.0005835963, 0.0005835926, 0.0005836007, 
    0.0005836019, 0.0005836061, 0.0005836041, 0.0005836099, 0.0005836113, 
    0.0005836124, 0.000583611, 0.0005836111, 0.000583612, 0.0005836106, 
    0.000583612, 0.0005836096, 0.000583612, 0.0005836056, 0.0005836072, 
    0.0005836065, 0.0005836057, 0.0005836081, 0.0005836106, 0.0005836107, 
    0.0005836115, 0.0005836107, 0.0005836099, 0.0005835883, 0.0005836115, 
    0.0005836032, 0.0005836055, 0.0005836058, 0.000583605, 0.0005836111, 
    0.0005836089, 0.000583612, 0.0005836104, 0.0005836131, 0.0005836117, 
    0.0005836115, 0.0005836127, 0.0005836117, 0.000583609, 0.0005836068, 
    0.0005836051, 0.0005836055, 0.0005836074, 0.0005836108, 0.0005836111, 
    0.0005836104, 0.0005836129, 0.0005836094, 0.0005836121, 0.000583611, 
    0.0005836108, 0.0005836079, 0.0005836127, 0.0005836066, 0.0005836072, 
    0.0005836088, 0.0005836122, 0.0005836101, 0.0005836109, 0.0005836104, 
    0.0005836108, 0.0005836105, 0.0005836088, 0.0005836083, 0.0005836071, 
    0.000583606, 0.0005836069, 0.0005836079, 0.0005836109, 0.0005836106, 
    0.0005836135, 0.0005836143, 0.0005835867, 0.0005835841, 0.0005835883, 
    0.0005835847, 0.0005835911, 0.0005836101, 0.0005835847, 0.0005836089, 
    0.0005836099, 0.0005836117, 0.000583613, 0.0005836108, 0.0005836134, 
    0.0005836105, 0.0005836074, 0.0005836067, 0.0005836052, 0.0005836067, 
    0.0005836066, 0.0005836081, 0.0005836076, 0.000583611, 0.0005836092, 
    0.0005836115, 0.0005836134, 0.000583588, 0.0005835912, 0.0005835944, 
    0.0005835959, 0.0005835964, 0.0005835965 ;

 QBOT =
  0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_NODYNLNDUSE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_R =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  81.23011, 81.22916, 81.22935, 81.22859, 81.229, 81.22852, 81.2299, 
    81.22913, 81.22962, 81.23001, 81.22716, 81.22855, 81.22562, 81.22652, 
    81.22382, 81.22577, 81.2235, 81.22384, 81.22276, 81.22307, 81.2188, 
    81.22261, 81.21806, 81.219, 81.21886, 81.22265, 81.22826, 81.22734, 
    81.22832, 81.22819, 81.22824, 81.229, 81.22939, 81.23016, 81.23003, 
    81.22945, 81.22813, 81.22856, 81.22742, 81.22745, 81.22619, 81.22675, 
    81.22462, 81.22522, 81.22305, 81.2235, 81.22308, 81.22321, 81.22308, 
    81.22373, 81.22345, 81.22443, 81.22665, 81.22601, 81.22794, 81.22913, 
    81.22987, 81.23042, 81.23034, 81.2302, 81.22945, 81.22872, 81.22817, 
    81.22781, 81.22745, 81.2264, 81.22581, 81.2245, 81.22472, 81.22433, 
    81.22354, 81.22291, 81.22301, 81.22273, 81.22433, 81.22314, 81.22485, 
    81.22449, 81.22742, 81.22844, 81.22894, 81.22931, 81.23029, 81.22961, 
    81.22988, 81.22924, 81.22884, 81.22903, 81.2278, 81.22828, 81.22578, 
    81.22685, 81.22359, 81.22468, 81.22343, 81.22426, 81.22312, 81.22378, 
    81.22263, 81.21946, 81.22255, 81.21896, 81.22382, 81.22308, 81.22904, 
    81.22901, 81.22886, 81.22953, 81.22957, 81.23017, 81.22963, 81.22941, 
    81.22881, 81.22847, 81.22813, 81.22741, 81.22661, 81.22546, 81.22463, 
    81.22367, 81.22441, 81.22372, 81.22445, 81.2246, 81.21956, 81.22345, 
    81.21906, 81.21914, 81.22273, 81.21912, 81.22899, 81.22917, 81.22983, 
    81.22931, 81.23024, 81.22973, 81.22944, 81.22829, 81.22802, 81.22779, 
    81.22732, 81.22672, 81.22569, 81.22477, 81.22352, 81.22358, 81.22356, 
    81.22337, 81.22384, 81.2233, 81.22321, 81.22344, 81.21915, 81.21954, 
    81.21914, 81.21939, 81.22911, 81.2288, 81.22897, 81.22865, 81.22888, 
    81.22789, 81.22759, 81.22617, 81.22674, 81.22582, 81.22665, 81.2265, 
    81.22582, 81.22659, 81.22483, 81.22605, 81.22337, 81.22502, 81.22329, 
    81.22353, 81.22314, 81.22279, 81.21943, 81.21864, 81.21881, 81.21813, 
    81.22832, 81.22793, 81.22795, 81.22752, 81.22721, 81.22652, 81.22542, 
    81.22583, 81.22506, 81.22491, 81.22607, 81.22537, 81.22765, 81.22729, 
    81.2275, 81.2283, 81.22575, 81.22707, 81.22462, 81.22533, 81.22285, 
    81.2243, 81.21892, 81.21806, 81.2172, 81.21626, 81.2277, 81.22797, 
    81.22747, 81.2268, 81.22615, 81.2253, 81.2252, 81.22504, 81.22462, 
    81.22427, 81.22501, 81.22379, 81.22724, 81.22563, 81.22808, 81.22736, 
    81.22684, 81.22706, 81.22588, 81.2256, 81.22449, 81.22505, 81.21828, 
    81.22274, 81.2155, 81.21672, 81.22807, 81.22769, 81.2264, 81.22701, 
    81.22523, 81.22479, 81.22443, 81.22358, 81.22353, 81.22326, 81.22369, 
    81.22327, 81.22529, 81.22457, 81.22653, 81.22607, 81.22628, 81.22652, 
    81.22578, 81.225, 81.22496, 81.22472, 81.22366, 81.22522, 81.21812, 
    81.22342, 81.22729, 81.22659, 81.22646, 81.22674, 81.22484, 81.22553, 
    81.22326, 81.22376, 81.22294, 81.22335, 81.22341, 81.22433, 81.22467, 
    81.2255, 81.22617, 81.22669, 81.22657, 81.226, 81.22495, 81.22353, 
    81.22375, 81.223, 81.22536, 81.22455, 81.22487, 81.22363, 81.22585, 
    81.22436, 81.22623, 81.22606, 81.22555, 81.22451, 81.22385, 81.22361, 
    81.22375, 81.22491, 81.22503, 81.22556, 81.22571, 81.2261, 81.22643, 
    81.22613, 81.22582, 81.22491, 81.22369, 81.22279, 81.22256, 81.21864, 
    81.21948, 81.21812, 81.21932, 81.21721, 81.22385, 81.21931, 81.22552, 
    81.2252, 81.22466, 81.22295, 81.22363, 81.22282, 81.22504, 81.22599, 
    81.22621, 81.22667, 81.2262, 81.22624, 81.22579, 81.22594, 81.22488, 
    81.22544, 81.22342, 81.22283, 81.21822, 81.21718, 81.21609, 81.21562, 
    81.21548, 81.21542 ;

 RH2M_R =
  81.23011, 81.22916, 81.22935, 81.22859, 81.229, 81.22852, 81.2299, 
    81.22913, 81.22962, 81.23001, 81.22716, 81.22855, 81.22562, 81.22652, 
    81.22382, 81.22577, 81.2235, 81.22384, 81.22276, 81.22307, 81.2188, 
    81.22261, 81.21806, 81.219, 81.21886, 81.22265, 81.22826, 81.22734, 
    81.22832, 81.22819, 81.22824, 81.229, 81.22939, 81.23016, 81.23003, 
    81.22945, 81.22813, 81.22856, 81.22742, 81.22745, 81.22619, 81.22675, 
    81.22462, 81.22522, 81.22305, 81.2235, 81.22308, 81.22321, 81.22308, 
    81.22373, 81.22345, 81.22443, 81.22665, 81.22601, 81.22794, 81.22913, 
    81.22987, 81.23042, 81.23034, 81.2302, 81.22945, 81.22872, 81.22817, 
    81.22781, 81.22745, 81.2264, 81.22581, 81.2245, 81.22472, 81.22433, 
    81.22354, 81.22291, 81.22301, 81.22273, 81.22433, 81.22314, 81.22485, 
    81.22449, 81.22742, 81.22844, 81.22894, 81.22931, 81.23029, 81.22961, 
    81.22988, 81.22924, 81.22884, 81.22903, 81.2278, 81.22828, 81.22578, 
    81.22685, 81.22359, 81.22468, 81.22343, 81.22426, 81.22312, 81.22378, 
    81.22263, 81.21946, 81.22255, 81.21896, 81.22382, 81.22308, 81.22904, 
    81.22901, 81.22886, 81.22953, 81.22957, 81.23017, 81.22963, 81.22941, 
    81.22881, 81.22847, 81.22813, 81.22741, 81.22661, 81.22546, 81.22463, 
    81.22367, 81.22441, 81.22372, 81.22445, 81.2246, 81.21956, 81.22345, 
    81.21906, 81.21914, 81.22273, 81.21912, 81.22899, 81.22917, 81.22983, 
    81.22931, 81.23024, 81.22973, 81.22944, 81.22829, 81.22802, 81.22779, 
    81.22732, 81.22672, 81.22569, 81.22477, 81.22352, 81.22358, 81.22356, 
    81.22337, 81.22384, 81.2233, 81.22321, 81.22344, 81.21915, 81.21954, 
    81.21914, 81.21939, 81.22911, 81.2288, 81.22897, 81.22865, 81.22888, 
    81.22789, 81.22759, 81.22617, 81.22674, 81.22582, 81.22665, 81.2265, 
    81.22582, 81.22659, 81.22483, 81.22605, 81.22337, 81.22502, 81.22329, 
    81.22353, 81.22314, 81.22279, 81.21943, 81.21864, 81.21881, 81.21813, 
    81.22832, 81.22793, 81.22795, 81.22752, 81.22721, 81.22652, 81.22542, 
    81.22583, 81.22506, 81.22491, 81.22607, 81.22537, 81.22765, 81.22729, 
    81.2275, 81.2283, 81.22575, 81.22707, 81.22462, 81.22533, 81.22285, 
    81.2243, 81.21892, 81.21806, 81.2172, 81.21626, 81.2277, 81.22797, 
    81.22747, 81.2268, 81.22615, 81.2253, 81.2252, 81.22504, 81.22462, 
    81.22427, 81.22501, 81.22379, 81.22724, 81.22563, 81.22808, 81.22736, 
    81.22684, 81.22706, 81.22588, 81.2256, 81.22449, 81.22505, 81.21828, 
    81.22274, 81.2155, 81.21672, 81.22807, 81.22769, 81.2264, 81.22701, 
    81.22523, 81.22479, 81.22443, 81.22358, 81.22353, 81.22326, 81.22369, 
    81.22327, 81.22529, 81.22457, 81.22653, 81.22607, 81.22628, 81.22652, 
    81.22578, 81.225, 81.22496, 81.22472, 81.22366, 81.22522, 81.21812, 
    81.22342, 81.22729, 81.22659, 81.22646, 81.22674, 81.22484, 81.22553, 
    81.22326, 81.22376, 81.22294, 81.22335, 81.22341, 81.22433, 81.22467, 
    81.2255, 81.22617, 81.22669, 81.22657, 81.226, 81.22495, 81.22353, 
    81.22375, 81.223, 81.22536, 81.22455, 81.22487, 81.22363, 81.22585, 
    81.22436, 81.22623, 81.22606, 81.22555, 81.22451, 81.22385, 81.22361, 
    81.22375, 81.22491, 81.22503, 81.22556, 81.22571, 81.2261, 81.22643, 
    81.22613, 81.22582, 81.22491, 81.22369, 81.22279, 81.22256, 81.21864, 
    81.21948, 81.21812, 81.21932, 81.21721, 81.22385, 81.21931, 81.22552, 
    81.2252, 81.22466, 81.22295, 81.22363, 81.22282, 81.22504, 81.22599, 
    81.22621, 81.22667, 81.2262, 81.22624, 81.22579, 81.22594, 81.22488, 
    81.22544, 81.22342, 81.22283, 81.21822, 81.21718, 81.21609, 81.21562, 
    81.21548, 81.21542 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RSCANOPY =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SABG =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004381193, 0.0004399699, 0.00043961, 0.0004411027, 0.0004402746, 
    0.0004412519, 0.0004384942, 0.000440043, 0.0004390542, 0.0004382854, 
    0.0004439988, 0.0004411688, 0.0004469388, 0.0004451337, 0.000449668, 
    0.0004466577, 0.000450275, 0.0004495811, 0.0004516694, 0.000451071, 
    0.000453742, 0.0004519454, 0.0004551266, 0.000453313, 0.0004535966, 
    0.0004518858, 0.0004417388, 0.0004436469, 0.0004416256, 0.0004418977, 
    0.0004417756, 0.0004402914, 0.0004395435, 0.0004379773, 0.0004382616, 
    0.0004394119, 0.0004420197, 0.0004411344, 0.0004433654, 0.000443315, 
    0.0004457988, 0.0004446789, 0.0004488537, 0.000447667, 0.000451096, 
    0.0004502335, 0.0004510553, 0.0004508061, 0.0004510584, 0.0004497937, 
    0.0004503354, 0.0004492226, 0.0004448892, 0.000446163, 0.0004423637, 
    0.0004400791, 0.0004385619, 0.0004374853, 0.0004376373, 0.0004379275, 
    0.0004394185, 0.0004408205, 0.0004418889, 0.0004426035, 0.0004433076, 
    0.000445439, 0.0004465673, 0.0004490935, 0.0004486376, 0.0004494098, 
    0.0004501477, 0.0004513864, 0.0004511825, 0.0004517281, 0.0004493892, 
    0.0004509436, 0.0004483775, 0.0004490793, 0.0004434994, 0.0004413735, 
    0.0004404697, 0.0004396787, 0.0004377543, 0.0004390832, 0.0004385593, 
    0.0004398055, 0.0004405974, 0.0004402057, 0.000442623, 0.0004416831, 
    0.0004466341, 0.0004445015, 0.0004500617, 0.000448731, 0.0004503804, 
    0.0004495388, 0.0004509808, 0.0004496829, 0.0004519311, 0.0004524209, 
    0.000452086, 0.0004533714, 0.0004496106, 0.0004510547, 0.000440195, 
    0.0004402589, 0.0004405564, 0.0004392481, 0.0004391681, 0.0004379692, 
    0.0004390359, 0.0004394901, 0.0004406432, 0.0004413252, 0.0004419735, 
    0.0004433991, 0.0004449912, 0.0004472176, 0.0004488172, 0.0004498894, 
    0.0004492319, 0.0004498123, 0.0004491633, 0.0004488592, 0.0004522373, 
    0.0004503403, 0.0004531864, 0.000453029, 0.0004517407, 0.0004530466, 
    0.0004403036, 0.000439936, 0.0004386597, 0.0004396584, 0.0004378385, 
    0.0004388572, 0.0004394427, 0.0004417026, 0.0004421991, 0.0004426595, 
    0.0004435688, 0.0004447357, 0.000446783, 0.0004485642, 0.0004501904, 
    0.0004500712, 0.0004501131, 0.0004504762, 0.0004495764, 0.0004506239, 
    0.0004507996, 0.0004503399, 0.0004530077, 0.0004522456, 0.0004530254, 
    0.0004525291, 0.0004400554, 0.0004406738, 0.0004403395, 0.000440968, 
    0.0004405251, 0.000442494, 0.0004430842, 0.0004458464, 0.0004447128, 
    0.000446517, 0.0004448959, 0.0004451832, 0.0004465755, 0.0004449834, 
    0.0004484658, 0.0004461046, 0.0004504903, 0.0004481323, 0.0004506379, 
    0.0004501829, 0.0004509361, 0.0004516108, 0.0004524596, 0.0004540256, 
    0.0004536629, 0.0004549726, 0.0004415959, 0.000442398, 0.0004423274, 
    0.0004431669, 0.0004437878, 0.0004451337, 0.0004472922, 0.0004464804, 
    0.0004479706, 0.0004482697, 0.0004460056, 0.0004473956, 0.0004429344, 
    0.000443655, 0.000443226, 0.0004416583, 0.0004466669, 0.0004440963, 
    0.000448843, 0.0004474504, 0.0004515144, 0.0004494932, 0.0004534632, 
    0.0004551602, 0.0004567575, 0.0004586239, 0.0004428359, 0.0004422907, 
    0.0004432667, 0.0004446171, 0.0004458701, 0.000447536, 0.0004477064, 
    0.0004480183, 0.0004488267, 0.0004495064, 0.0004481169, 0.0004496766, 
    0.000443822, 0.00044689, 0.0004420838, 0.000443531, 0.0004445367, 
    0.0004440956, 0.0004463869, 0.0004469269, 0.0004491214, 0.000447987, 
    0.0004547412, 0.0004517528, 0.0004600451, 0.0004577277, 0.0004421001, 
    0.0004428338, 0.0004453873, 0.0004441723, 0.000447647, 0.0004485024, 
    0.0004491976, 0.0004500864, 0.0004501823, 0.0004507089, 0.0004498458, 
    0.0004506747, 0.0004475389, 0.0004489402, 0.0004450949, 0.0004460307, 
    0.0004456001, 0.0004451278, 0.0004465853, 0.0004481381, 0.0004481713, 
    0.0004486691, 0.000450072, 0.0004476601, 0.0004551265, 0.0004505152, 
    0.0004436338, 0.0004450469, 0.0004452488, 0.0004447014, 0.0004484165, 
    0.0004470703, 0.0004506961, 0.0004497161, 0.0004513216, 0.0004505238, 
    0.0004504063, 0.0004493815, 0.0004487434, 0.0004471316, 0.00044582, 
    0.0004447801, 0.0004450218, 0.0004461641, 0.000448233, 0.0004501903, 
    0.0004497614, 0.0004511989, 0.000447394, 0.0004489894, 0.0004483726, 
    0.0004499806, 0.0004464586, 0.0004494585, 0.0004456917, 0.0004460219, 
    0.0004470434, 0.0004490984, 0.000449553, 0.0004500384, 0.0004497388, 
    0.0004482859, 0.0004480478, 0.0004470182, 0.0004467339, 0.0004459495, 
    0.0004452999, 0.0004458933, 0.0004465163, 0.0004482861, 0.0004498809, 
    0.0004516197, 0.0004520452, 0.0004540768, 0.000452423, 0.0004551519, 
    0.0004528316, 0.0004568482, 0.0004496323, 0.0004527646, 0.0004470899, 
    0.0004477012, 0.0004488068, 0.0004513428, 0.0004499737, 0.0004515748, 
    0.0004480385, 0.0004462036, 0.0004457289, 0.0004448433, 0.0004457491, 
    0.0004456754, 0.0004465422, 0.0004462635, 0.0004483447, 0.0004472267, 
    0.0004504026, 0.0004515615, 0.0004548347, 0.000456841, 0.0004588835, 
    0.0004597852, 0.0004600596, 0.0004601743 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.516111e-14, 3.525612e-14, 3.523766e-14, 3.531423e-14, 3.527177e-14, 
    3.532189e-14, 3.518039e-14, 3.525988e-14, 3.520915e-14, 3.516968e-14, 
    3.546258e-14, 3.531764e-14, 3.561299e-14, 3.552072e-14, 3.575234e-14, 
    3.559862e-14, 3.578331e-14, 3.574794e-14, 3.585442e-14, 3.582393e-14, 
    3.59599e-14, 3.586848e-14, 3.603035e-14, 3.59381e-14, 3.595252e-14, 
    3.586546e-14, 3.534686e-14, 3.544453e-14, 3.534106e-14, 3.5355e-14, 
    3.534875e-14, 3.527264e-14, 3.523424e-14, 3.515386e-14, 3.516847e-14, 
    3.522751e-14, 3.536126e-14, 3.53159e-14, 3.543024e-14, 3.542766e-14, 
    3.555475e-14, 3.549747e-14, 3.571082e-14, 3.565024e-14, 3.58252e-14, 
    3.578123e-14, 3.582313e-14, 3.581044e-14, 3.58233e-14, 3.575881e-14, 
    3.578644e-14, 3.572968e-14, 3.550819e-14, 3.557334e-14, 3.537889e-14, 
    3.526171e-14, 3.518387e-14, 3.512857e-14, 3.513639e-14, 3.515129e-14, 
    3.522786e-14, 3.529981e-14, 3.535459e-14, 3.539121e-14, 3.542729e-14, 
    3.553631e-14, 3.559402e-14, 3.572305e-14, 3.569981e-14, 3.57392e-14, 
    3.577686e-14, 3.584001e-14, 3.582962e-14, 3.585742e-14, 3.573818e-14, 
    3.581744e-14, 3.568656e-14, 3.572237e-14, 3.543699e-14, 3.532815e-14, 
    3.528176e-14, 3.524121e-14, 3.51424e-14, 3.521064e-14, 3.518375e-14, 
    3.524774e-14, 3.528837e-14, 3.526828e-14, 3.539221e-14, 3.534405e-14, 
    3.559744e-14, 3.548839e-14, 3.577247e-14, 3.570458e-14, 3.578873e-14, 
    3.574581e-14, 3.581934e-14, 3.575317e-14, 3.586778e-14, 3.58927e-14, 
    3.587567e-14, 3.594111e-14, 3.574949e-14, 3.582312e-14, 3.526771e-14, 
    3.527099e-14, 3.528626e-14, 3.521911e-14, 3.521501e-14, 3.515346e-14, 
    3.520824e-14, 3.523155e-14, 3.529073e-14, 3.53257e-14, 3.535894e-14, 
    3.543197e-14, 3.551345e-14, 3.562728e-14, 3.570898e-14, 3.57637e-14, 
    3.573016e-14, 3.575977e-14, 3.572666e-14, 3.571114e-14, 3.588336e-14, 
    3.578669e-14, 3.59317e-14, 3.592369e-14, 3.585808e-14, 3.592459e-14, 
    3.527329e-14, 3.525444e-14, 3.518891e-14, 3.52402e-14, 3.514675e-14, 
    3.519906e-14, 3.522911e-14, 3.534503e-14, 3.537051e-14, 3.539409e-14, 
    3.544067e-14, 3.55004e-14, 3.560508e-14, 3.569606e-14, 3.577905e-14, 
    3.577298e-14, 3.577512e-14, 3.579363e-14, 3.574774e-14, 3.580117e-14, 
    3.581012e-14, 3.578669e-14, 3.592261e-14, 3.588381e-14, 3.592352e-14, 
    3.589826e-14, 3.526057e-14, 3.52923e-14, 3.527515e-14, 3.530738e-14, 
    3.528467e-14, 3.538559e-14, 3.541582e-14, 3.555718e-14, 3.549922e-14, 
    3.559148e-14, 3.55086e-14, 3.552329e-14, 3.559444e-14, 3.551309e-14, 
    3.569103e-14, 3.55704e-14, 3.579436e-14, 3.5674e-14, 3.580189e-14, 
    3.57787e-14, 3.58171e-14, 3.585147e-14, 3.589472e-14, 3.597441e-14, 
    3.595596e-14, 3.602258e-14, 3.533958e-14, 3.538068e-14, 3.537708e-14, 
    3.542009e-14, 3.545188e-14, 3.552076e-14, 3.56311e-14, 3.558963e-14, 
    3.566577e-14, 3.568104e-14, 3.556537e-14, 3.563639e-14, 3.540819e-14, 
    3.544508e-14, 3.542313e-14, 3.534281e-14, 3.559917e-14, 3.546769e-14, 
    3.571033e-14, 3.563922e-14, 3.584657e-14, 3.57435e-14, 3.59458e-14, 
    3.603208e-14, 3.611329e-14, 3.620797e-14, 3.540312e-14, 3.53752e-14, 
    3.542521e-14, 3.549431e-14, 3.555842e-14, 3.564356e-14, 3.565228e-14, 
    3.566821e-14, 3.570949e-14, 3.574417e-14, 3.567323e-14, 3.575286e-14, 
    3.54536e-14, 3.561058e-14, 3.536463e-14, 3.543874e-14, 3.549024e-14, 
    3.546767e-14, 3.558489e-14, 3.561249e-14, 3.572454e-14, 3.566665e-14, 
    3.601078e-14, 3.585871e-14, 3.628005e-14, 3.616252e-14, 3.536544e-14, 
    3.540304e-14, 3.553373e-14, 3.547157e-14, 3.564925e-14, 3.569292e-14, 
    3.572842e-14, 3.577375e-14, 3.577865e-14, 3.58055e-14, 3.57615e-14, 
    3.580377e-14, 3.564374e-14, 3.571529e-14, 3.551882e-14, 3.556667e-14, 
    3.554467e-14, 3.552051e-14, 3.559504e-14, 3.567434e-14, 3.567606e-14, 
    3.570147e-14, 3.577297e-14, 3.564997e-14, 3.603033e-14, 3.579559e-14, 
    3.544401e-14, 3.55163e-14, 3.552666e-14, 3.549866e-14, 3.568854e-14, 
    3.561979e-14, 3.580485e-14, 3.575488e-14, 3.583674e-14, 3.579607e-14, 
    3.579009e-14, 3.573782e-14, 3.570525e-14, 3.562294e-14, 3.55559e-14, 
    3.550273e-14, 3.55151e-14, 3.55735e-14, 3.56792e-14, 3.577909e-14, 
    3.575721e-14, 3.583053e-14, 3.563638e-14, 3.571783e-14, 3.568635e-14, 
    3.576841e-14, 3.558852e-14, 3.574164e-14, 3.554933e-14, 3.556622e-14, 
    3.561842e-14, 3.572333e-14, 3.574657e-14, 3.577132e-14, 3.575605e-14, 
    3.568188e-14, 3.566974e-14, 3.561716e-14, 3.560262e-14, 3.556254e-14, 
    3.552933e-14, 3.555967e-14, 3.559151e-14, 3.568193e-14, 3.576331e-14, 
    3.585196e-14, 3.587365e-14, 3.5977e-14, 3.589284e-14, 3.603163e-14, 
    3.591358e-14, 3.611785e-14, 3.575055e-14, 3.591017e-14, 3.562081e-14, 
    3.565204e-14, 3.570846e-14, 3.583779e-14, 3.576803e-14, 3.584963e-14, 
    3.566927e-14, 3.55755e-14, 3.555126e-14, 3.550595e-14, 3.55523e-14, 
    3.554853e-14, 3.559285e-14, 3.557861e-14, 3.568493e-14, 3.562784e-14, 
    3.578993e-14, 3.584899e-14, 3.601559e-14, 3.611753e-14, 3.622121e-14, 
    3.626692e-14, 3.628083e-14, 3.628664e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.169146e-14, 1.172309e-14, 1.171694e-14, 1.174243e-14, 1.17283e-14, 
    1.174498e-14, 1.169788e-14, 1.172434e-14, 1.170745e-14, 1.169432e-14, 
    1.179181e-14, 1.174357e-14, 1.184187e-14, 1.181116e-14, 1.188826e-14, 
    1.183709e-14, 1.189857e-14, 1.188679e-14, 1.192224e-14, 1.191209e-14, 
    1.195735e-14, 1.192692e-14, 1.19808e-14, 1.195009e-14, 1.195489e-14, 
    1.192591e-14, 1.175329e-14, 1.17858e-14, 1.175136e-14, 1.1756e-14, 
    1.175392e-14, 1.172859e-14, 1.171581e-14, 1.168905e-14, 1.169391e-14, 
    1.171357e-14, 1.175809e-14, 1.174299e-14, 1.178104e-14, 1.178018e-14, 
    1.182249e-14, 1.180342e-14, 1.187444e-14, 1.185428e-14, 1.191251e-14, 
    1.189788e-14, 1.191182e-14, 1.19076e-14, 1.191188e-14, 1.189041e-14, 
    1.189961e-14, 1.188071e-14, 1.180699e-14, 1.182868e-14, 1.176395e-14, 
    1.172495e-14, 1.169904e-14, 1.168063e-14, 1.168324e-14, 1.16882e-14, 
    1.171368e-14, 1.173763e-14, 1.175586e-14, 1.176805e-14, 1.178006e-14, 
    1.181635e-14, 1.183556e-14, 1.187851e-14, 1.187077e-14, 1.188388e-14, 
    1.189642e-14, 1.191744e-14, 1.191398e-14, 1.192324e-14, 1.188355e-14, 
    1.190993e-14, 1.186636e-14, 1.187828e-14, 1.178329e-14, 1.174706e-14, 
    1.173162e-14, 1.171812e-14, 1.168524e-14, 1.170795e-14, 1.1699e-14, 
    1.17203e-14, 1.173382e-14, 1.172714e-14, 1.176839e-14, 1.175236e-14, 
    1.18367e-14, 1.18004e-14, 1.189496e-14, 1.187236e-14, 1.190037e-14, 
    1.188608e-14, 1.191056e-14, 1.188853e-14, 1.192668e-14, 1.193498e-14, 
    1.192931e-14, 1.195109e-14, 1.188731e-14, 1.191182e-14, 1.172695e-14, 
    1.172804e-14, 1.173312e-14, 1.171077e-14, 1.17094e-14, 1.168892e-14, 
    1.170715e-14, 1.171491e-14, 1.173461e-14, 1.174625e-14, 1.175731e-14, 
    1.178162e-14, 1.180874e-14, 1.184663e-14, 1.187383e-14, 1.189204e-14, 
    1.188087e-14, 1.189073e-14, 1.187971e-14, 1.187455e-14, 1.193187e-14, 
    1.189969e-14, 1.194796e-14, 1.194529e-14, 1.192345e-14, 1.194559e-14, 
    1.17288e-14, 1.172253e-14, 1.170072e-14, 1.171779e-14, 1.168668e-14, 
    1.170409e-14, 1.17141e-14, 1.175268e-14, 1.176116e-14, 1.176901e-14, 
    1.178452e-14, 1.18044e-14, 1.183924e-14, 1.186953e-14, 1.189715e-14, 
    1.189513e-14, 1.189584e-14, 1.1902e-14, 1.188673e-14, 1.190451e-14, 
    1.190749e-14, 1.189969e-14, 1.194494e-14, 1.193202e-14, 1.194524e-14, 
    1.193683e-14, 1.172457e-14, 1.173513e-14, 1.172942e-14, 1.174015e-14, 
    1.173259e-14, 1.176618e-14, 1.177624e-14, 1.18233e-14, 1.1804e-14, 
    1.183471e-14, 1.180713e-14, 1.181202e-14, 1.18357e-14, 1.180862e-14, 
    1.186785e-14, 1.18277e-14, 1.190224e-14, 1.186218e-14, 1.190475e-14, 
    1.189703e-14, 1.190982e-14, 1.192126e-14, 1.193565e-14, 1.196218e-14, 
    1.195604e-14, 1.197821e-14, 1.175087e-14, 1.176455e-14, 1.176335e-14, 
    1.177767e-14, 1.178825e-14, 1.181117e-14, 1.18479e-14, 1.18341e-14, 
    1.185944e-14, 1.186453e-14, 1.182602e-14, 1.184966e-14, 1.177371e-14, 
    1.178598e-14, 1.177868e-14, 1.175194e-14, 1.183727e-14, 1.179351e-14, 
    1.187427e-14, 1.185061e-14, 1.191962e-14, 1.188531e-14, 1.195266e-14, 
    1.198138e-14, 1.200841e-14, 1.203992e-14, 1.177202e-14, 1.176273e-14, 
    1.177937e-14, 1.180237e-14, 1.182371e-14, 1.185205e-14, 1.185495e-14, 
    1.186025e-14, 1.187399e-14, 1.188554e-14, 1.186192e-14, 1.188843e-14, 
    1.178882e-14, 1.184107e-14, 1.175921e-14, 1.178387e-14, 1.180102e-14, 
    1.17935e-14, 1.183252e-14, 1.184171e-14, 1.187901e-14, 1.185974e-14, 
    1.197428e-14, 1.192366e-14, 1.206392e-14, 1.202479e-14, 1.175948e-14, 
    1.177199e-14, 1.181549e-14, 1.17948e-14, 1.185394e-14, 1.186848e-14, 
    1.18803e-14, 1.189538e-14, 1.189702e-14, 1.190595e-14, 1.189131e-14, 
    1.190538e-14, 1.185211e-14, 1.187593e-14, 1.181053e-14, 1.182646e-14, 
    1.181913e-14, 1.181109e-14, 1.18359e-14, 1.186229e-14, 1.186287e-14, 
    1.187133e-14, 1.189513e-14, 1.185418e-14, 1.198079e-14, 1.190265e-14, 
    1.178563e-14, 1.180969e-14, 1.181314e-14, 1.180382e-14, 1.186702e-14, 
    1.184414e-14, 1.190574e-14, 1.18891e-14, 1.191635e-14, 1.190282e-14, 
    1.190082e-14, 1.188343e-14, 1.187259e-14, 1.184518e-14, 1.182287e-14, 
    1.180517e-14, 1.180929e-14, 1.182873e-14, 1.186391e-14, 1.189716e-14, 
    1.188988e-14, 1.191428e-14, 1.184966e-14, 1.187677e-14, 1.186629e-14, 
    1.189361e-14, 1.183373e-14, 1.18847e-14, 1.182068e-14, 1.18263e-14, 
    1.184368e-14, 1.18786e-14, 1.188634e-14, 1.189457e-14, 1.188949e-14, 
    1.186481e-14, 1.186076e-14, 1.184326e-14, 1.183842e-14, 1.182508e-14, 
    1.181403e-14, 1.182412e-14, 1.183472e-14, 1.186482e-14, 1.189191e-14, 
    1.192142e-14, 1.192864e-14, 1.196304e-14, 1.193503e-14, 1.198122e-14, 
    1.194193e-14, 1.200992e-14, 1.188766e-14, 1.194079e-14, 1.184448e-14, 
    1.185487e-14, 1.187365e-14, 1.19167e-14, 1.189348e-14, 1.192064e-14, 
    1.186061e-14, 1.18294e-14, 1.182133e-14, 1.180625e-14, 1.182167e-14, 
    1.182042e-14, 1.183517e-14, 1.183043e-14, 1.186582e-14, 1.184682e-14, 
    1.190077e-14, 1.192043e-14, 1.197588e-14, 1.200982e-14, 1.204433e-14, 
    1.205955e-14, 1.206418e-14, 1.206611e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.178544e-11, -8.214632e-11, -8.207617e-11, -8.236724e-11, -8.220578e-11, 
    -8.239637e-11, -8.185861e-11, -8.216063e-11, -8.196783e-11, 
    -8.181793e-11, -8.293211e-11, -8.238023e-11, -8.350552e-11, -8.31535e-11, 
    -8.403786e-11, -8.345073e-11, -8.415626e-11, -8.402094e-11, 
    -8.442827e-11, -8.431158e-11, -8.483258e-11, -8.448213e-11, 
    -8.510268e-11, -8.47489e-11, -8.480423e-11, -8.447057e-11, -8.249131e-11, 
    -8.28634e-11, -8.246925e-11, -8.252232e-11, -8.249851e-11, -8.220911e-11, 
    -8.206325e-11, -8.175786e-11, -8.181331e-11, -8.203762e-11, 
    -8.254617e-11, -8.237355e-11, -8.280865e-11, -8.279882e-11, 
    -8.328323e-11, -8.306482e-11, -8.387908e-11, -8.364764e-11, 
    -8.431645e-11, -8.414824e-11, -8.430855e-11, -8.425994e-11, 
    -8.430918e-11, -8.406249e-11, -8.416818e-11, -8.395112e-11, 
    -8.310572e-11, -8.335416e-11, -8.261321e-11, -8.21677e-11, -8.187185e-11, 
    -8.166191e-11, -8.169158e-11, -8.174816e-11, -8.203893e-11, 
    -8.231234e-11, -8.25207e-11, -8.266007e-11, -8.279741e-11, -8.321308e-11, 
    -8.343314e-11, -8.392586e-11, -8.383696e-11, -8.398758e-11, 
    -8.413151e-11, -8.437313e-11, -8.433337e-11, -8.443982e-11, 
    -8.398363e-11, -8.42868e-11, -8.378631e-11, -8.392319e-11, -8.283468e-11, 
    -8.242013e-11, -8.224387e-11, -8.208965e-11, -8.171441e-11, 
    -8.197353e-11, -8.187138e-11, -8.211443e-11, -8.226885e-11, 
    -8.219248e-11, -8.266389e-11, -8.248061e-11, -8.344618e-11, 
    -8.303026e-11, -8.411472e-11, -8.385521e-11, -8.417693e-11, 
    -8.401276e-11, -8.429405e-11, -8.404089e-11, -8.447944e-11, 
    -8.457496e-11, -8.450968e-11, -8.476039e-11, -8.402686e-11, 
    -8.430854e-11, -8.219034e-11, -8.220279e-11, -8.226082e-11, 
    -8.200571e-11, -8.199011e-11, -8.175634e-11, -8.196435e-11, 
    -8.205293e-11, -8.227781e-11, -8.241082e-11, -8.253727e-11, 
    -8.281529e-11, -8.31258e-11, -8.356003e-11, -8.387203e-11, -8.408117e-11, 
    -8.395293e-11, -8.406614e-11, -8.393958e-11, -8.388026e-11, 
    -8.453917e-11, -8.416916e-11, -8.472433e-11, -8.469362e-11, 
    -8.444235e-11, -8.469708e-11, -8.221154e-11, -8.213986e-11, 
    -8.189097e-11, -8.208575e-11, -8.173089e-11, -8.192951e-11, 
    -8.204372e-11, -8.248442e-11, -8.258128e-11, -8.267106e-11, -8.28484e-11, 
    -8.3076e-11, -8.347528e-11, -8.38227e-11, -8.413989e-11, -8.411664e-11, 
    -8.412483e-11, -8.419568e-11, -8.402017e-11, -8.42245e-11, -8.425878e-11, 
    -8.416912e-11, -8.468951e-11, -8.454085e-11, -8.469297e-11, 
    -8.459617e-11, -8.216316e-11, -8.228378e-11, -8.22186e-11, -8.234115e-11, 
    -8.225481e-11, -8.263876e-11, -8.275388e-11, -8.32926e-11, -8.307151e-11, 
    -8.342339e-11, -8.310726e-11, -8.316327e-11, -8.343484e-11, 
    -8.312435e-11, -8.380353e-11, -8.334304e-11, -8.419843e-11, 
    -8.373853e-11, -8.422725e-11, -8.413852e-11, -8.428545e-11, 
    -8.441703e-11, -8.458262e-11, -8.488809e-11, -8.481735e-11, 
    -8.507283e-11, -8.24636e-11, -8.262005e-11, -8.260628e-11, -8.277002e-11, 
    -8.289111e-11, -8.315359e-11, -8.357458e-11, -8.341627e-11, 
    -8.370692e-11, -8.376527e-11, -8.332371e-11, -8.35948e-11, -8.272476e-11, 
    -8.286531e-11, -8.278164e-11, -8.247594e-11, -8.345274e-11, 
    -8.295142e-11, -8.387718e-11, -8.360558e-11, -8.439827e-11, 
    -8.400403e-11, -8.477841e-11, -8.510943e-11, -8.542105e-11, 
    -8.578516e-11, -8.270545e-11, -8.259914e-11, -8.27895e-11, -8.305285e-11, 
    -8.329724e-11, -8.362214e-11, -8.36554e-11, -8.371626e-11, -8.387394e-11, 
    -8.40065e-11, -8.37355e-11, -8.403974e-11, -8.289788e-11, -8.349626e-11, 
    -8.255894e-11, -8.284116e-11, -8.303733e-11, -8.295128e-11, 
    -8.339818e-11, -8.350351e-11, -8.393154e-11, -8.371028e-11, 
    -8.502772e-11, -8.444481e-11, -8.606244e-11, -8.561035e-11, 
    -8.256199e-11, -8.270509e-11, -8.320309e-11, -8.296614e-11, 
    -8.364384e-11, -8.381066e-11, -8.394629e-11, -8.411964e-11, 
    -8.413837e-11, -8.424108e-11, -8.407276e-11, -8.423444e-11, 
    -8.362284e-11, -8.389614e-11, -8.314618e-11, -8.332871e-11, 
    -8.324474e-11, -8.315263e-11, -8.343691e-11, -8.373976e-11, 
    -8.374625e-11, -8.384336e-11, -8.411698e-11, -8.364659e-11, 
    -8.510292e-11, -8.420346e-11, -8.286112e-11, -8.313672e-11, 
    -8.317611e-11, -8.306934e-11, -8.379394e-11, -8.353138e-11, 
    -8.423858e-11, -8.404745e-11, -8.436062e-11, -8.4205e-11, -8.41821e-11, 
    -8.398223e-11, -8.385779e-11, -8.354342e-11, -8.328764e-11, 
    -8.308483e-11, -8.313199e-11, -8.335477e-11, -8.375829e-11, 
    -8.414006e-11, -8.405642e-11, -8.433682e-11, -8.35947e-11, -8.390587e-11, 
    -8.37856e-11, -8.409921e-11, -8.341206e-11, -8.399714e-11, -8.326251e-11, 
    -8.332692e-11, -8.352617e-11, -8.392696e-11, -8.401566e-11, 
    -8.411034e-11, -8.405193e-11, -8.376853e-11, -8.372211e-11, 
    -8.352133e-11, -8.346588e-11, -8.33129e-11, -8.318624e-11, -8.330196e-11, 
    -8.342349e-11, -8.376866e-11, -8.407974e-11, -8.44189e-11, -8.450192e-11, 
    -8.48982e-11, -8.45756e-11, -8.510793e-11, -8.465531e-11, -8.543886e-11, 
    -8.403108e-11, -8.464204e-11, -8.353524e-11, -8.365447e-11, 
    -8.387011e-11, -8.436477e-11, -8.409774e-11, -8.441003e-11, -8.37203e-11, 
    -8.336245e-11, -8.326988e-11, -8.309716e-11, -8.327384e-11, 
    -8.325947e-11, -8.342853e-11, -8.33742e-11, -8.378012e-11, -8.356208e-11, 
    -8.418152e-11, -8.440758e-11, -8.504605e-11, -8.543745e-11, 
    -8.583592e-11, -8.601184e-11, -8.606538e-11, -8.608777e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -1.971184e-12, -1.97988e-12, -1.978189e-12, -1.985203e-12, -1.981312e-12, 
    -1.985905e-12, -1.972947e-12, -1.980225e-12, -1.975579e-12, 
    -1.971967e-12, -1.998815e-12, -1.985516e-12, -2.012632e-12, 
    -2.004149e-12, -2.025459e-12, -2.011312e-12, -2.028312e-12, 
    -2.025052e-12, -2.034867e-12, -2.032055e-12, -2.044609e-12, 
    -2.036165e-12, -2.051118e-12, -2.042593e-12, -2.043926e-12, 
    -2.035886e-12, -1.988193e-12, -1.997159e-12, -1.987661e-12, -1.98894e-12, 
    -1.988366e-12, -1.981393e-12, -1.977878e-12, -1.970519e-12, 
    -1.971855e-12, -1.97726e-12, -1.989515e-12, -1.985355e-12, -1.99584e-12, 
    -1.995603e-12, -2.007276e-12, -2.002012e-12, -2.021633e-12, 
    -2.016057e-12, -2.032172e-12, -2.028119e-12, -2.031982e-12, 
    -2.030811e-12, -2.031997e-12, -2.026053e-12, -2.0286e-12, -2.023369e-12, 
    -2.002998e-12, -2.008985e-12, -1.99113e-12, -1.980395e-12, -1.973266e-12, 
    -1.968207e-12, -1.968922e-12, -1.970285e-12, -1.977292e-12, -1.98388e-12, 
    -1.988901e-12, -1.992259e-12, -1.995569e-12, -2.005585e-12, 
    -2.010888e-12, -2.022761e-12, -2.020618e-12, -2.024248e-12, 
    -2.027716e-12, -2.033538e-12, -2.03258e-12, -2.035145e-12, -2.024152e-12, 
    -2.031458e-12, -2.019398e-12, -2.022696e-12, -1.996467e-12, 
    -1.986477e-12, -1.98223e-12, -1.978514e-12, -1.969472e-12, -1.975716e-12, 
    -1.973254e-12, -1.979111e-12, -1.982832e-12, -1.980992e-12, 
    -1.992351e-12, -1.987935e-12, -2.011202e-12, -2.00118e-12, -2.027311e-12, 
    -2.021058e-12, -2.02881e-12, -2.024855e-12, -2.031633e-12, -2.025533e-12, 
    -2.0361e-12, -2.038402e-12, -2.036828e-12, -2.04287e-12, -2.025194e-12, 
    -2.031982e-12, -1.98094e-12, -1.98124e-12, -1.982639e-12, -1.976491e-12, 
    -1.976115e-12, -1.970483e-12, -1.975495e-12, -1.977629e-12, 
    -1.983048e-12, -1.986253e-12, -1.9893e-12, -1.996e-12, -2.003482e-12, 
    -2.013945e-12, -2.021463e-12, -2.026503e-12, -2.023413e-12, 
    -2.026141e-12, -2.023091e-12, -2.021662e-12, -2.037539e-12, 
    -2.028623e-12, -2.042001e-12, -2.041261e-12, -2.035206e-12, 
    -2.041344e-12, -1.981451e-12, -1.979724e-12, -1.973727e-12, -1.97842e-12, 
    -1.969869e-12, -1.974655e-12, -1.977407e-12, -1.988027e-12, 
    -1.990361e-12, -1.992524e-12, -1.996797e-12, -2.002282e-12, 
    -2.011903e-12, -2.020275e-12, -2.027918e-12, -2.027358e-12, 
    -2.027555e-12, -2.029262e-12, -2.025033e-12, -2.029956e-12, 
    -2.030783e-12, -2.028622e-12, -2.041162e-12, -2.03758e-12, -2.041245e-12, 
    -2.038913e-12, -1.980286e-12, -1.983192e-12, -1.981621e-12, 
    -1.984575e-12, -1.982494e-12, -1.991746e-12, -1.99452e-12, -2.007501e-12, 
    -2.002174e-12, -2.010653e-12, -2.003035e-12, -2.004385e-12, 
    -2.010929e-12, -2.003447e-12, -2.019813e-12, -2.008717e-12, 
    -2.029329e-12, -2.018246e-12, -2.030023e-12, -2.027885e-12, 
    -2.031425e-12, -2.034596e-12, -2.038586e-12, -2.045947e-12, 
    -2.044242e-12, -2.050398e-12, -1.987525e-12, -1.991295e-12, 
    -1.990963e-12, -1.994909e-12, -1.997827e-12, -2.004152e-12, 
    -2.014296e-12, -2.010481e-12, -2.017485e-12, -2.018891e-12, 
    -2.008251e-12, -2.014783e-12, -1.993818e-12, -1.997205e-12, 
    -1.995189e-12, -1.987822e-12, -2.01136e-12, -1.99928e-12, -2.021588e-12, 
    -2.015043e-12, -2.034144e-12, -2.024644e-12, -2.043304e-12, -2.05128e-12, 
    -2.058789e-12, -2.067563e-12, -1.993353e-12, -1.990791e-12, 
    -1.995378e-12, -2.001724e-12, -2.007613e-12, -2.015442e-12, 
    -2.016243e-12, -2.01771e-12, -2.021509e-12, -2.024704e-12, -2.018173e-12, 
    -2.025505e-12, -1.99799e-12, -2.012409e-12, -1.989822e-12, -1.996623e-12, 
    -2.00135e-12, -1.999277e-12, -2.010045e-12, -2.012583e-12, -2.022897e-12, 
    -2.017566e-12, -2.049311e-12, -2.035265e-12, -2.074244e-12, 
    -2.063351e-12, -1.989896e-12, -1.993344e-12, -2.005344e-12, 
    -1.999635e-12, -2.015965e-12, -2.019985e-12, -2.023253e-12, -2.02743e-12, 
    -2.027881e-12, -2.030356e-12, -2.0263e-12, -2.030196e-12, -2.015459e-12, 
    -2.022044e-12, -2.003973e-12, -2.008371e-12, -2.006348e-12, 
    -2.004128e-12, -2.010978e-12, -2.018276e-12, -2.018433e-12, 
    -2.020772e-12, -2.027366e-12, -2.016031e-12, -2.051123e-12, -2.02945e-12, 
    -1.997104e-12, -2.003745e-12, -2.004694e-12, -2.002122e-12, 
    -2.019582e-12, -2.013255e-12, -2.030296e-12, -2.02569e-12, -2.033237e-12, 
    -2.029487e-12, -2.028935e-12, -2.024119e-12, -2.02112e-12, -2.013545e-12, 
    -2.007382e-12, -2.002495e-12, -2.003631e-12, -2.008999e-12, 
    -2.018723e-12, -2.027922e-12, -2.025907e-12, -2.032663e-12, 
    -2.014781e-12, -2.022279e-12, -2.019381e-12, -2.026938e-12, -2.01038e-12, 
    -2.024478e-12, -2.006776e-12, -2.008328e-12, -2.013129e-12, 
    -2.022787e-12, -2.024924e-12, -2.027206e-12, -2.025798e-12, -2.01897e-12, 
    -2.017851e-12, -2.013013e-12, -2.011677e-12, -2.00799e-12, -2.004938e-12, 
    -2.007727e-12, -2.010655e-12, -2.018973e-12, -2.026468e-12, 
    -2.034641e-12, -2.036641e-12, -2.04619e-12, -2.038417e-12, -2.051244e-12, 
    -2.040338e-12, -2.059218e-12, -2.025296e-12, -2.040018e-12, 
    -2.013348e-12, -2.016221e-12, -2.021417e-12, -2.033337e-12, 
    -2.026902e-12, -2.034428e-12, -2.017807e-12, -2.009184e-12, 
    -2.006954e-12, -2.002792e-12, -2.007049e-12, -2.006703e-12, 
    -2.010777e-12, -2.009467e-12, -2.019249e-12, -2.013995e-12, 
    -2.028921e-12, -2.034368e-12, -2.049753e-12, -2.059184e-12, 
    -2.068786e-12, -2.073025e-12, -2.074315e-12, -2.074855e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.798018e-15, 3.808292e-15, 3.806296e-15, 3.814575e-15, 3.809985e-15, 
    3.815403e-15, 3.800103e-15, 3.808698e-15, 3.803213e-15, 3.798945e-15, 
    3.830615e-15, 3.814944e-15, 3.84688e-15, 3.836903e-15, 3.861948e-15, 
    3.845326e-15, 3.865297e-15, 3.861472e-15, 3.872986e-15, 3.869689e-15, 
    3.884392e-15, 3.874507e-15, 3.89201e-15, 3.882035e-15, 3.883594e-15, 
    3.87418e-15, 3.818103e-15, 3.828665e-15, 3.817476e-15, 3.818983e-15, 
    3.818308e-15, 3.810078e-15, 3.805926e-15, 3.797235e-15, 3.798814e-15, 
    3.805199e-15, 3.819661e-15, 3.814756e-15, 3.827119e-15, 3.82684e-15, 
    3.840582e-15, 3.834389e-15, 3.857459e-15, 3.850909e-15, 3.869827e-15, 
    3.865072e-15, 3.869603e-15, 3.86823e-15, 3.869621e-15, 3.862647e-15, 
    3.865636e-15, 3.859498e-15, 3.835549e-15, 3.842592e-15, 3.821567e-15, 
    3.808897e-15, 3.80048e-15, 3.794501e-15, 3.795346e-15, 3.796957e-15, 
    3.805236e-15, 3.813016e-15, 3.818939e-15, 3.822899e-15, 3.8268e-15, 
    3.838589e-15, 3.844829e-15, 3.858781e-15, 3.856267e-15, 3.860528e-15, 
    3.8646e-15, 3.871428e-15, 3.870304e-15, 3.873311e-15, 3.860417e-15, 
    3.868988e-15, 3.854835e-15, 3.858707e-15, 3.827849e-15, 3.81608e-15, 
    3.811064e-15, 3.80668e-15, 3.795996e-15, 3.803374e-15, 3.800466e-15, 
    3.807386e-15, 3.811779e-15, 3.809607e-15, 3.823007e-15, 3.817799e-15, 
    3.845199e-15, 3.833407e-15, 3.864125e-15, 3.856784e-15, 3.865884e-15, 
    3.861242e-15, 3.869193e-15, 3.862037e-15, 3.87443e-15, 3.877126e-15, 
    3.875284e-15, 3.88236e-15, 3.861641e-15, 3.869602e-15, 3.809546e-15, 
    3.8099e-15, 3.811551e-15, 3.80429e-15, 3.803847e-15, 3.797191e-15, 
    3.803114e-15, 3.805635e-15, 3.812034e-15, 3.815816e-15, 3.819409e-15, 
    3.827307e-15, 3.836117e-15, 3.848425e-15, 3.85726e-15, 3.863177e-15, 
    3.859549e-15, 3.862751e-15, 3.859171e-15, 3.857493e-15, 3.876115e-15, 
    3.865663e-15, 3.881343e-15, 3.880476e-15, 3.873382e-15, 3.880574e-15, 
    3.810149e-15, 3.80811e-15, 3.801025e-15, 3.80657e-15, 3.796466e-15, 
    3.802122e-15, 3.805371e-15, 3.817906e-15, 3.82066e-15, 3.82321e-15, 
    3.828247e-15, 3.834706e-15, 3.846024e-15, 3.855863e-15, 3.864837e-15, 
    3.86418e-15, 3.864411e-15, 3.866414e-15, 3.861451e-15, 3.867228e-15, 
    3.868196e-15, 3.865663e-15, 3.88036e-15, 3.876164e-15, 3.880458e-15, 
    3.877726e-15, 3.808773e-15, 3.812203e-15, 3.81035e-15, 3.813834e-15, 
    3.811378e-15, 3.822291e-15, 3.82556e-15, 3.840845e-15, 3.834578e-15, 
    3.844554e-15, 3.835593e-15, 3.837181e-15, 3.844874e-15, 3.836078e-15, 
    3.855319e-15, 3.842274e-15, 3.866491e-15, 3.853476e-15, 3.867306e-15, 
    3.864798e-15, 3.868951e-15, 3.872668e-15, 3.877343e-15, 3.885961e-15, 
    3.883966e-15, 3.89117e-15, 3.817316e-15, 3.821761e-15, 3.821371e-15, 
    3.826022e-15, 3.829459e-15, 3.836907e-15, 3.848839e-15, 3.844354e-15, 
    3.852587e-15, 3.854238e-15, 3.841731e-15, 3.84941e-15, 3.824735e-15, 
    3.828724e-15, 3.826351e-15, 3.817666e-15, 3.845385e-15, 3.831169e-15, 
    3.857405e-15, 3.849717e-15, 3.872137e-15, 3.860992e-15, 3.882868e-15, 
    3.892198e-15, 3.900978e-15, 3.911217e-15, 3.824187e-15, 3.821168e-15, 
    3.826575e-15, 3.834047e-15, 3.84098e-15, 3.850186e-15, 3.851128e-15, 
    3.852851e-15, 3.857314e-15, 3.861065e-15, 3.853393e-15, 3.862005e-15, 
    3.829645e-15, 3.846619e-15, 3.820025e-15, 3.828038e-15, 3.833608e-15, 
    3.831167e-15, 3.843842e-15, 3.846826e-15, 3.858942e-15, 3.852682e-15, 
    3.889894e-15, 3.873449e-15, 3.919012e-15, 3.906302e-15, 3.820113e-15, 
    3.824178e-15, 3.838309e-15, 3.831589e-15, 3.850801e-15, 3.855523e-15, 
    3.859362e-15, 3.864263e-15, 3.864794e-15, 3.867696e-15, 3.862939e-15, 
    3.867509e-15, 3.850205e-15, 3.857942e-15, 3.836698e-15, 3.841872e-15, 
    3.839492e-15, 3.836881e-15, 3.844939e-15, 3.853514e-15, 3.8537e-15, 
    3.856447e-15, 3.864179e-15, 3.850879e-15, 3.892008e-15, 3.866625e-15, 
    3.828608e-15, 3.836425e-15, 3.837545e-15, 3.834518e-15, 3.855049e-15, 
    3.847615e-15, 3.867626e-15, 3.862223e-15, 3.871075e-15, 3.866677e-15, 
    3.866029e-15, 3.860378e-15, 3.856857e-15, 3.847955e-15, 3.840707e-15, 
    3.834957e-15, 3.836295e-15, 3.84261e-15, 3.854039e-15, 3.86484e-15, 
    3.862475e-15, 3.870403e-15, 3.849409e-15, 3.858216e-15, 3.854812e-15, 
    3.863686e-15, 3.844234e-15, 3.860791e-15, 3.839996e-15, 3.841822e-15, 
    3.847467e-15, 3.858811e-15, 3.861324e-15, 3.864e-15, 3.86235e-15, 
    3.854329e-15, 3.853017e-15, 3.847331e-15, 3.845759e-15, 3.841425e-15, 
    3.837833e-15, 3.841114e-15, 3.844557e-15, 3.854334e-15, 3.863134e-15, 
    3.87272e-15, 3.875066e-15, 3.886241e-15, 3.87714e-15, 3.892149e-15, 
    3.879384e-15, 3.901472e-15, 3.861755e-15, 3.879014e-15, 3.847725e-15, 
    3.851102e-15, 3.857203e-15, 3.871188e-15, 3.863645e-15, 3.872468e-15, 
    3.852965e-15, 3.842826e-15, 3.840205e-15, 3.835306e-15, 3.840317e-15, 
    3.83991e-15, 3.844702e-15, 3.843163e-15, 3.854658e-15, 3.848485e-15, 
    3.866013e-15, 3.872399e-15, 3.890414e-15, 3.901437e-15, 3.912648e-15, 
    3.917591e-15, 3.919096e-15, 3.919724e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.562789e-09, -8.600542e-09, -8.593203e-09, -8.623654e-09, -8.606762e-09, 
    -8.626701e-09, -8.570444e-09, -8.60204e-09, -8.58187e-09, -8.566189e-09, 
    -8.682747e-09, -8.625013e-09, -8.742733e-09, -8.705906e-09, 
    -8.798422e-09, -8.737001e-09, -8.810808e-09, -8.796652e-09, 
    -8.839263e-09, -8.827056e-09, -8.881558e-09, -8.844897e-09, 
    -8.909813e-09, -8.872805e-09, -8.878593e-09, -8.843688e-09, 
    -8.636633e-09, -8.675559e-09, -8.634326e-09, -8.639876e-09, 
    -8.637387e-09, -8.607111e-09, -8.591853e-09, -8.559905e-09, 
    -8.565705e-09, -8.589171e-09, -8.642373e-09, -8.624314e-09, 
    -8.669831e-09, -8.668803e-09, -8.719479e-09, -8.69663e-09, -8.781811e-09, 
    -8.757601e-09, -8.827565e-09, -8.809969e-09, -8.826738e-09, 
    -8.821654e-09, -8.826804e-09, -8.800998e-09, -8.812054e-09, 
    -8.789347e-09, -8.700908e-09, -8.726898e-09, -8.649386e-09, -8.60278e-09, 
    -8.571829e-09, -8.549866e-09, -8.552971e-09, -8.55889e-09, -8.589308e-09, 
    -8.617911e-09, -8.639708e-09, -8.654289e-09, -8.668656e-09, -8.71214e-09, 
    -8.735161e-09, -8.786706e-09, -8.777405e-09, -8.793163e-09, 
    -8.808219e-09, -8.833495e-09, -8.829335e-09, -8.840471e-09, 
    -8.792748e-09, -8.824464e-09, -8.772107e-09, -8.786427e-09, 
    -8.672555e-09, -8.629186e-09, -8.610748e-09, -8.594614e-09, 
    -8.555358e-09, -8.582466e-09, -8.57178e-09, -8.597206e-09, -8.613362e-09, 
    -8.605372e-09, -8.654688e-09, -8.635514e-09, -8.736525e-09, 
    -8.693015e-09, -8.806462e-09, -8.779314e-09, -8.81297e-09, -8.795796e-09, 
    -8.825222e-09, -8.79874e-09, -8.844616e-09, -8.854608e-09, -8.847779e-09, 
    -8.874006e-09, -8.797271e-09, -8.826738e-09, -8.605147e-09, -8.60645e-09, 
    -8.612521e-09, -8.585832e-09, -8.5842e-09, -8.559746e-09, -8.581506e-09, 
    -8.590773e-09, -8.614299e-09, -8.628213e-09, -8.641441e-09, 
    -8.670526e-09, -8.703009e-09, -8.748435e-09, -8.781074e-09, 
    -8.802952e-09, -8.789537e-09, -8.801381e-09, -8.788141e-09, 
    -8.781935e-09, -8.850865e-09, -8.812157e-09, -8.870234e-09, 
    -8.867022e-09, -8.840735e-09, -8.867383e-09, -8.607365e-09, 
    -8.599867e-09, -8.57383e-09, -8.594205e-09, -8.557082e-09, -8.577861e-09, 
    -8.589809e-09, -8.635913e-09, -8.646045e-09, -8.655437e-09, -8.67399e-09, 
    -8.6978e-09, -8.739568e-09, -8.775913e-09, -8.809095e-09, -8.806664e-09, 
    -8.80752e-09, -8.814932e-09, -8.796571e-09, -8.817945e-09, -8.821533e-09, 
    -8.812154e-09, -8.866591e-09, -8.851039e-09, -8.866953e-09, 
    -8.856827e-09, -8.602304e-09, -8.614922e-09, -8.608104e-09, 
    -8.620925e-09, -8.611892e-09, -8.652059e-09, -8.664101e-09, 
    -8.720458e-09, -8.697331e-09, -8.734141e-09, -8.70107e-09, -8.706929e-09, 
    -8.735339e-09, -8.702858e-09, -8.773908e-09, -8.725735e-09, -8.81522e-09, 
    -8.767109e-09, -8.818234e-09, -8.808952e-09, -8.824322e-09, 
    -8.838088e-09, -8.85541e-09, -8.887365e-09, -8.879965e-09, -8.906691e-09, 
    -8.633735e-09, -8.650101e-09, -8.648661e-09, -8.66579e-09, -8.678458e-09, 
    -8.705917e-09, -8.749957e-09, -8.733396e-09, -8.763802e-09, 
    -8.769906e-09, -8.723713e-09, -8.752073e-09, -8.661056e-09, 
    -8.675759e-09, -8.667005e-09, -8.635025e-09, -8.737211e-09, 
    -8.684767e-09, -8.781613e-09, -8.7532e-09, -8.836125e-09, -8.794883e-09, 
    -8.875892e-09, -8.91052e-09, -8.943118e-09, -8.981207e-09, -8.659034e-09, 
    -8.647913e-09, -8.667827e-09, -8.695378e-09, -8.720944e-09, 
    -8.754933e-09, -8.758412e-09, -8.764778e-09, -8.781273e-09, 
    -8.795142e-09, -8.766791e-09, -8.798619e-09, -8.679167e-09, 
    -8.741764e-09, -8.643708e-09, -8.673232e-09, -8.693754e-09, 
    -8.684752e-09, -8.731504e-09, -8.742522e-09, -8.7873e-09, -8.764153e-09, 
    -8.901972e-09, -8.840994e-09, -9.010214e-09, -8.962921e-09, 
    -8.644028e-09, -8.658997e-09, -8.711095e-09, -8.686307e-09, 
    -8.757203e-09, -8.774654e-09, -8.788843e-09, -8.806977e-09, 
    -8.808936e-09, -8.819681e-09, -8.802073e-09, -8.818986e-09, 
    -8.755006e-09, -8.783597e-09, -8.705141e-09, -8.724236e-09, 
    -8.715451e-09, -8.705817e-09, -8.735555e-09, -8.767237e-09, 
    -8.767915e-09, -8.778074e-09, -8.806698e-09, -8.75749e-09, -8.909838e-09, 
    -8.815745e-09, -8.67532e-09, -8.704152e-09, -8.708272e-09, -8.697103e-09, 
    -8.772904e-09, -8.745438e-09, -8.81942e-09, -8.799425e-09, -8.832187e-09, 
    -8.815906e-09, -8.813511e-09, -8.792602e-09, -8.779584e-09, 
    -8.746697e-09, -8.719939e-09, -8.698724e-09, -8.703656e-09, 
    -8.726962e-09, -8.769176e-09, -8.809113e-09, -8.800364e-09, 
    -8.829697e-09, -8.752062e-09, -8.784614e-09, -8.772032e-09, -8.80484e-09, 
    -8.732956e-09, -8.794163e-09, -8.717311e-09, -8.724049e-09, 
    -8.744893e-09, -8.78682e-09, -8.7961e-09, -8.806004e-09, -8.799893e-09, 
    -8.770248e-09, -8.765391e-09, -8.744387e-09, -8.738586e-09, 
    -8.722583e-09, -8.709332e-09, -8.721438e-09, -8.734151e-09, -8.77026e-09, 
    -8.802802e-09, -8.838283e-09, -8.846968e-09, -8.888422e-09, 
    -8.854676e-09, -8.910362e-09, -8.863014e-09, -8.944981e-09, 
    -8.797713e-09, -8.861625e-09, -8.745842e-09, -8.758315e-09, 
    -8.780874e-09, -8.83262e-09, -8.804686e-09, -8.837356e-09, -8.765201e-09, 
    -8.727766e-09, -8.718082e-09, -8.700013e-09, -8.718496e-09, 
    -8.716992e-09, -8.734679e-09, -8.728995e-09, -8.771459e-09, -8.74865e-09, 
    -8.81345e-09, -8.837098e-09, -8.903889e-09, -8.944833e-09, -8.986517e-09, 
    -9.004919e-09, -9.010521e-09, -9.012862e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.016115e-10, -1.020597e-10, -1.019726e-10, -1.023341e-10, -1.021336e-10, 
    -1.023702e-10, -1.017024e-10, -1.020775e-10, -1.018381e-10, 
    -1.016519e-10, -1.030356e-10, -1.023502e-10, -1.037477e-10, 
    -1.033105e-10, -1.044088e-10, -1.036796e-10, -1.045558e-10, 
    -1.043878e-10, -1.048937e-10, -1.047487e-10, -1.053958e-10, 
    -1.049605e-10, -1.057312e-10, -1.052919e-10, -1.053606e-10, 
    -1.049462e-10, -1.024881e-10, -1.029502e-10, -1.024608e-10, 
    -1.025267e-10, -1.024971e-10, -1.021377e-10, -1.019566e-10, 
    -1.015773e-10, -1.016462e-10, -1.019247e-10, -1.025563e-10, 
    -1.023419e-10, -1.028822e-10, -1.0287e-10, -1.034716e-10, -1.032004e-10, 
    -1.042116e-10, -1.039242e-10, -1.047548e-10, -1.045459e-10, -1.04745e-10, 
    -1.046846e-10, -1.047458e-10, -1.044394e-10, -1.045706e-10, 
    -1.043011e-10, -1.032512e-10, -1.035597e-10, -1.026395e-10, 
    -1.020863e-10, -1.017189e-10, -1.014581e-10, -1.01495e-10, -1.015652e-10, 
    -1.019263e-10, -1.022659e-10, -1.025246e-10, -1.026977e-10, 
    -1.028683e-10, -1.033845e-10, -1.036578e-10, -1.042697e-10, 
    -1.041593e-10, -1.043464e-10, -1.045251e-10, -1.048252e-10, 
    -1.047758e-10, -1.04908e-10, -1.043414e-10, -1.04718e-10, -1.040964e-10, 
    -1.042664e-10, -1.029146e-10, -1.023997e-10, -1.021809e-10, 
    -1.019893e-10, -1.015233e-10, -1.018451e-10, -1.017183e-10, 
    -1.020201e-10, -1.022119e-10, -1.02117e-10, -1.027025e-10, -1.024749e-10, 
    -1.03674e-10, -1.031575e-10, -1.045043e-10, -1.04182e-10, -1.045815e-10, 
    -1.043776e-10, -1.04727e-10, -1.044126e-10, -1.049572e-10, -1.050758e-10, 
    -1.049948e-10, -1.053061e-10, -1.043951e-10, -1.04745e-10, -1.021144e-10, 
    -1.021298e-10, -1.022019e-10, -1.018851e-10, -1.018657e-10, 
    -1.015754e-10, -1.018337e-10, -1.019437e-10, -1.02223e-10, -1.023882e-10, 
    -1.025452e-10, -1.028905e-10, -1.032761e-10, -1.038154e-10, 
    -1.042028e-10, -1.044626e-10, -1.043033e-10, -1.044439e-10, 
    -1.042867e-10, -1.042131e-10, -1.050314e-10, -1.045719e-10, 
    -1.052613e-10, -1.052232e-10, -1.049111e-10, -1.052275e-10, 
    -1.021407e-10, -1.020517e-10, -1.017426e-10, -1.019845e-10, 
    -1.015438e-10, -1.017905e-10, -1.019323e-10, -1.024796e-10, 
    -1.025999e-10, -1.027114e-10, -1.029316e-10, -1.032143e-10, 
    -1.037101e-10, -1.041416e-10, -1.045355e-10, -1.045066e-10, 
    -1.045168e-10, -1.046048e-10, -1.043868e-10, -1.046406e-10, 
    -1.046832e-10, -1.045718e-10, -1.052181e-10, -1.050335e-10, 
    -1.052224e-10, -1.051022e-10, -1.020806e-10, -1.022304e-10, 
    -1.021495e-10, -1.023017e-10, -1.021944e-10, -1.026713e-10, 
    -1.028142e-10, -1.034832e-10, -1.032087e-10, -1.036457e-10, 
    -1.032531e-10, -1.033226e-10, -1.036599e-10, -1.032743e-10, 
    -1.041178e-10, -1.035459e-10, -1.046082e-10, -1.040371e-10, -1.04644e-10, 
    -1.045338e-10, -1.047163e-10, -1.048797e-10, -1.050854e-10, 
    -1.054647e-10, -1.053769e-10, -1.056942e-10, -1.024537e-10, -1.02648e-10, 
    -1.026309e-10, -1.028343e-10, -1.029846e-10, -1.033106e-10, 
    -1.038334e-10, -1.036368e-10, -1.039978e-10, -1.040703e-10, 
    -1.035219e-10, -1.038586e-10, -1.027781e-10, -1.029526e-10, 
    -1.028487e-10, -1.024691e-10, -1.036821e-10, -1.030595e-10, 
    -1.042093e-10, -1.038719e-10, -1.048564e-10, -1.043668e-10, 
    -1.053285e-10, -1.057396e-10, -1.061266e-10, -1.065788e-10, 
    -1.027541e-10, -1.026221e-10, -1.028585e-10, -1.031855e-10, -1.03489e-10, 
    -1.038925e-10, -1.039338e-10, -1.040094e-10, -1.042052e-10, 
    -1.043699e-10, -1.040333e-10, -1.044111e-10, -1.029931e-10, 
    -1.037362e-10, -1.025721e-10, -1.029226e-10, -1.031662e-10, 
    -1.030594e-10, -1.036144e-10, -1.037452e-10, -1.042768e-10, -1.04002e-10, 
    -1.056381e-10, -1.049142e-10, -1.069232e-10, -1.063617e-10, 
    -1.025759e-10, -1.027536e-10, -1.033721e-10, -1.030778e-10, 
    -1.039195e-10, -1.041266e-10, -1.042951e-10, -1.045104e-10, 
    -1.045336e-10, -1.046612e-10, -1.044521e-10, -1.046529e-10, 
    -1.038934e-10, -1.042328e-10, -1.033014e-10, -1.035281e-10, 
    -1.034238e-10, -1.033094e-10, -1.036625e-10, -1.040386e-10, 
    -1.040466e-10, -1.041672e-10, -1.045071e-10, -1.039229e-10, 
    -1.057315e-10, -1.046145e-10, -1.029474e-10, -1.032897e-10, 
    -1.033386e-10, -1.03206e-10, -1.041059e-10, -1.037798e-10, -1.046581e-10, 
    -1.044207e-10, -1.048096e-10, -1.046164e-10, -1.045879e-10, 
    -1.043397e-10, -1.041852e-10, -1.037947e-10, -1.034771e-10, 
    -1.032252e-10, -1.032838e-10, -1.035605e-10, -1.040616e-10, 
    -1.045357e-10, -1.044319e-10, -1.047801e-10, -1.038584e-10, 
    -1.042449e-10, -1.040955e-10, -1.04485e-10, -1.036316e-10, -1.043582e-10, 
    -1.034459e-10, -1.035259e-10, -1.037733e-10, -1.042711e-10, 
    -1.043812e-10, -1.044988e-10, -1.044263e-10, -1.040743e-10, 
    -1.040167e-10, -1.037673e-10, -1.036985e-10, -1.035085e-10, 
    -1.033512e-10, -1.034949e-10, -1.036458e-10, -1.040745e-10, 
    -1.044608e-10, -1.04882e-10, -1.049851e-10, -1.054773e-10, -1.050766e-10, 
    -1.057377e-10, -1.051756e-10, -1.061487e-10, -1.044004e-10, 
    -1.051591e-10, -1.037846e-10, -1.039327e-10, -1.042005e-10, 
    -1.048148e-10, -1.044832e-10, -1.04871e-10, -1.040144e-10, -1.0357e-10, 
    -1.034551e-10, -1.032405e-10, -1.0346e-10, -1.034421e-10, -1.036521e-10, 
    -1.035846e-10, -1.040887e-10, -1.038179e-10, -1.045872e-10, -1.04868e-10, 
    -1.056609e-10, -1.06147e-10, -1.066419e-10, -1.068604e-10, -1.069268e-10, 
    -1.069547e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.427539e-12, -8.464725e-12, -8.457497e-12, -8.48749e-12, -8.470853e-12, 
    -8.490492e-12, -8.435079e-12, -8.466201e-12, -8.446334e-12, 
    -8.430888e-12, -8.545698e-12, -8.488829e-12, -8.604784e-12, -8.56851e-12, 
    -8.659639e-12, -8.599139e-12, -8.671839e-12, -8.657896e-12, 
    -8.699868e-12, -8.687844e-12, -8.74153e-12, -8.705418e-12, -8.769363e-12, 
    -8.732908e-12, -8.73861e-12, -8.704227e-12, -8.500275e-12, -8.538617e-12, 
    -8.498003e-12, -8.50347e-12, -8.501018e-12, -8.471196e-12, -8.456167e-12, 
    -8.424698e-12, -8.430412e-12, -8.453525e-12, -8.505929e-12, 
    -8.488141e-12, -8.532976e-12, -8.531963e-12, -8.581879e-12, 
    -8.559373e-12, -8.643277e-12, -8.61943e-12, -8.688346e-12, -8.671014e-12, 
    -8.687532e-12, -8.682523e-12, -8.687597e-12, -8.662177e-12, 
    -8.673067e-12, -8.650701e-12, -8.563587e-12, -8.589188e-12, 
    -8.512837e-12, -8.466929e-12, -8.436443e-12, -8.41481e-12, -8.417868e-12, 
    -8.423698e-12, -8.453661e-12, -8.481833e-12, -8.503304e-12, 
    -8.517666e-12, -8.531818e-12, -8.57465e-12, -8.597326e-12, -8.648098e-12, 
    -8.638937e-12, -8.654458e-12, -8.669289e-12, -8.694187e-12, 
    -8.690089e-12, -8.701058e-12, -8.65405e-12, -8.685291e-12, -8.633718e-12, 
    -8.647823e-12, -8.535658e-12, -8.49294e-12, -8.474778e-12, -8.458886e-12, 
    -8.420219e-12, -8.446921e-12, -8.436395e-12, -8.461439e-12, 
    -8.477353e-12, -8.469482e-12, -8.518059e-12, -8.499173e-12, -8.59867e-12, 
    -8.555811e-12, -8.667559e-12, -8.640817e-12, -8.67397e-12, -8.657053e-12, 
    -8.686038e-12, -8.659952e-12, -8.705142e-12, -8.714984e-12, 
    -8.708257e-12, -8.734092e-12, -8.658505e-12, -8.687531e-12, 
    -8.469262e-12, -8.470545e-12, -8.476525e-12, -8.450237e-12, 
    -8.448629e-12, -8.424541e-12, -8.445976e-12, -8.455103e-12, 
    -8.478275e-12, -8.491981e-12, -8.505011e-12, -8.53366e-12, -8.565656e-12, 
    -8.610401e-12, -8.642551e-12, -8.664102e-12, -8.650887e-12, 
    -8.662553e-12, -8.649512e-12, -8.643399e-12, -8.711296e-12, 
    -8.673169e-12, -8.730377e-12, -8.727212e-12, -8.701319e-12, 
    -8.727568e-12, -8.471447e-12, -8.46406e-12, -8.438414e-12, -8.458484e-12, 
    -8.421919e-12, -8.442385e-12, -8.454153e-12, -8.499567e-12, 
    -8.509545e-12, -8.518798e-12, -8.537072e-12, -8.560525e-12, 
    -8.601667e-12, -8.637467e-12, -8.670152e-12, -8.667757e-12, 
    -8.668601e-12, -8.675901e-12, -8.657816e-12, -8.678871e-12, 
    -8.682404e-12, -8.673165e-12, -8.726788e-12, -8.711469e-12, 
    -8.727144e-12, -8.71717e-12, -8.466461e-12, -8.47889e-12, -8.472174e-12, 
    -8.484803e-12, -8.475906e-12, -8.51547e-12, -8.527332e-12, -8.582844e-12, 
    -8.560062e-12, -8.596321e-12, -8.563746e-12, -8.569517e-12, 
    -8.597501e-12, -8.565507e-12, -8.635492e-12, -8.588042e-12, 
    -8.676185e-12, -8.628795e-12, -8.679155e-12, -8.670011e-12, 
    -8.685152e-12, -8.698711e-12, -8.715774e-12, -8.74725e-12, -8.739962e-12, 
    -8.766287e-12, -8.49742e-12, -8.513541e-12, -8.512123e-12, -8.528995e-12, 
    -8.541473e-12, -8.56852e-12, -8.611901e-12, -8.595588e-12, -8.625538e-12, 
    -8.631549e-12, -8.586049e-12, -8.613985e-12, -8.524331e-12, 
    -8.538814e-12, -8.530192e-12, -8.498691e-12, -8.599345e-12, 
    -8.547687e-12, -8.643082e-12, -8.615095e-12, -8.696777e-12, 
    -8.656153e-12, -8.735949e-12, -8.770058e-12, -8.802169e-12, 
    -8.839689e-12, -8.522341e-12, -8.511387e-12, -8.531001e-12, 
    -8.558139e-12, -8.583322e-12, -8.616802e-12, -8.620228e-12, -8.6265e-12, 
    -8.642748e-12, -8.656408e-12, -8.628482e-12, -8.659832e-12, -8.54217e-12, 
    -8.603829e-12, -8.507244e-12, -8.536325e-12, -8.55654e-12, -8.547673e-12, 
    -8.593724e-12, -8.604577e-12, -8.648683e-12, -8.625884e-12, 
    -8.761639e-12, -8.701573e-12, -8.868261e-12, -8.821675e-12, 
    -8.507559e-12, -8.522304e-12, -8.573621e-12, -8.549204e-12, 
    -8.619038e-12, -8.636227e-12, -8.650203e-12, -8.668066e-12, 
    -8.669995e-12, -8.68058e-12, -8.663236e-12, -8.679895e-12, -8.616873e-12, 
    -8.645036e-12, -8.567757e-12, -8.586565e-12, -8.577913e-12, 
    -8.568421e-12, -8.597714e-12, -8.628921e-12, -8.62959e-12, -8.639597e-12, 
    -8.667791e-12, -8.619321e-12, -8.769388e-12, -8.676703e-12, 
    -8.538383e-12, -8.566782e-12, -8.57084e-12, -8.559839e-12, -8.634504e-12, 
    -8.607449e-12, -8.680322e-12, -8.660627e-12, -8.692898e-12, 
    -8.676861e-12, -8.674502e-12, -8.653907e-12, -8.641084e-12, 
    -8.608689e-12, -8.582333e-12, -8.561435e-12, -8.566294e-12, 
    -8.589251e-12, -8.63083e-12, -8.67017e-12, -8.661552e-12, -8.690445e-12, 
    -8.613974e-12, -8.646038e-12, -8.633644e-12, -8.665961e-12, 
    -8.595154e-12, -8.655444e-12, -8.579744e-12, -8.586381e-12, 
    -8.606912e-12, -8.648211e-12, -8.657352e-12, -8.667108e-12, 
    -8.661088e-12, -8.631887e-12, -8.627103e-12, -8.606413e-12, -8.6007e-12, 
    -8.584936e-12, -8.571885e-12, -8.583808e-12, -8.596331e-12, -8.6319e-12, 
    -8.663954e-12, -8.698904e-12, -8.707457e-12, -8.748292e-12, -8.71505e-12, 
    -8.769903e-12, -8.723264e-12, -8.804004e-12, -8.658941e-12, 
    -8.721896e-12, -8.607847e-12, -8.620133e-12, -8.642354e-12, 
    -8.693325e-12, -8.665809e-12, -8.697989e-12, -8.626916e-12, 
    -8.590042e-12, -8.580503e-12, -8.562705e-12, -8.58091e-12, -8.57943e-12, 
    -8.596852e-12, -8.591253e-12, -8.63308e-12, -8.610612e-12, -8.674442e-12, 
    -8.697736e-12, -8.763527e-12, -8.803859e-12, -8.84492e-12, -8.863047e-12, 
    -8.868564e-12, -8.87087e-12 ;

 SMIN_NH4 =
  0.0004368965, 0.0004387366, 0.0004383788, 0.0004398629, 0.0004390396, 
    0.0004400112, 0.0004372693, 0.0004388092, 0.0004378261, 0.0004370617, 
    0.0004427424, 0.0004399286, 0.0004456654, 0.0004438708, 0.0004483787, 
    0.0004453859, 0.0004489821, 0.0004482923, 0.0004503683, 0.0004497735, 
    0.0004524288, 0.0004506427, 0.0004538051, 0.0004520022, 0.0004522842, 
    0.0004505835, 0.0004404954, 0.0004423925, 0.0004403828, 0.0004406534, 
    0.0004405319, 0.0004390563, 0.0004383127, 0.0004367554, 0.000437038, 
    0.0004381818, 0.0004407746, 0.0004398944, 0.0004421126, 0.0004420625, 
    0.0004445319, 0.0004434185, 0.0004475691, 0.0004463893, 0.0004497982, 
    0.0004489409, 0.0004497579, 0.0004495101, 0.0004497609, 0.0004485036, 
    0.0004490422, 0.0004479358, 0.0004436277, 0.000444894, 0.0004411167, 
    0.0004388452, 0.0004373366, 0.0004362661, 0.0004364173, 0.0004367058, 
    0.0004381884, 0.0004395823, 0.0004406446, 0.0004413551, 0.0004420552, 
    0.0004441743, 0.000445296, 0.0004478075, 0.0004473543, 0.000448122, 
    0.0004488555, 0.0004500869, 0.0004498842, 0.0004504267, 0.0004481015, 
    0.0004496468, 0.0004470956, 0.0004477934, 0.0004422458, 0.0004401321, 
    0.0004392335, 0.000438447, 0.0004365336, 0.0004378549, 0.000437334, 
    0.0004385732, 0.0004393605, 0.000438971, 0.0004413745, 0.00044044, 
    0.0004453624, 0.0004432421, 0.00044877, 0.0004474472, 0.0004490869, 
    0.0004482502, 0.0004496838, 0.0004483935, 0.0004506285, 0.0004511154, 
    0.0004507825, 0.0004520603, 0.0004483216, 0.0004497573, 0.0004389604, 
    0.0004390239, 0.0004393198, 0.0004380189, 0.0004379393, 0.0004367473, 
    0.0004378078, 0.0004382595, 0.000439406, 0.0004400841, 0.0004407287, 
    0.0004421461, 0.000443729, 0.0004459425, 0.0004475329, 0.0004485988, 
    0.0004479451, 0.0004485221, 0.000447877, 0.0004475745, 0.0004509329, 
    0.000449047, 0.0004518764, 0.0004517199, 0.0004504392, 0.0004517374, 
    0.0004390684, 0.0004387028, 0.0004374338, 0.0004384269, 0.0004366174, 
    0.0004376302, 0.0004382124, 0.0004404593, 0.000440953, 0.0004414108, 
    0.0004423149, 0.0004434751, 0.0004455104, 0.0004472813, 0.000448898, 
    0.0004487794, 0.0004488211, 0.0004491822, 0.0004482876, 0.0004493289, 
    0.0004495036, 0.0004490467, 0.0004516988, 0.0004509412, 0.0004517164, 
    0.000451223, 0.0004388216, 0.0004394365, 0.0004391041, 0.000439729, 
    0.0004392886, 0.0004412462, 0.000441833, 0.0004445793, 0.0004434522, 
    0.000445246, 0.0004436343, 0.0004439199, 0.0004453042, 0.0004437213, 
    0.0004471834, 0.000444836, 0.0004491961, 0.0004468519, 0.0004493429, 
    0.0004488906, 0.0004496393, 0.00045031, 0.0004511539, 0.0004527107, 
    0.0004523501, 0.0004536521, 0.0004403533, 0.0004411508, 0.0004410806, 
    0.0004419153, 0.0004425326, 0.0004438707, 0.0004460167, 0.0004452096, 
    0.0004466911, 0.0004469885, 0.0004447376, 0.0004461195, 0.0004416841, 
    0.0004424006, 0.000441974, 0.0004404153, 0.000445395, 0.0004428393, 
    0.0004475585, 0.0004461739, 0.0004502143, 0.0004482049, 0.0004521516, 
    0.0004538386, 0.0004554264, 0.0004572816, 0.0004415861, 0.0004410441, 
    0.0004420145, 0.0004433571, 0.0004446028, 0.000446259, 0.0004464285, 
    0.0004467386, 0.0004475423, 0.000448218, 0.0004468366, 0.0004483872, 
    0.0004425666, 0.0004456169, 0.0004408384, 0.0004422772, 0.0004432772, 
    0.0004428386, 0.0004451167, 0.0004456535, 0.0004478352, 0.0004467074, 
    0.000453422, 0.0004504512, 0.0004586944, 0.0004563908, 0.0004408546, 
    0.0004415841, 0.0004441229, 0.0004429149, 0.0004463695, 0.0004472198, 
    0.000447911, 0.0004487946, 0.0004488899, 0.0004494135, 0.0004485555, 
    0.0004493795, 0.000446262, 0.0004476551, 0.0004438321, 0.0004447625, 
    0.0004443344, 0.0004438648, 0.0004453139, 0.0004468577, 0.0004468907, 
    0.0004473856, 0.0004487803, 0.0004463825, 0.0004538051, 0.0004492209, 
    0.0004423795, 0.0004437844, 0.0004439852, 0.0004434409, 0.0004471344, 
    0.0004457961, 0.0004494007, 0.0004484264, 0.0004500226, 0.0004492294, 
    0.0004491126, 0.0004480939, 0.0004474595, 0.000445857, 0.000444553, 
    0.0004435192, 0.0004437595, 0.0004448952, 0.000446952, 0.0004488979, 
    0.0004484715, 0.0004499006, 0.0004461179, 0.000447704, 0.0004470908, 
    0.0004486894, 0.0004451879, 0.0004481704, 0.0004444255, 0.0004447538, 
    0.0004457694, 0.0004478123, 0.0004482643, 0.0004487469, 0.000448449, 
    0.0004470046, 0.0004467679, 0.0004457443, 0.0004454616, 0.0004446818, 
    0.000444036, 0.0004446259, 0.0004452453, 0.0004470048, 0.0004485903, 
    0.0004503189, 0.000450742, 0.0004527616, 0.0004511175, 0.0004538303, 
    0.0004515237, 0.0004555165, 0.0004483431, 0.0004514571, 0.0004458156, 
    0.0004464233, 0.0004475225, 0.0004500436, 0.0004486825, 0.0004502743, 
    0.0004467586, 0.0004449344, 0.0004444625, 0.000443582, 0.0004444825, 
    0.0004444093, 0.000445271, 0.000444994, 0.0004470631, 0.0004459516, 
    0.0004491089, 0.0004502611, 0.0004535149, 0.0004555094, 0.0004575397, 
    0.000458436, 0.0004587088, 0.0004588228 ;

 SMIN_NH4_vr =
  0.002871801, 0.002876779, 0.002875805, 0.002879816, 0.002877589, 
    0.002880208, 0.002872796, 0.002876954, 0.002874296, 0.002872224, 
    0.00288756, 0.00287997, 0.002895438, 0.0028906, 0.00290273, 0.002894677, 
    0.00290435, 0.002902492, 0.00290807, 0.002906468, 0.002913589, 
    0.002908799, 0.002917274, 0.002912442, 0.002913193, 0.002908625, 
    0.002881523, 0.002886638, 0.002881213, 0.002881943, 0.002881612, 
    0.002877621, 0.002875607, 0.002871393, 0.002872154, 0.002875247, 
    0.002882249, 0.002879868, 0.002885854, 0.00288572, 0.00289237, 
    0.00288937, 0.002900544, 0.002897365, 0.002906531, 0.002904222, 
    0.002906416, 0.002905746, 0.002906416, 0.002903037, 0.002904478, 
    0.002901505, 0.002889969, 0.002893377, 0.002883189, 0.002877045, 
    0.002872965, 0.002870069, 0.002870472, 0.002871253, 0.002875259, 
    0.002879023, 0.002881892, 0.002883805, 0.002885691, 0.002891402, 
    0.002894422, 0.002901177, 0.002899959, 0.002902017, 0.00290399, 
    0.002907293, 0.002906748, 0.0029082, 0.002901948, 0.002906101, 
    0.002899237, 0.002901114, 0.002886228, 0.002880524, 0.002878092, 
    0.002875964, 0.002870784, 0.002874359, 0.002872946, 0.002876294, 
    0.002878421, 0.002877364, 0.002883854, 0.002881326, 0.002894596, 
    0.002888884, 0.002903763, 0.002900202, 0.002904607, 0.002902359, 
    0.002906204, 0.002902738, 0.002908736, 0.002910044, 0.002909143, 
    0.002912575, 0.002902526, 0.002906384, 0.002877352, 0.002877524, 
    0.00287832, 0.002874798, 0.002874582, 0.002871353, 0.002874218, 
    0.00287544, 0.002878536, 0.002880363, 0.0028821, 0.002885927, 0.00289019, 
    0.002896149, 0.002900429, 0.002903291, 0.002901532, 0.002903079, 
    0.002901343, 0.002900525, 0.002909546, 0.00290448, 0.002912073, 
    0.002911654, 0.00290821, 0.002911692, 0.002877639, 0.002876646, 
    0.002873213, 0.002875894, 0.002870996, 0.002873736, 0.002875305, 
    0.002881373, 0.002882704, 0.00288394, 0.002886376, 0.0028895, 
    0.002894982, 0.002899745, 0.002904092, 0.002903769, 0.002903879, 
    0.002904845, 0.002902439, 0.002905233, 0.002905698, 0.002904471, 
    0.002911588, 0.002909556, 0.002911632, 0.002910304, 0.002876964, 
    0.002878621, 0.002877719, 0.002879408, 0.002878211, 0.002883498, 
    0.002885077, 0.002892478, 0.002889438, 0.002894272, 0.002889924, 
    0.002890693, 0.002894416, 0.002890151, 0.002899471, 0.002893145, 
    0.002904879, 0.002898567, 0.002905268, 0.002904047, 0.002906056, 
    0.002907857, 0.002910118, 0.002914294, 0.002913321, 0.002916812, 
    0.002881094, 0.002883242, 0.002883053, 0.002885301, 0.002886962, 
    0.002890571, 0.002896348, 0.002894171, 0.002898155, 0.002898956, 
    0.00289289, 0.00289661, 0.002884651, 0.002886578, 0.002885428, 
    0.002881215, 0.002894643, 0.002887751, 0.002900462, 0.002896732, 
    0.002907591, 0.002902191, 0.002912786, 0.002917307, 0.002921559, 
    0.002926515, 0.002884415, 0.002882947, 0.002885563, 0.002889183, 
    0.002892535, 0.002896996, 0.002897449, 0.002898279, 0.002900438, 
    0.002902256, 0.002898534, 0.002902702, 0.00288702, 0.00289524, 
    0.002882352, 0.002886234, 0.002888926, 0.002887745, 0.002893882, 
    0.002895323, 0.002901189, 0.002898157, 0.002916181, 0.002908213, 
    0.002930286, 0.002924128, 0.002882433, 0.002884397, 0.002891239, 
    0.002887984, 0.002897286, 0.002899574, 0.002901427, 0.002903803, 
    0.002904053, 0.00290546, 0.002903148, 0.002905364, 0.002896972, 
    0.002900722, 0.002890425, 0.002892926, 0.002891772, 0.002890502, 
    0.002894402, 0.002898557, 0.002898644, 0.00289997, 0.002903712, 
    0.002897266, 0.002917193, 0.002904887, 0.00288654, 0.002890322, 
    0.002890861, 0.002889395, 0.002899336, 0.002895734, 0.002905426, 
    0.002902803, 0.002907089, 0.002904958, 0.002904637, 0.0029019, 
    0.002900187, 0.002895874, 0.002892356, 0.002889571, 0.002890212, 
    0.002893272, 0.002898803, 0.002904037, 0.002902887, 0.002906724, 
    0.002896548, 0.002900815, 0.002899159, 0.00290346, 0.0028941, 0.00290212, 
    0.002892043, 0.002892923, 0.002895654, 0.00290115, 0.002902362, 
    0.002903659, 0.002902852, 0.002898967, 0.002898326, 0.002895567, 
    0.002894801, 0.002892702, 0.002890955, 0.002892545, 0.002894206, 
    0.002898945, 0.002903204, 0.002907844, 0.00290898, 0.00291439, 
    0.00290998, 0.002917245, 0.002911058, 0.002921758, 0.002902579, 
    0.002910945, 0.002895779, 0.002897411, 0.002900365, 0.002907136, 
    0.002903478, 0.002907753, 0.0028983, 0.002893382, 0.002892108, 
    0.002889736, 0.002892157, 0.00289196, 0.002894278, 0.002893527, 
    0.002899093, 0.002896103, 0.002904588, 0.002907683, 0.00291641, 
    0.002921746, 0.002927179, 0.002929569, 0.002930297, 0.002930598,
  0.001605606, 0.001611716, 0.001610529, 0.001615453, 0.001612722, 
    0.001615945, 0.001606846, 0.001611957, 0.001608695, 0.001606157, 
    0.001624997, 0.001615672, 0.001634675, 0.001628737, 0.001643645, 
    0.001633751, 0.001645639, 0.001643361, 0.001650217, 0.001648254, 
    0.001657012, 0.001651122, 0.001661549, 0.001655607, 0.001656536, 
    0.001650928, 0.001617551, 0.001623836, 0.001617178, 0.001618075, 
    0.001617673, 0.001612778, 0.001610309, 0.00160514, 0.001606079, 
    0.001609876, 0.001618478, 0.00161556, 0.001622915, 0.001622749, 
    0.001630927, 0.001627241, 0.001640972, 0.001637072, 0.001648335, 
    0.001645505, 0.001648202, 0.001647385, 0.001648213, 0.001644061, 
    0.00164584, 0.001642185, 0.001627931, 0.001632123, 0.001619612, 
    0.001612076, 0.00160707, 0.001603514, 0.001604017, 0.001604975, 
    0.001609898, 0.001614525, 0.001618049, 0.001620404, 0.001622725, 
    0.001629741, 0.001633454, 0.001641759, 0.001640263, 0.001642799, 
    0.001645223, 0.001649289, 0.00164862, 0.00165041, 0.001642733, 
    0.001647836, 0.00163941, 0.001641715, 0.001623351, 0.001616348, 
    0.001613365, 0.001610757, 0.001604403, 0.001608791, 0.001607061, 
    0.001611177, 0.001613789, 0.001612497, 0.001620469, 0.001617371, 
    0.001633674, 0.001626657, 0.00164494, 0.00164057, 0.001645988, 
    0.001643224, 0.001647958, 0.001643697, 0.001651077, 0.001652684, 
    0.001651585, 0.001655801, 0.001643461, 0.001648202, 0.001612461, 
    0.001612672, 0.001613654, 0.001609336, 0.001609072, 0.001605114, 
    0.001608636, 0.001610135, 0.001613941, 0.001616191, 0.001618328, 
    0.001623027, 0.001628269, 0.001635595, 0.001640853, 0.001644376, 
    0.001642216, 0.001644123, 0.001641991, 0.001640992, 0.001652082, 
    0.001645856, 0.001655195, 0.001654679, 0.001650453, 0.001654737, 
    0.00161282, 0.001611607, 0.001607393, 0.001610691, 0.001604683, 
    0.001608046, 0.001609979, 0.001617434, 0.001619073, 0.00162059, 
    0.001623586, 0.001627429, 0.001634166, 0.001640022, 0.001645364, 
    0.001644973, 0.001645111, 0.001646303, 0.001643348, 0.001646788, 
    0.001647365, 0.001645856, 0.00165461, 0.001652111, 0.001654668, 
    0.001653041, 0.001612001, 0.001614042, 0.001612939, 0.001615012, 
    0.001613551, 0.001620043, 0.001621988, 0.001631084, 0.001627353, 
    0.00163329, 0.001627957, 0.001628902, 0.001633482, 0.001628246, 
    0.001639698, 0.001631934, 0.001646349, 0.001638602, 0.001646834, 
    0.001645341, 0.001647814, 0.001650027, 0.001652813, 0.001657946, 
    0.001656758, 0.001661048, 0.001617083, 0.001619727, 0.001619495, 
    0.001622262, 0.001624307, 0.001628739, 0.001635841, 0.001633171, 
    0.001638072, 0.001639055, 0.00163161, 0.001636181, 0.001621497, 
    0.001623871, 0.001622458, 0.001617291, 0.001633785, 0.001625325, 
    0.00164094, 0.001636363, 0.001649712, 0.001643076, 0.001656103, 
    0.001661661, 0.001666892, 0.001672994, 0.001621171, 0.001619375, 
    0.001622591, 0.001627038, 0.001631163, 0.001636642, 0.001637203, 
    0.001638229, 0.001640886, 0.001643118, 0.001638552, 0.001643678, 
    0.001624419, 0.00163452, 0.001618695, 0.001623462, 0.001626776, 
    0.001625324, 0.001632866, 0.001634643, 0.001641855, 0.001638128, 
    0.001660289, 0.001650493, 0.001677639, 0.001670065, 0.001618747, 
    0.001621165, 0.001629574, 0.001625574, 0.001637008, 0.001639819, 
    0.001642104, 0.001645023, 0.001645338, 0.001647067, 0.001644234, 
    0.001646955, 0.001636654, 0.00164126, 0.001628614, 0.001631694, 
    0.001630278, 0.001628723, 0.001633519, 0.001638624, 0.001638734, 
    0.00164037, 0.001644974, 0.001637055, 0.001661549, 0.00164643, 
    0.001623801, 0.001628453, 0.001629119, 0.001627317, 0.001639538, 
    0.001635112, 0.001647025, 0.001643808, 0.001649079, 0.00164646, 
    0.001646074, 0.00164271, 0.001640614, 0.001635315, 0.001631001, 
    0.001627579, 0.001628375, 0.001632133, 0.001638936, 0.001645366, 
    0.001643958, 0.001648678, 0.00163618, 0.001641423, 0.001639397, 
    0.001644679, 0.0016331, 0.001642957, 0.001630578, 0.001631664, 
    0.001635024, 0.001641777, 0.001643273, 0.001644866, 0.001643883, 
    0.001639109, 0.001638327, 0.001634943, 0.001634008, 0.001631428, 
    0.001629291, 0.001631243, 0.001633292, 0.001639112, 0.001644351, 
    0.001650059, 0.001651455, 0.001658113, 0.001652693, 0.001661633, 
    0.00165403, 0.001667187, 0.00164353, 0.001653809, 0.001635178, 
    0.001637188, 0.00164082, 0.001649147, 0.001644654, 0.001649909, 
    0.001638297, 0.001632262, 0.001630702, 0.001627787, 0.001630769, 
    0.001630526, 0.001633378, 0.001632462, 0.001639305, 0.00163563, 
    0.001646064, 0.001649868, 0.001660598, 0.001667166, 0.001673846, 
    0.001676792, 0.001677688, 0.001678063,
  0.001508832, 0.001515505, 0.001514208, 0.001519587, 0.001516604, 
    0.001520126, 0.001510186, 0.001515769, 0.001512205, 0.001509433, 
    0.001530017, 0.001519827, 0.001540595, 0.001534103, 0.001550404, 
    0.001539585, 0.001552584, 0.001550093, 0.001557591, 0.001555444, 
    0.001565028, 0.001558583, 0.001569993, 0.00156349, 0.001564507, 
    0.00155837, 0.00152188, 0.001528749, 0.001521472, 0.001522452, 
    0.001522013, 0.001516665, 0.001513969, 0.001508323, 0.001509348, 
    0.001513495, 0.001522893, 0.001519704, 0.00152774, 0.001527558, 
    0.001536497, 0.001532468, 0.00154748, 0.001543215, 0.001555533, 
    0.001552437, 0.001555388, 0.001554493, 0.0015554, 0.001550858, 
    0.001552804, 0.001548807, 0.001533222, 0.001537804, 0.001524131, 
    0.0015159, 0.00151043, 0.001506547, 0.001507096, 0.001508143, 0.00151352, 
    0.001518573, 0.001522423, 0.001524997, 0.001527532, 0.001535202, 
    0.001539261, 0.001548341, 0.001546704, 0.001549478, 0.001552129, 
    0.001556577, 0.001555845, 0.001557804, 0.001549406, 0.001554988, 
    0.001545771, 0.001548292, 0.001528219, 0.001520565, 0.001517307, 
    0.001514457, 0.001507518, 0.001512311, 0.001510422, 0.001514915, 
    0.00151777, 0.001516358, 0.001525067, 0.001521682, 0.001539501, 
    0.00153183, 0.00155182, 0.00154704, 0.001552965, 0.001549942, 
    0.001555121, 0.00155046, 0.001558533, 0.001560291, 0.001559089, 
    0.001563701, 0.001550202, 0.001555388, 0.001516319, 0.001516549, 
    0.001517621, 0.001512906, 0.001512617, 0.001508294, 0.001512141, 
    0.001513779, 0.001517935, 0.001520393, 0.001522728, 0.001527862, 
    0.001533592, 0.0015416, 0.00154735, 0.001551202, 0.00154884, 0.001550925, 
    0.001548594, 0.001547502, 0.001559632, 0.001552822, 0.001563038, 
    0.001562473, 0.00155785, 0.001562537, 0.001516711, 0.001515386, 
    0.001510784, 0.001514385, 0.001507823, 0.001511497, 0.001513608, 
    0.001521752, 0.001523541, 0.001525199, 0.001528474, 0.001532674, 
    0.001540038, 0.001546441, 0.001552283, 0.001551855, 0.001552006, 
    0.00155331, 0.001550079, 0.001553841, 0.001554472, 0.001552821, 
    0.001562398, 0.001559663, 0.001562461, 0.001560681, 0.001515816, 
    0.001518045, 0.001516841, 0.001519106, 0.00151751, 0.001524603, 
    0.001526728, 0.001536669, 0.001532591, 0.001539081, 0.001533251, 
    0.001534284, 0.001539292, 0.001533566, 0.001546088, 0.001537599, 
    0.001553361, 0.00154489, 0.001553892, 0.001552258, 0.001554963, 
    0.001557385, 0.001560432, 0.001566049, 0.001564749, 0.001569445, 
    0.001521368, 0.001524257, 0.001524003, 0.001527027, 0.001529262, 
    0.001534105, 0.001541869, 0.00153895, 0.001544308, 0.001545383, 
    0.001537243, 0.001542241, 0.001526191, 0.001528785, 0.001527241, 
    0.001521596, 0.001539622, 0.001530374, 0.001547445, 0.00154244, 
    0.001557039, 0.001549781, 0.001564033, 0.001570117, 0.001575842, 
    0.001582525, 0.001525834, 0.001523871, 0.001527386, 0.001532246, 
    0.001536755, 0.001542745, 0.001543358, 0.00154448, 0.001547385, 
    0.001549827, 0.001544834, 0.001550439, 0.001529386, 0.001540425, 
    0.001523129, 0.001528339, 0.00153196, 0.001530372, 0.001538617, 
    0.001540559, 0.001548446, 0.00154437, 0.001568615, 0.001557895, 
    0.001587612, 0.001579317, 0.001523185, 0.001525828, 0.001535018, 
    0.001530646, 0.001543145, 0.001546219, 0.001548718, 0.00155191, 
    0.001552255, 0.001554146, 0.001551047, 0.001554024, 0.001542758, 
    0.001547794, 0.001533969, 0.001537335, 0.001535787, 0.001534088, 
    0.001539331, 0.001544912, 0.001545032, 0.001546822, 0.00155186, 
    0.001543196, 0.001569996, 0.001553452, 0.001528708, 0.001533794, 
    0.001534521, 0.001532551, 0.001545911, 0.001541072, 0.0015541, 
    0.001550581, 0.001556347, 0.001553482, 0.00155306, 0.00154938, 
    0.001547088, 0.001541294, 0.001536578, 0.001532837, 0.001533707, 
    0.001537816, 0.001545254, 0.001552286, 0.001550746, 0.001555908, 
    0.00154224, 0.001547973, 0.001545757, 0.001551534, 0.001538872, 
    0.001549653, 0.001536115, 0.001537303, 0.001540976, 0.001548361, 
    0.001549996, 0.001551739, 0.001550663, 0.001545443, 0.001544588, 
    0.001540887, 0.001539865, 0.001537044, 0.001534708, 0.001536842, 
    0.001539083, 0.001545445, 0.001551175, 0.001557419, 0.001558947, 
    0.001566234, 0.001560302, 0.001570088, 0.001561767, 0.001576167, 
    0.001550279, 0.001561524, 0.001541144, 0.001543341, 0.001547314, 
    0.001556422, 0.001551507, 0.001557256, 0.001544554, 0.001537957, 
    0.001536251, 0.001533064, 0.001536323, 0.001536058, 0.001539176, 
    0.001538174, 0.001545657, 0.001541638, 0.00155305, 0.00155721, 
    0.001568952, 0.001576142, 0.001583457, 0.001586684, 0.001587666, 
    0.001588076,
  0.001433686, 0.001440472, 0.001439153, 0.001444626, 0.00144159, 
    0.001445174, 0.001435062, 0.001440742, 0.001437116, 0.001434297, 
    0.001455244, 0.00144487, 0.001466018, 0.001459404, 0.001476016, 
    0.001464989, 0.001478239, 0.001475698, 0.001483346, 0.001481155, 
    0.001490936, 0.001484357, 0.001496004, 0.001489365, 0.001490404, 
    0.00148414, 0.001446958, 0.001453953, 0.001446544, 0.001447541, 
    0.001447094, 0.001441653, 0.001438911, 0.001433167, 0.00143421, 
    0.001438428, 0.00144799, 0.001444745, 0.001452923, 0.001452739, 
    0.001461841, 0.001457737, 0.001473034, 0.001468687, 0.001481247, 
    0.001478089, 0.001481098, 0.001480186, 0.00148111, 0.001476478, 
    0.001478463, 0.001474387, 0.001458506, 0.001463174, 0.00144925, 
    0.001440875, 0.001435311, 0.001431362, 0.001431921, 0.001432985, 
    0.001438453, 0.001443594, 0.001447511, 0.001450131, 0.001452712, 
    0.001460524, 0.001464658, 0.001473913, 0.001472243, 0.001475072, 
    0.001477774, 0.001482311, 0.001481564, 0.001483563, 0.001474997, 
    0.00148069, 0.001471292, 0.001473863, 0.001453413, 0.00144562, 
    0.001442307, 0.001439407, 0.00143235, 0.001437223, 0.001435302, 
    0.001439872, 0.001442776, 0.00144134, 0.001450202, 0.001446757, 
    0.001464903, 0.001457088, 0.001477459, 0.001472586, 0.001478627, 
    0.001475545, 0.001480826, 0.001476073, 0.001484307, 0.0014861, 
    0.001484874, 0.00148958, 0.001475809, 0.001481098, 0.0014413, 
    0.001441534, 0.001442625, 0.001437828, 0.001437535, 0.001433139, 
    0.001437051, 0.001438716, 0.001442945, 0.001445445, 0.001447822, 
    0.001453048, 0.001458883, 0.001467042, 0.001472902, 0.001476829, 
    0.001474421, 0.001476547, 0.00147417, 0.001473056, 0.001485428, 
    0.001478481, 0.001488904, 0.001488327, 0.00148361, 0.001488392, 
    0.001441699, 0.001440351, 0.001435671, 0.001439333, 0.00143266, 
    0.001436395, 0.001438543, 0.001446829, 0.001448649, 0.001450337, 
    0.00145367, 0.001457947, 0.001465449, 0.001471975, 0.001477932, 
    0.001477495, 0.001477649, 0.001478979, 0.001475684, 0.00147952, 
    0.001480164, 0.001478481, 0.00148825, 0.00148546, 0.001488315, 
    0.001486498, 0.001440789, 0.001443057, 0.001441831, 0.001444136, 
    0.001442512, 0.00144973, 0.001451894, 0.001462018, 0.001457863, 
    0.001464475, 0.001458535, 0.001459587, 0.00146469, 0.001458856, 
    0.001471615, 0.001462965, 0.001479031, 0.001470395, 0.001479572, 
    0.001477906, 0.001480665, 0.001483135, 0.001486244, 0.001491977, 
    0.00149065, 0.001495444, 0.001446437, 0.001449378, 0.00144912, 
    0.001452197, 0.001454473, 0.001459405, 0.001467315, 0.001464341, 
    0.001469801, 0.001470897, 0.001462602, 0.001467695, 0.001451347, 
    0.001453988, 0.001452415, 0.001446669, 0.001465026, 0.001455607, 
    0.001472998, 0.001467897, 0.001482783, 0.001475381, 0.001489919, 
    0.001496131, 0.001501977, 0.001508807, 0.001450983, 0.001448985, 
    0.001452563, 0.001457513, 0.001462105, 0.001468208, 0.001468833, 
    0.001469976, 0.001472937, 0.001475427, 0.001470338, 0.001476051, 
    0.001454601, 0.001465844, 0.00144823, 0.001453534, 0.001457221, 
    0.001455604, 0.001464001, 0.00146598, 0.001474019, 0.001469864, 
    0.001494598, 0.001483657, 0.001514007, 0.001505528, 0.001448287, 
    0.001450977, 0.001460336, 0.001455883, 0.001468616, 0.001471749, 
    0.001474296, 0.001477552, 0.001477903, 0.001479832, 0.001476671, 
    0.001479707, 0.001468221, 0.001473355, 0.001459266, 0.001462696, 
    0.001461118, 0.001459387, 0.001464728, 0.001470418, 0.001470539, 
    0.001472363, 0.001477502, 0.001468667, 0.001496009, 0.001479126, 
    0.001453909, 0.001459089, 0.001459829, 0.001457822, 0.001471435, 
    0.001466503, 0.001479785, 0.001476196, 0.001482076, 0.001479154, 
    0.001478724, 0.001474971, 0.001472634, 0.001466729, 0.001461924, 
    0.001458113, 0.001458999, 0.001463185, 0.001470766, 0.001477935, 
    0.001476365, 0.001481629, 0.001467693, 0.001473537, 0.001471278, 
    0.001477168, 0.001464262, 0.001475252, 0.001461452, 0.001462662, 
    0.001466405, 0.001473933, 0.001475599, 0.001477377, 0.00147628, 
    0.001470958, 0.001470086, 0.001466314, 0.001465273, 0.001462399, 
    0.001460019, 0.001462193, 0.001464476, 0.00147096, 0.001476802, 
    0.00148317, 0.001484729, 0.001492167, 0.001486112, 0.001496103, 
    0.001487609, 0.001502312, 0.001475889, 0.00148736, 0.001466576, 
    0.001468815, 0.001472866, 0.001482154, 0.00147714, 0.001483004, 
    0.001470052, 0.00146333, 0.001461591, 0.001458345, 0.001461665, 
    0.001461395, 0.001464571, 0.00146355, 0.001471176, 0.00146708, 
    0.001478713, 0.001482958, 0.001494942, 0.001502285, 0.001509759, 
    0.001513058, 0.001514061, 0.001514481,
  0.001344946, 0.001351194, 0.001349979, 0.001355021, 0.001352224, 
    0.001355526, 0.001346212, 0.001351442, 0.001348103, 0.001345508, 
    0.001364814, 0.001355246, 0.001374761, 0.001368652, 0.001384006, 
    0.00137381, 0.001386063, 0.001383711, 0.00139079, 0.001388762, 
    0.001397823, 0.001391727, 0.001402524, 0.001396367, 0.00139733, 
    0.001391526, 0.00135717, 0.001363622, 0.001356788, 0.001357708, 
    0.001357295, 0.001352282, 0.001349756, 0.001344468, 0.001345428, 
    0.001349312, 0.001358122, 0.00135513, 0.001362671, 0.0013625, 
    0.001370903, 0.001367113, 0.001381247, 0.001377227, 0.001388846, 
    0.001385923, 0.001388709, 0.001387864, 0.00138872, 0.001384433, 
    0.00138627, 0.001382498, 0.001367823, 0.001372133, 0.001359283, 
    0.001351565, 0.001346442, 0.001342808, 0.001343321, 0.001344301, 
    0.001349335, 0.00135407, 0.00135768, 0.001360095, 0.001362476, 
    0.001369687, 0.001373505, 0.00138206, 0.001380515, 0.001383132, 
    0.001385632, 0.001389832, 0.001389141, 0.001390991, 0.001383063, 
    0.001388331, 0.001379635, 0.001382013, 0.001363124, 0.001355937, 
    0.001352885, 0.001350213, 0.001343716, 0.001348202, 0.001346434, 
    0.001350641, 0.001353316, 0.001351993, 0.001360161, 0.001356985, 
    0.001373731, 0.001366514, 0.001385341, 0.001380832, 0.001386421, 
    0.001383569, 0.001388457, 0.001384058, 0.00139168, 0.001393341, 
    0.001392206, 0.001396567, 0.001383814, 0.001388709, 0.001351956, 
    0.001352172, 0.001353177, 0.001348759, 0.001348489, 0.001344442, 
    0.001348043, 0.001349577, 0.001353471, 0.001355776, 0.001357967, 
    0.001362786, 0.001368172, 0.001375707, 0.001381124, 0.001384757, 
    0.001382529, 0.001384496, 0.001382297, 0.001381267, 0.001392719, 
    0.001386287, 0.001395939, 0.001395405, 0.001391036, 0.001395465, 
    0.001352323, 0.001351082, 0.001346773, 0.001350145, 0.001344002, 
    0.00134744, 0.001349418, 0.001357052, 0.001358729, 0.001360286, 
    0.00136336, 0.001367307, 0.001374235, 0.001380268, 0.001385778, 
    0.001385374, 0.001385516, 0.001386747, 0.001383698, 0.001387248, 
    0.001387844, 0.001386286, 0.001395333, 0.001392748, 0.001395394, 
    0.00139371, 0.001351485, 0.001353575, 0.001352446, 0.001354569, 
    0.001353073, 0.001359726, 0.001361722, 0.001371066, 0.00136723, 
    0.001373335, 0.00136785, 0.001368821, 0.001373535, 0.001368146, 
    0.001379935, 0.001371941, 0.001386795, 0.001378807, 0.001387296, 
    0.001385754, 0.001388307, 0.001390595, 0.001393474, 0.001398789, 
    0.001397558, 0.001402004, 0.00135669, 0.001359402, 0.001359163, 
    0.001362001, 0.001364101, 0.001368653, 0.001375959, 0.001373211, 
    0.001378257, 0.00137927, 0.001371605, 0.00137631, 0.001361217, 
    0.001363654, 0.001362203, 0.001356904, 0.001373845, 0.001365147, 
    0.001381214, 0.001376497, 0.001390269, 0.001383418, 0.00139688, 
    0.001402642, 0.001408067, 0.001414412, 0.001360882, 0.001359039, 
    0.001362339, 0.001366906, 0.001371146, 0.001376785, 0.001377362, 
    0.001378419, 0.001381157, 0.00138346, 0.001378753, 0.001384038, 
    0.00136422, 0.0013746, 0.001358342, 0.001363235, 0.001366637, 
    0.001365144, 0.001372897, 0.001374725, 0.001382158, 0.001378315, 
    0.00140122, 0.001391079, 0.001419246, 0.001411366, 0.001358395, 
    0.001360875, 0.001369512, 0.001365402, 0.001377161, 0.001380058, 
    0.001382414, 0.001385426, 0.001385751, 0.001387537, 0.001384611, 
    0.001387421, 0.001376797, 0.001381543, 0.001368524, 0.001371691, 
    0.001370234, 0.001368636, 0.001373569, 0.001378828, 0.00137894, 
    0.001380626, 0.001385382, 0.001377209, 0.00140253, 0.001386885, 
    0.00136358, 0.001368361, 0.001369044, 0.001367192, 0.001379768, 
    0.001375209, 0.001387493, 0.001384171, 0.001389614, 0.001386909, 
    0.001386511, 0.001383038, 0.001380877, 0.001375418, 0.001370979, 
    0.00136746, 0.001368278, 0.001372144, 0.001379149, 0.001385781, 
    0.001384328, 0.001389201, 0.001376308, 0.001381712, 0.001379623, 
    0.001385071, 0.001373138, 0.0013833, 0.001370543, 0.00137166, 
    0.001375119, 0.001382079, 0.001383619, 0.001385265, 0.001384249, 
    0.001379327, 0.001378521, 0.001375035, 0.001374072, 0.001371417, 
    0.001369219, 0.001371227, 0.001373337, 0.001379329, 0.001384733, 
    0.001390628, 0.001392071, 0.001398966, 0.001393353, 0.001402617, 
    0.001394741, 0.001408379, 0.001383888, 0.001394509, 0.001375276, 
    0.001377346, 0.001381092, 0.001389687, 0.001385045, 0.001390474, 
    0.001378489, 0.001372278, 0.001370671, 0.001367674, 0.001370739, 
    0.00137049, 0.001373424, 0.001372481, 0.001379528, 0.001375742, 
    0.001386502, 0.001390431, 0.001401538, 0.001408353, 0.001415296, 
    0.001418363, 0.001419297, 0.001419687,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.222765e-06, 1.23331e-06, 1.231256e-06, 1.239789e-06, 1.235052e-06, 
    1.240644e-06, 1.224898e-06, 1.233729e-06, 1.228088e-06, 1.223711e-06, 
    1.256432e-06, 1.240169e-06, 1.273445e-06, 1.262986e-06, 1.289345e-06, 
    1.271814e-06, 1.292895e-06, 1.288837e-06, 1.30107e-06, 1.297559e-06, 
    1.31327e-06, 1.302691e-06, 1.321453e-06, 1.31074e-06, 1.312412e-06, 
    1.302342e-06, 1.243434e-06, 1.254402e-06, 1.242786e-06, 1.244346e-06, 
    1.243646e-06, 1.235149e-06, 1.230878e-06, 1.22196e-06, 1.223576e-06, 
    1.230128e-06, 1.245047e-06, 1.239972e-06, 1.252784e-06, 1.252494e-06, 
    1.266835e-06, 1.260358e-06, 1.284591e-06, 1.277679e-06, 1.297705e-06, 
    1.292653e-06, 1.297467e-06, 1.296006e-06, 1.297486e-06, 1.290081e-06, 
    1.293251e-06, 1.286745e-06, 1.261571e-06, 1.268943e-06, 1.247022e-06, 
    1.233935e-06, 1.225284e-06, 1.219165e-06, 1.220028e-06, 1.221677e-06, 
    1.230166e-06, 1.238175e-06, 1.244297e-06, 1.248401e-06, 1.252452e-06, 
    1.264753e-06, 1.27129e-06, 1.28599e-06, 1.283331e-06, 1.287837e-06, 
    1.292151e-06, 1.299409e-06, 1.298213e-06, 1.301416e-06, 1.287718e-06, 
    1.296813e-06, 1.281816e-06, 1.285909e-06, 1.253554e-06, 1.241341e-06, 
    1.236168e-06, 1.23165e-06, 1.220693e-06, 1.228254e-06, 1.22527e-06, 
    1.232374e-06, 1.236899e-06, 1.23466e-06, 1.248513e-06, 1.243118e-06, 
    1.271678e-06, 1.259334e-06, 1.291648e-06, 1.283876e-06, 1.293514e-06, 
    1.288591e-06, 1.297031e-06, 1.289434e-06, 1.302609e-06, 1.305488e-06, 
    1.303519e-06, 1.311086e-06, 1.289012e-06, 1.297466e-06, 1.234598e-06, 
    1.234963e-06, 1.236664e-06, 1.229194e-06, 1.228738e-06, 1.221915e-06, 
    1.227985e-06, 1.230574e-06, 1.237162e-06, 1.241066e-06, 1.244784e-06, 
    1.252979e-06, 1.262164e-06, 1.275067e-06, 1.284379e-06, 1.290641e-06, 
    1.286799e-06, 1.29019e-06, 1.286399e-06, 1.284625e-06, 1.304409e-06, 
    1.29328e-06, 1.309996e-06, 1.309068e-06, 1.301491e-06, 1.309172e-06, 
    1.235219e-06, 1.233119e-06, 1.225842e-06, 1.231535e-06, 1.221173e-06, 
    1.226967e-06, 1.230305e-06, 1.24323e-06, 1.246079e-06, 1.248724e-06, 
    1.253956e-06, 1.260688e-06, 1.272543e-06, 1.282904e-06, 1.292402e-06, 
    1.291704e-06, 1.29195e-06, 1.294076e-06, 1.288812e-06, 1.29494e-06, 
    1.29597e-06, 1.293278e-06, 1.308943e-06, 1.304458e-06, 1.309048e-06, 
    1.306126e-06, 1.233801e-06, 1.237337e-06, 1.235425e-06, 1.239021e-06, 
    1.236487e-06, 1.247772e-06, 1.251166e-06, 1.267112e-06, 1.260555e-06, 
    1.270999e-06, 1.261614e-06, 1.263274e-06, 1.271339e-06, 1.26212e-06, 
    1.282331e-06, 1.268609e-06, 1.294158e-06, 1.280389e-06, 1.295023e-06, 
    1.292359e-06, 1.296771e-06, 1.300729e-06, 1.305717e-06, 1.314947e-06, 
    1.312806e-06, 1.320545e-06, 1.242617e-06, 1.247221e-06, 1.246816e-06, 
    1.251642e-06, 1.255218e-06, 1.262988e-06, 1.2755e-06, 1.270787e-06, 
    1.279446e-06, 1.281188e-06, 1.268035e-06, 1.276102e-06, 1.250306e-06, 
    1.254455e-06, 1.251984e-06, 1.242978e-06, 1.271871e-06, 1.256999e-06, 
    1.284532e-06, 1.276422e-06, 1.300163e-06, 1.288328e-06, 1.311629e-06, 
    1.321655e-06, 1.331129e-06, 1.342243e-06, 1.249738e-06, 1.246605e-06, 
    1.252217e-06, 1.260003e-06, 1.26725e-06, 1.276917e-06, 1.277909e-06, 
    1.279725e-06, 1.284435e-06, 1.288403e-06, 1.280299e-06, 1.289398e-06, 
    1.255417e-06, 1.273166e-06, 1.24542e-06, 1.253741e-06, 1.259541e-06, 
    1.256995e-06, 1.270247e-06, 1.273381e-06, 1.286157e-06, 1.279544e-06, 
    1.319176e-06, 1.301564e-06, 1.350739e-06, 1.336901e-06, 1.245511e-06, 
    1.249726e-06, 1.264455e-06, 1.257436e-06, 1.277564e-06, 1.282544e-06, 
    1.2866e-06, 1.291794e-06, 1.292355e-06, 1.295439e-06, 1.290388e-06, 
    1.295239e-06, 1.276937e-06, 1.285099e-06, 1.262766e-06, 1.268182e-06, 
    1.265689e-06, 1.262957e-06, 1.271398e-06, 1.280424e-06, 1.280618e-06, 
    1.283519e-06, 1.291712e-06, 1.277643e-06, 1.321457e-06, 1.294306e-06, 
    1.254332e-06, 1.262487e-06, 1.263654e-06, 1.26049e-06, 1.282044e-06, 
    1.274212e-06, 1.295364e-06, 1.289629e-06, 1.299031e-06, 1.294355e-06, 
    1.293667e-06, 1.287675e-06, 1.283951e-06, 1.274569e-06, 1.266962e-06, 
    1.260947e-06, 1.262344e-06, 1.268956e-06, 1.280977e-06, 1.292404e-06, 
    1.289896e-06, 1.298314e-06, 1.276096e-06, 1.285388e-06, 1.281792e-06, 
    1.291178e-06, 1.270661e-06, 1.288123e-06, 1.266218e-06, 1.26813e-06, 
    1.274056e-06, 1.286021e-06, 1.288676e-06, 1.291514e-06, 1.289763e-06, 
    1.281284e-06, 1.279898e-06, 1.273911e-06, 1.272261e-06, 1.267712e-06, 
    1.263953e-06, 1.267387e-06, 1.270999e-06, 1.281287e-06, 1.290595e-06, 
    1.300783e-06, 1.303283e-06, 1.315251e-06, 1.305504e-06, 1.321608e-06, 
    1.307909e-06, 1.33167e-06, 1.289139e-06, 1.307511e-06, 1.274327e-06, 
    1.27788e-06, 1.28432e-06, 1.299156e-06, 1.291136e-06, 1.300518e-06, 
    1.279844e-06, 1.269185e-06, 1.266435e-06, 1.261312e-06, 1.266552e-06, 
    1.266125e-06, 1.271149e-06, 1.269533e-06, 1.281629e-06, 1.275124e-06, 
    1.293648e-06, 1.300442e-06, 1.319731e-06, 1.331627e-06, 1.343795e-06, 
    1.349185e-06, 1.350828e-06, 1.351515e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  7.717309e-06, 7.75199e-06, 7.745231e-06, 7.773217e-06, 7.757685e-06, 
    7.775997e-06, 7.724302e-06, 7.753305e-06, 7.73478e-06, 7.720369e-06, 
    7.827509e-06, 7.774403e-06, 7.882823e-06, 7.848861e-06, 7.934218e-06, 
    7.877507e-06, 7.945659e-06, 7.932575e-06, 7.971967e-06, 7.960664e-06, 
    8.011064e-06, 7.977156e-06, 8.037227e-06, 8.002959e-06, 8.008301e-06, 
    7.975996e-06, 7.785155e-06, 7.820949e-06, 7.783016e-06, 7.78812e-06, 
    7.785823e-06, 7.757965e-06, 7.74393e-06, 7.714595e-06, 7.719908e-06, 
    7.741453e-06, 7.790355e-06, 7.77374e-06, 7.815617e-06, 7.814673e-06, 
    7.861342e-06, 7.840285e-06, 7.918856e-06, 7.896493e-06, 7.961126e-06, 
    7.944844e-06, 7.960342e-06, 7.95563e-06, 7.96038e-06, 7.936525e-06, 
    7.946725e-06, 7.925748e-06, 7.844323e-06, 7.868267e-06, 7.796855e-06, 
    7.75396e-06, 7.725537e-06, 7.705382e-06, 7.708212e-06, 7.713643e-06, 
    7.741563e-06, 7.767846e-06, 7.787893e-06, 7.801296e-06, 7.814513e-06, 
    7.854546e-06, 7.875778e-06, 7.92335e-06, 7.914767e-06, 7.9293e-06, 
    7.943217e-06, 7.966571e-06, 7.962723e-06, 7.973004e-06, 7.928882e-06, 
    7.95819e-06, 7.909805e-06, 7.923028e-06, 7.818141e-06, 7.778258e-06, 
    7.761279e-06, 7.746453e-06, 7.710396e-06, 7.735283e-06, 7.725459e-06, 
    7.748809e-06, 7.763653e-06, 7.756299e-06, 7.801655e-06, 7.783998e-06, 
    7.877024e-06, 7.836918e-06, 7.941604e-06, 7.91651e-06, 7.947597e-06, 
    7.93173e-06, 7.958902e-06, 7.934432e-06, 7.976824e-06, 7.986071e-06, 
    7.979731e-06, 8.004014e-06, 7.933023e-06, 7.960255e-06, 7.756139e-06, 
    7.757338e-06, 7.76291e-06, 7.738362e-06, 7.736861e-06, 7.714398e-06, 
    7.734368e-06, 7.742878e-06, 7.764496e-06, 7.777276e-06, 7.789432e-06, 
    7.816205e-06, 7.84611e-06, 7.887991e-06, 7.918125e-06, 7.938328e-06, 
    7.925931e-06, 7.936859e-06, 7.924623e-06, 7.91888e-06, 7.982582e-06, 
    7.946785e-06, 8.000497e-06, 7.997527e-06, 7.973183e-06, 7.997838e-06, 
    7.758163e-06, 7.75126e-06, 7.727333e-06, 7.746042e-06, 7.711938e-06, 
    7.731012e-06, 7.74197e-06, 7.784343e-06, 7.793666e-06, 7.802308e-06, 
    7.819381e-06, 7.8413e-06, 7.879802e-06, 7.913337e-06, 7.943996e-06, 
    7.941737e-06, 7.942524e-06, 7.949358e-06, 7.932387e-06, 7.952129e-06, 
    7.955428e-06, 7.946765e-06, 7.997104e-06, 7.982716e-06, 7.997431e-06, 
    7.988048e-06, 7.753492e-06, 7.765076e-06, 7.758797e-06, 7.770584e-06, 
    7.762259e-06, 7.799198e-06, 7.81027e-06, 7.862182e-06, 7.840865e-06, 
    7.874798e-06, 7.844297e-06, 7.849696e-06, 7.875856e-06, 7.845926e-06, 
    7.911451e-06, 7.866977e-06, 7.949615e-06, 7.905132e-06, 7.952386e-06, 
    7.943795e-06, 7.957993e-06, 7.97072e-06, 7.986735e-06, 8.016305e-06, 
    8.009441e-06, 8.034193e-06, 7.782367e-06, 7.797405e-06, 7.796086e-06, 
    7.811838e-06, 7.82349e-06, 7.848795e-06, 7.889396e-06, 7.874109e-06, 
    7.902157e-06, 7.90779e-06, 7.865153e-06, 7.891306e-06, 7.807405e-06, 
    7.820921e-06, 7.81287e-06, 7.783422e-06, 7.877546e-06, 7.829186e-06, 
    7.918523e-06, 7.89228e-06, 7.96888e-06, 7.93075e-06, 8.005663e-06, 
    8.037714e-06, 8.067939e-06, 8.103236e-06, 7.805625e-06, 7.79538e-06, 
    7.8137e-06, 7.839062e-06, 7.862621e-06, 7.893977e-06, 7.897182e-06, 
    7.903043e-06, 7.918267e-06, 7.931078e-06, 7.904872e-06, 7.934268e-06, 
    7.824031e-06, 7.881748e-06, 7.791396e-06, 7.818561e-06, 7.837456e-06, 
    7.82917e-06, 7.872259e-06, 7.882409e-06, 7.923724e-06, 7.902362e-06, 
    8.029769e-06, 7.973333e-06, 8.13016e-06, 8.08626e-06, 7.791794e-06, 
    7.805559e-06, 7.853529e-06, 7.830694e-06, 7.896053e-06, 7.912162e-06, 
    7.925252e-06, 7.942002e-06, 7.9438e-06, 7.953731e-06, 7.937443e-06, 
    7.953076e-06, 7.893955e-06, 7.920357e-06, 7.847962e-06, 7.865547e-06, 
    7.85745e-06, 7.848555e-06, 7.875965e-06, 7.905189e-06, 7.905818e-06, 
    7.915179e-06, 7.941572e-06, 7.896166e-06, 8.036996e-06, 7.94991e-06, 
    7.820579e-06, 7.84711e-06, 7.850912e-06, 7.840624e-06, 7.910522e-06, 
    7.885172e-06, 7.953491e-06, 7.935001e-06, 7.965274e-06, 7.950222e-06, 
    7.947989e-06, 7.928672e-06, 7.916627e-06, 7.886266e-06, 7.861568e-06, 
    7.842021e-06, 7.846548e-06, 7.868029e-06, 7.906957e-06, 7.943855e-06, 
    7.935756e-06, 7.962867e-06, 7.891138e-06, 7.921186e-06, 7.909546e-06, 
    7.939862e-06, 7.873666e-06, 7.930128e-06, 7.859235e-06, 7.865434e-06, 
    7.884645e-06, 7.92334e-06, 7.931912e-06, 7.941059e-06, 7.9354e-06, 
    7.90801e-06, 7.903521e-06, 7.884127e-06, 7.878759e-06, 7.864009e-06, 
    7.851773e-06, 7.862933e-06, 7.874633e-06, 7.907963e-06, 7.938006e-06, 
    7.970796e-06, 7.978831e-06, 8.017159e-06, 7.985926e-06, 8.037438e-06, 
    7.993591e-06, 8.069524e-06, 7.933402e-06, 7.992505e-06, 7.885526e-06, 
    7.897024e-06, 7.917833e-06, 7.965638e-06, 7.939821e-06, 7.970013e-06, 
    7.903341e-06, 7.868775e-06, 7.85985e-06, 7.843194e-06, 7.860215e-06, 
    7.858831e-06, 7.875131e-06, 7.869877e-06, 7.909046e-06, 7.887998e-06, 
    7.947819e-06, 7.969679e-06, 8.031497e-06, 8.069422e-06, 8.108103e-06, 
    8.125172e-06, 8.130371e-06, 8.132535e-06,
  4.029571e-06, 4.060347e-06, 4.054359e-06, 4.07923e-06, 4.065429e-06, 
    4.081723e-06, 4.035807e-06, 4.061568e-06, 4.045117e-06, 4.032343e-06, 
    4.127653e-06, 4.080342e-06, 4.177049e-06, 4.146708e-06, 4.223094e-06, 
    4.172317e-06, 4.233362e-06, 4.221634e-06, 4.256989e-06, 4.24685e-06, 
    4.29218e-06, 4.261672e-06, 4.315757e-06, 4.284892e-06, 4.289712e-06, 
    4.260666e-06, 4.089853e-06, 4.121749e-06, 4.087964e-06, 4.092507e-06, 
    4.09047e-06, 4.065711e-06, 4.053252e-06, 4.027228e-06, 4.031949e-06, 
    4.051068e-06, 4.09455e-06, 4.079774e-06, 4.117066e-06, 4.116222e-06, 
    4.157883e-06, 4.139079e-06, 4.209346e-06, 4.189331e-06, 4.247272e-06, 
    4.232671e-06, 4.246585e-06, 4.242365e-06, 4.24664e-06, 4.225234e-06, 
    4.2344e-06, 4.215585e-06, 4.142597e-06, 4.163995e-06, 4.100296e-06, 
    4.062166e-06, 4.036934e-06, 4.019061e-06, 4.021585e-06, 4.026399e-06, 
    4.05118e-06, 4.074538e-06, 4.092372e-06, 4.104317e-06, 4.116101e-06, 
    4.151829e-06, 4.170803e-06, 4.213394e-06, 4.205702e-06, 4.218741e-06, 
    4.23122e-06, 4.252195e-06, 4.248741e-06, 4.25799e-06, 4.218401e-06, 
    4.244695e-06, 4.201321e-06, 4.213166e-06, 4.119282e-06, 4.083759e-06, 
    4.068675e-06, 4.055509e-06, 4.023527e-06, 4.045601e-06, 4.036893e-06, 
    4.057627e-06, 4.07082e-06, 4.064294e-06, 4.104644e-06, 4.088938e-06, 
    4.171928e-06, 4.136104e-06, 4.229764e-06, 4.207281e-06, 4.235161e-06, 
    4.220927e-06, 4.245325e-06, 4.223365e-06, 4.261437e-06, 4.269747e-06, 
    4.264065e-06, 4.285897e-06, 4.222148e-06, 4.246583e-06, 4.06411e-06, 
    4.065174e-06, 4.070135e-06, 4.048346e-06, 4.047015e-06, 4.027097e-06, 
    4.044821e-06, 4.052375e-06, 4.071587e-06, 4.082963e-06, 4.09379e-06, 
    4.117634e-06, 4.144322e-06, 4.181758e-06, 4.208736e-06, 4.226856e-06, 
    4.215744e-06, 4.225553e-06, 4.214587e-06, 4.209451e-06, 4.266633e-06, 
    4.234484e-06, 4.282756e-06, 4.28008e-06, 4.258209e-06, 4.280382e-06, 
    4.065922e-06, 4.059799e-06, 4.038564e-06, 4.055179e-06, 4.024931e-06, 
    4.041848e-06, 4.051587e-06, 4.089261e-06, 4.097561e-06, 4.105257e-06, 
    4.120478e-06, 4.14004e-06, 4.174442e-06, 4.204465e-06, 4.231948e-06, 
    4.229933e-06, 4.230642e-06, 4.236787e-06, 4.221567e-06, 4.239288e-06, 
    4.242262e-06, 4.234483e-06, 4.279722e-06, 4.266782e-06, 4.280023e-06, 
    4.271597e-06, 4.06179e-06, 4.072096e-06, 4.066525e-06, 4.077002e-06, 
    4.069618e-06, 4.102483e-06, 4.112357e-06, 4.158685e-06, 4.139654e-06, 
    4.169964e-06, 4.142731e-06, 4.14755e-06, 4.170944e-06, 4.144202e-06, 
    4.202803e-06, 4.16303e-06, 4.237026e-06, 4.197176e-06, 4.239527e-06, 
    4.231829e-06, 4.24458e-06, 4.25601e-06, 4.270417e-06, 4.297026e-06, 
    4.29086e-06, 4.313152e-06, 4.087482e-06, 4.100882e-06, 4.099706e-06, 
    4.113749e-06, 4.124145e-06, 4.146719e-06, 4.183017e-06, 4.169355e-06, 
    4.194455e-06, 4.199499e-06, 4.161374e-06, 4.184762e-06, 4.109862e-06, 
    4.121924e-06, 4.114744e-06, 4.088535e-06, 4.172495e-06, 4.129322e-06, 
    4.209182e-06, 4.185696e-06, 4.254379e-06, 4.220164e-06, 4.287466e-06, 
    4.316341e-06, 4.343605e-06, 4.375519e-06, 4.108207e-06, 4.099093e-06, 
    4.115421e-06, 4.138044e-06, 4.15909e-06, 4.187126e-06, 4.190001e-06, 
    4.195261e-06, 4.208903e-06, 4.220384e-06, 4.19692e-06, 4.223265e-06, 
    4.124714e-06, 4.176253e-06, 4.095645e-06, 4.119849e-06, 4.136711e-06, 
    4.129316e-06, 4.167796e-06, 4.176883e-06, 4.213886e-06, 4.194745e-06, 
    4.309203e-06, 4.258419e-06, 4.399893e-06, 4.360185e-06, 4.095909e-06, 
    4.108178e-06, 4.150977e-06, 4.130593e-06, 4.189002e-06, 4.203425e-06, 
    4.215168e-06, 4.230189e-06, 4.231816e-06, 4.240727e-06, 4.226127e-06, 
    4.240152e-06, 4.187185e-06, 4.210824e-06, 4.146082e-06, 4.161802e-06, 
    4.154569e-06, 4.146637e-06, 4.171136e-06, 4.197288e-06, 4.197855e-06, 
    4.206253e-06, 4.229938e-06, 4.18924e-06, 4.315759e-06, 4.237443e-06, 
    4.121571e-06, 4.145259e-06, 4.148656e-06, 4.13947e-06, 4.201978e-06, 
    4.179287e-06, 4.24051e-06, 4.223933e-06, 4.25111e-06, 4.237596e-06, 
    4.235609e-06, 4.218281e-06, 4.207504e-06, 4.180325e-06, 4.158262e-06, 
    4.140803e-06, 4.14486e-06, 4.164048e-06, 4.198891e-06, 4.231959e-06, 
    4.224706e-06, 4.249042e-06, 4.184757e-06, 4.211664e-06, 4.201254e-06, 
    4.228419e-06, 4.16899e-06, 4.219554e-06, 4.1561e-06, 4.161651e-06, 
    4.178837e-06, 4.213486e-06, 4.221178e-06, 4.229383e-06, 4.22432e-06, 
    4.199779e-06, 4.195766e-06, 4.178421e-06, 4.173633e-06, 4.160443e-06, 
    4.14953e-06, 4.159498e-06, 4.169974e-06, 4.199792e-06, 4.226728e-06, 
    4.256172e-06, 4.263392e-06, 4.297898e-06, 4.269795e-06, 4.316195e-06, 
    4.276719e-06, 4.345147e-06, 4.222503e-06, 4.275576e-06, 4.179622e-06, 
    4.189922e-06, 4.208566e-06, 4.251462e-06, 4.228291e-06, 4.255397e-06, 
    4.19561e-06, 4.164707e-06, 4.156735e-06, 4.141862e-06, 4.157076e-06, 
    4.155838e-06, 4.170413e-06, 4.165728e-06, 4.200784e-06, 4.18194e-06, 
    4.235557e-06, 4.255185e-06, 4.310811e-06, 4.345035e-06, 4.379986e-06, 
    4.395445e-06, 4.400154e-06, 4.402123e-06,
  3.819898e-06, 3.853829e-06, 3.847224e-06, 3.874663e-06, 3.859433e-06, 
    3.877414e-06, 3.826769e-06, 3.855177e-06, 3.837032e-06, 3.82295e-06, 
    3.928147e-06, 3.875889e-06, 3.982765e-06, 3.9492e-06, 4.033751e-06, 
    3.977531e-06, 4.045129e-06, 4.032129e-06, 4.071319e-06, 4.060076e-06, 
    4.110373e-06, 4.076514e-06, 4.136552e-06, 4.102279e-06, 4.107631e-06, 
    4.075398e-06, 3.886385e-06, 3.921623e-06, 3.884301e-06, 3.889317e-06, 
    3.887067e-06, 3.859745e-06, 3.846006e-06, 3.817313e-06, 3.822516e-06, 
    3.843595e-06, 3.891573e-06, 3.875261e-06, 3.916437e-06, 3.915505e-06, 
    3.961557e-06, 3.940765e-06, 4.018517e-06, 3.996353e-06, 4.060545e-06, 
    4.04436e-06, 4.059784e-06, 4.055105e-06, 4.059845e-06, 4.036119e-06, 
    4.046276e-06, 4.025427e-06, 3.944655e-06, 3.968319e-06, 3.897917e-06, 
    3.855841e-06, 3.828012e-06, 3.808314e-06, 3.811096e-06, 3.816401e-06, 
    3.843719e-06, 3.869482e-06, 3.889166e-06, 3.902355e-06, 3.915371e-06, 
    3.954869e-06, 3.975853e-06, 4.023002e-06, 4.01448e-06, 4.028926e-06, 
    4.042752e-06, 4.066005e-06, 4.062174e-06, 4.072432e-06, 4.028547e-06, 
    4.057689e-06, 4.009628e-06, 4.022748e-06, 3.918899e-06, 3.879659e-06, 
    3.863021e-06, 3.848492e-06, 3.813235e-06, 3.837567e-06, 3.827967e-06, 
    3.850826e-06, 3.86538e-06, 3.85818e-06, 3.902716e-06, 3.885375e-06, 
    3.977098e-06, 3.937478e-06, 4.041138e-06, 4.016229e-06, 4.047119e-06, 
    4.031344e-06, 4.058387e-06, 4.034046e-06, 4.076253e-06, 4.085472e-06, 
    4.07917e-06, 4.103392e-06, 4.032698e-06, 4.059782e-06, 3.857977e-06, 
    3.859151e-06, 3.864624e-06, 3.840593e-06, 3.839126e-06, 3.81717e-06, 
    3.836705e-06, 3.845036e-06, 3.866226e-06, 3.87878e-06, 3.890732e-06, 
    3.917065e-06, 3.946564e-06, 3.987974e-06, 4.017842e-06, 4.037914e-06, 
    4.025602e-06, 4.036471e-06, 4.024321e-06, 4.018632e-06, 4.082018e-06, 
    4.046371e-06, 4.099905e-06, 4.096936e-06, 4.072675e-06, 4.09727e-06, 
    3.859976e-06, 3.853222e-06, 3.829808e-06, 3.848126e-06, 3.814782e-06, 
    3.833429e-06, 3.844169e-06, 3.885734e-06, 3.894896e-06, 3.903394e-06, 
    3.920207e-06, 3.941828e-06, 3.979877e-06, 4.013113e-06, 4.043557e-06, 
    4.041323e-06, 4.04211e-06, 4.048922e-06, 4.032055e-06, 4.051694e-06, 
    4.054992e-06, 4.046368e-06, 4.096538e-06, 4.08218e-06, 4.096873e-06, 
    4.087522e-06, 3.855417e-06, 3.866788e-06, 3.860641e-06, 3.872202e-06, 
    3.864055e-06, 3.900334e-06, 3.91124e-06, 3.962448e-06, 3.941401e-06, 
    3.974923e-06, 3.944801e-06, 3.950131e-06, 3.976013e-06, 3.946428e-06, 
    4.011274e-06, 3.967256e-06, 4.049186e-06, 4.005047e-06, 4.051959e-06, 
    4.043425e-06, 4.05756e-06, 4.070236e-06, 4.086213e-06, 4.115749e-06, 
    4.108902e-06, 4.133657e-06, 3.883767e-06, 3.898564e-06, 3.897263e-06, 
    3.912773e-06, 3.92426e-06, 3.949211e-06, 3.989366e-06, 3.974246e-06, 
    4.002025e-06, 4.007612e-06, 3.965417e-06, 3.991298e-06, 3.908482e-06, 
    3.921809e-06, 3.913874e-06, 3.884932e-06, 3.977725e-06, 3.929984e-06, 
    4.018335e-06, 3.99233e-06, 4.068427e-06, 4.030504e-06, 4.105135e-06, 
    4.137205e-06, 4.167497e-06, 4.202998e-06, 3.906652e-06, 3.896586e-06, 
    3.91462e-06, 3.939624e-06, 3.962893e-06, 3.993914e-06, 3.997095e-06, 
    4.002919e-06, 4.018025e-06, 4.030744e-06, 4.004759e-06, 4.033935e-06, 
    3.924898e-06, 3.981881e-06, 3.892781e-06, 3.919517e-06, 3.938149e-06, 
    3.929974e-06, 3.972521e-06, 3.982576e-06, 4.023548e-06, 4.002347e-06, 
    4.129277e-06, 4.072911e-06, 4.230124e-06, 4.185938e-06, 3.893071e-06, 
    3.906619e-06, 3.953922e-06, 3.931385e-06, 3.99599e-06, 4.011959e-06, 
    4.024964e-06, 4.04161e-06, 4.043411e-06, 4.05329e-06, 4.037107e-06, 
    4.052651e-06, 3.99398e-06, 4.020154e-06, 3.948506e-06, 3.965892e-06, 
    3.95789e-06, 3.94912e-06, 3.976216e-06, 4.005166e-06, 4.00579e-06, 
    4.015092e-06, 4.041346e-06, 3.996252e-06, 4.136567e-06, 4.049662e-06, 
    3.921414e-06, 3.947602e-06, 3.951354e-06, 3.941195e-06, 4.010357e-06, 
    3.985238e-06, 4.053049e-06, 4.034675e-06, 4.0648e-06, 4.049818e-06, 
    4.047616e-06, 4.028414e-06, 4.016476e-06, 3.986387e-06, 3.961977e-06, 
    3.942669e-06, 3.947155e-06, 3.968378e-06, 4.006941e-06, 4.043572e-06, 
    4.035535e-06, 4.062507e-06, 3.99129e-06, 4.021086e-06, 4.009557e-06, 
    4.039648e-06, 3.973844e-06, 4.029837e-06, 3.959584e-06, 3.965723e-06, 
    3.98474e-06, 4.023107e-06, 4.031623e-06, 4.040716e-06, 4.035105e-06, 
    4.007923e-06, 4.003479e-06, 3.984278e-06, 3.978981e-06, 3.964386e-06, 
    3.952319e-06, 3.963343e-06, 3.974933e-06, 4.007936e-06, 4.037775e-06, 
    4.070415e-06, 4.078422e-06, 4.116724e-06, 4.085531e-06, 4.137053e-06, 
    4.093224e-06, 4.169223e-06, 4.033099e-06, 4.091946e-06, 3.985607e-06, 
    3.997007e-06, 4.017656e-06, 4.065196e-06, 4.039506e-06, 4.06956e-06, 
    4.003306e-06, 3.969109e-06, 3.960286e-06, 3.943841e-06, 3.960663e-06, 
    3.959294e-06, 3.975417e-06, 3.970233e-06, 4.009034e-06, 3.988172e-06, 
    4.047559e-06, 4.069323e-06, 4.131058e-06, 4.169091e-06, 4.207962e-06, 
    4.225169e-06, 4.230412e-06, 4.232605e-06,
  3.894142e-06, 3.931183e-06, 3.923969e-06, 3.953942e-06, 3.937302e-06, 
    3.956948e-06, 3.901638e-06, 3.932657e-06, 3.912842e-06, 3.89747e-06, 
    4.012422e-06, 3.955282e-06, 4.0722e-06, 4.035449e-06, 4.128075e-06, 
    4.06647e-06, 4.140551e-06, 4.126292e-06, 4.169281e-06, 4.156943e-06, 
    4.212162e-06, 4.174981e-06, 4.240923e-06, 4.20327e-06, 4.209149e-06, 
    4.173757e-06, 3.96675e-06, 4.005286e-06, 3.964472e-06, 3.969955e-06, 
    3.967495e-06, 3.937645e-06, 3.922643e-06, 3.891318e-06, 3.896996e-06, 
    3.920009e-06, 3.972422e-06, 3.954593e-06, 3.999603e-06, 3.998583e-06, 
    4.048975e-06, 4.026217e-06, 4.111369e-06, 4.08708e-06, 4.157458e-06, 
    4.139704e-06, 4.156623e-06, 4.15149e-06, 4.15669e-06, 4.130667e-06, 
    4.141807e-06, 4.118944e-06, 4.030474e-06, 4.056378e-06, 3.979356e-06, 
    3.933385e-06, 3.902996e-06, 3.8815e-06, 3.884535e-06, 3.890325e-06, 
    3.920144e-06, 3.94828e-06, 3.969788e-06, 3.984206e-06, 3.998437e-06, 
    4.04166e-06, 4.064631e-06, 4.116288e-06, 4.106943e-06, 4.122781e-06, 
    4.13794e-06, 4.163449e-06, 4.159246e-06, 4.170503e-06, 4.122364e-06, 
    4.154327e-06, 4.101625e-06, 4.116007e-06, 4.002307e-06, 3.959399e-06, 
    3.941227e-06, 3.925355e-06, 3.88687e-06, 3.913427e-06, 3.902948e-06, 
    3.927903e-06, 3.943799e-06, 3.935933e-06, 3.9846e-06, 3.965645e-06, 
    4.065994e-06, 4.022622e-06, 4.13617e-06, 4.108861e-06, 4.142729e-06, 
    4.125431e-06, 4.155092e-06, 4.128392e-06, 4.174696e-06, 4.184815e-06, 
    4.177898e-06, 4.204489e-06, 4.126915e-06, 4.156623e-06, 3.935712e-06, 
    3.936995e-06, 3.942971e-06, 3.916731e-06, 3.915129e-06, 3.891162e-06, 
    3.912485e-06, 3.921582e-06, 3.944721e-06, 3.958439e-06, 3.971501e-06, 
    4.000292e-06, 4.032565e-06, 4.077904e-06, 4.110628e-06, 4.132634e-06, 
    4.119134e-06, 4.131052e-06, 4.11773e-06, 4.111494e-06, 4.181023e-06, 
    4.141911e-06, 4.20066e-06, 4.197399e-06, 4.170771e-06, 4.197767e-06, 
    3.937895e-06, 3.930518e-06, 3.904956e-06, 3.924954e-06, 3.888556e-06, 
    3.90891e-06, 3.920635e-06, 3.96604e-06, 3.976051e-06, 3.985343e-06, 
    4.003727e-06, 4.02738e-06, 4.069035e-06, 4.105446e-06, 4.138823e-06, 
    4.136373e-06, 4.137235e-06, 4.144707e-06, 4.12621e-06, 4.147748e-06, 
    4.151368e-06, 4.141906e-06, 4.196963e-06, 4.181199e-06, 4.19733e-06, 
    4.187063e-06, 3.932916e-06, 3.945336e-06, 3.938622e-06, 3.951252e-06, 
    3.942352e-06, 3.982e-06, 3.993925e-06, 4.049952e-06, 4.026914e-06, 
    4.063611e-06, 4.030634e-06, 4.036468e-06, 4.064809e-06, 4.032413e-06, 
    4.103434e-06, 4.055218e-06, 4.144998e-06, 4.096613e-06, 4.148039e-06, 
    4.138678e-06, 4.154183e-06, 4.168092e-06, 4.185626e-06, 4.218065e-06, 
    4.210543e-06, 4.23774e-06, 3.963888e-06, 3.980063e-06, 3.978638e-06, 
    3.995597e-06, 4.008161e-06, 4.035459e-06, 4.079427e-06, 4.062867e-06, 
    4.093295e-06, 4.099416e-06, 4.053198e-06, 4.081545e-06, 3.990906e-06, 
    4.005483e-06, 3.996801e-06, 3.965163e-06, 4.066679e-06, 4.014425e-06, 
    4.11117e-06, 4.082674e-06, 4.166107e-06, 4.124512e-06, 4.206405e-06, 
    4.241645e-06, 4.274944e-06, 4.314012e-06, 3.988905e-06, 3.977899e-06, 
    3.997616e-06, 4.024972e-06, 4.050436e-06, 4.084408e-06, 4.087893e-06, 
    4.094275e-06, 4.110829e-06, 4.124772e-06, 4.096293e-06, 4.128271e-06, 
    4.008866e-06, 4.07123e-06, 3.973742e-06, 4.002976e-06, 4.023357e-06, 
    4.014411e-06, 4.060976e-06, 4.071988e-06, 4.116886e-06, 4.093647e-06, 
    4.232934e-06, 4.171032e-06, 4.343875e-06, 4.295235e-06, 3.974057e-06, 
    3.988867e-06, 4.040618e-06, 4.015955e-06, 4.086682e-06, 4.104182e-06, 
    4.118435e-06, 4.136689e-06, 4.138663e-06, 4.149499e-06, 4.131749e-06, 
    4.148797e-06, 4.084481e-06, 4.113163e-06, 4.034687e-06, 4.05372e-06, 
    4.044959e-06, 4.035359e-06, 4.065023e-06, 4.09674e-06, 4.09742e-06, 
    4.107616e-06, 4.136412e-06, 4.08697e-06, 4.240953e-06, 4.145531e-06, 
    4.005047e-06, 4.033703e-06, 4.037805e-06, 4.026687e-06, 4.102426e-06, 
    4.074904e-06, 4.149235e-06, 4.129083e-06, 4.162127e-06, 4.145691e-06, 
    4.143275e-06, 4.122217e-06, 4.109132e-06, 4.076164e-06, 4.049434e-06, 
    4.028299e-06, 4.033209e-06, 4.056442e-06, 4.098685e-06, 4.138841e-06, 
    4.130029e-06, 4.159611e-06, 4.081533e-06, 4.114186e-06, 4.101551e-06, 
    4.134536e-06, 4.062427e-06, 4.12379e-06, 4.046812e-06, 4.053534e-06, 
    4.074359e-06, 4.116404e-06, 4.125736e-06, 4.135709e-06, 4.129554e-06, 
    4.09976e-06, 4.094889e-06, 4.073852e-06, 4.068053e-06, 4.05207e-06, 
    4.03886e-06, 4.050929e-06, 4.063621e-06, 4.099772e-06, 4.132484e-06, 
    4.16829e-06, 4.177076e-06, 4.219142e-06, 4.184885e-06, 4.241487e-06, 
    4.193339e-06, 4.276853e-06, 4.127362e-06, 4.191929e-06, 4.075308e-06, 
    4.087796e-06, 4.110429e-06, 4.162566e-06, 4.134381e-06, 4.167353e-06, 
    4.094698e-06, 4.057244e-06, 4.047582e-06, 4.029582e-06, 4.047994e-06, 
    4.046495e-06, 4.064148e-06, 4.058471e-06, 4.100976e-06, 4.078117e-06, 
    4.143214e-06, 4.167093e-06, 4.234886e-06, 4.276701e-06, 4.31947e-06, 
    4.338417e-06, 4.344191e-06, 4.346606e-06,
  4.133135e-06, 4.171723e-06, 4.164205e-06, 4.195447e-06, 4.178099e-06, 
    4.198581e-06, 4.140941e-06, 4.17326e-06, 4.152611e-06, 4.136599e-06, 
    4.256462e-06, 4.196844e-06, 4.318896e-06, 4.280498e-06, 4.377331e-06, 
    4.312909e-06, 4.390388e-06, 4.375463e-06, 4.420467e-06, 4.407547e-06, 
    4.465407e-06, 4.426438e-06, 4.495569e-06, 4.456082e-06, 4.462247e-06, 
    4.425156e-06, 4.208801e-06, 4.249014e-06, 4.206426e-06, 4.212145e-06, 
    4.209578e-06, 4.178458e-06, 4.162826e-06, 4.130193e-06, 4.136106e-06, 
    4.160079e-06, 4.214718e-06, 4.196123e-06, 4.243073e-06, 4.242009e-06, 
    4.294625e-06, 4.270856e-06, 4.35985e-06, 4.334448e-06, 4.408086e-06, 
    4.389499e-06, 4.407212e-06, 4.401837e-06, 4.407282e-06, 4.380041e-06, 
    4.391701e-06, 4.367774e-06, 4.275302e-06, 4.302361e-06, 4.221949e-06, 
    4.174021e-06, 4.142356e-06, 4.119971e-06, 4.123131e-06, 4.12916e-06, 
    4.16022e-06, 4.189542e-06, 4.211968e-06, 4.227008e-06, 4.241856e-06, 
    4.28699e-06, 4.310986e-06, 4.364998e-06, 4.35522e-06, 4.371791e-06, 
    4.387653e-06, 4.414361e-06, 4.409958e-06, 4.421749e-06, 4.371352e-06, 
    4.404809e-06, 4.349657e-06, 4.364701e-06, 4.245905e-06, 4.201135e-06, 
    4.182194e-06, 4.16565e-06, 4.125562e-06, 4.153223e-06, 4.142306e-06, 
    4.168302e-06, 4.18487e-06, 4.176671e-06, 4.22742e-06, 4.207649e-06, 
    4.31241e-06, 4.267104e-06, 4.385801e-06, 4.357226e-06, 4.392666e-06, 
    4.37456e-06, 4.40561e-06, 4.37766e-06, 4.426141e-06, 4.436741e-06, 
    4.429495e-06, 4.457359e-06, 4.376114e-06, 4.407213e-06, 4.176442e-06, 
    4.177778e-06, 4.184008e-06, 4.156665e-06, 4.154995e-06, 4.130031e-06, 
    4.152239e-06, 4.161717e-06, 4.185832e-06, 4.200134e-06, 4.213755e-06, 
    4.243793e-06, 4.277487e-06, 4.324857e-06, 4.359075e-06, 4.382099e-06, 
    4.367972e-06, 4.380443e-06, 4.366504e-06, 4.359979e-06, 4.432768e-06, 
    4.39181e-06, 4.453345e-06, 4.449927e-06, 4.42203e-06, 4.450312e-06, 
    4.178717e-06, 4.171028e-06, 4.144397e-06, 4.16523e-06, 4.127318e-06, 
    4.148515e-06, 4.160733e-06, 4.208062e-06, 4.218501e-06, 4.228195e-06, 
    4.247378e-06, 4.27207e-06, 4.315587e-06, 4.353656e-06, 4.388576e-06, 
    4.386012e-06, 4.386915e-06, 4.394737e-06, 4.375377e-06, 4.39792e-06, 
    4.401711e-06, 4.391804e-06, 4.44947e-06, 4.432951e-06, 4.449854e-06, 
    4.439094e-06, 4.173527e-06, 4.186473e-06, 4.179474e-06, 4.192641e-06, 
    4.183363e-06, 4.22471e-06, 4.237152e-06, 4.295649e-06, 4.271584e-06, 
    4.309918e-06, 4.275469e-06, 4.281561e-06, 4.311175e-06, 4.277326e-06, 
    4.351553e-06, 4.301151e-06, 4.395041e-06, 4.344421e-06, 4.398225e-06, 
    4.388425e-06, 4.404656e-06, 4.419223e-06, 4.43759e-06, 4.471593e-06, 
    4.463705e-06, 4.492228e-06, 4.205816e-06, 4.222687e-06, 4.2212e-06, 
    4.238893e-06, 4.252006e-06, 4.280506e-06, 4.326448e-06, 4.309139e-06, 
    4.340946e-06, 4.347348e-06, 4.299036e-06, 4.328663e-06, 4.234e-06, 
    4.249214e-06, 4.240151e-06, 4.207146e-06, 4.313125e-06, 4.258548e-06, 
    4.359642e-06, 4.329841e-06, 4.417145e-06, 4.373603e-06, 4.459367e-06, 
    4.496329e-06, 4.531272e-06, 4.572315e-06, 4.231911e-06, 4.220428e-06, 
    4.241e-06, 4.269558e-06, 4.296152e-06, 4.331656e-06, 4.335297e-06, 
    4.341971e-06, 4.359284e-06, 4.373871e-06, 4.344084e-06, 4.377533e-06, 
    4.252749e-06, 4.317881e-06, 4.216093e-06, 4.246598e-06, 4.267871e-06, 
    4.258531e-06, 4.307162e-06, 4.318671e-06, 4.365622e-06, 4.341314e-06, 
    4.487191e-06, 4.422306e-06, 4.603706e-06, 4.552585e-06, 4.216421e-06, 
    4.231871e-06, 4.285896e-06, 4.260141e-06, 4.334031e-06, 4.352332e-06, 
    4.367241e-06, 4.386345e-06, 4.388409e-06, 4.399753e-06, 4.381173e-06, 
    4.399018e-06, 4.331731e-06, 4.361726e-06, 4.2797e-06, 4.299582e-06, 
    4.290428e-06, 4.280402e-06, 4.311392e-06, 4.344552e-06, 4.34526e-06, 
    4.355925e-06, 4.386065e-06, 4.334332e-06, 4.49561e-06, 4.395609e-06, 
    4.248755e-06, 4.278676e-06, 4.282957e-06, 4.271346e-06, 4.350496e-06, 
    4.32172e-06, 4.399476e-06, 4.378382e-06, 4.412975e-06, 4.395766e-06, 
    4.393237e-06, 4.371198e-06, 4.35751e-06, 4.323038e-06, 4.295105e-06, 
    4.273029e-06, 4.278156e-06, 4.302427e-06, 4.346585e-06, 4.388597e-06, 
    4.379374e-06, 4.41034e-06, 4.328649e-06, 4.362797e-06, 4.349581e-06, 
    4.38409e-06, 4.30868e-06, 4.372854e-06, 4.292365e-06, 4.299387e-06, 
    4.32115e-06, 4.36512e-06, 4.37488e-06, 4.385319e-06, 4.378875e-06, 
    4.347708e-06, 4.342614e-06, 4.32062e-06, 4.31456e-06, 4.297857e-06, 
    4.284058e-06, 4.296665e-06, 4.309928e-06, 4.347721e-06, 4.381943e-06, 
    4.419431e-06, 4.428633e-06, 4.472728e-06, 4.436818e-06, 4.496171e-06, 
    4.445685e-06, 4.533286e-06, 4.376587e-06, 4.444201e-06, 4.322141e-06, 
    4.335196e-06, 4.358868e-06, 4.413439e-06, 4.383927e-06, 4.418452e-06, 
    4.342414e-06, 4.303267e-06, 4.293169e-06, 4.27437e-06, 4.293599e-06, 
    4.292033e-06, 4.310477e-06, 4.304545e-06, 4.348979e-06, 4.325078e-06, 
    4.393174e-06, 4.418178e-06, 4.489234e-06, 4.533121e-06, 4.578048e-06, 
    4.597965e-06, 4.604037e-06, 4.606577e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.778224, 5.778204, 5.778208, 5.778193, 5.778201, 5.778191, 5.77822, 
    5.778203, 5.778214, 5.778222, 5.778162, 5.778192, 5.778132, 5.778151, 
    5.778103, 5.778135, 5.778097, 5.778104, 5.778083, 5.778089, 5.778061, 
    5.77808, 5.778047, 5.778066, 5.778063, 5.77808, 5.778186, 5.778166, 
    5.778187, 5.778184, 5.778185, 5.778201, 5.778209, 5.778225, 5.778222, 
    5.77821, 5.778183, 5.778192, 5.778169, 5.77817, 5.778144, 5.778155, 
    5.778112, 5.778124, 5.778089, 5.778098, 5.778089, 5.778091, 5.778089, 
    5.778102, 5.778097, 5.778108, 5.778153, 5.77814, 5.77818, 5.778203, 
    5.778219, 5.77823, 5.778229, 5.778225, 5.77821, 5.778195, 5.778184, 
    5.778177, 5.77817, 5.778148, 5.778136, 5.77811, 5.778114, 5.778106, 
    5.778099, 5.778086, 5.778088, 5.778082, 5.778106, 5.77809, 5.778117, 
    5.77811, 5.778168, 5.77819, 5.778199, 5.778207, 5.778227, 5.778214, 
    5.778219, 5.778206, 5.778198, 5.778202, 5.778177, 5.778186, 5.778135, 
    5.778157, 5.7781, 5.778113, 5.778096, 5.778105, 5.77809, 5.778103, 
    5.77808, 5.778075, 5.778078, 5.778065, 5.778104, 5.778089, 5.778202, 
    5.778202, 5.778198, 5.778212, 5.778213, 5.778225, 5.778214, 5.778209, 
    5.778197, 5.77819, 5.778183, 5.778169, 5.778152, 5.778129, 5.778112, 
    5.778101, 5.778108, 5.778102, 5.778109, 5.778112, 5.778077, 5.778097, 
    5.778067, 5.778069, 5.778082, 5.778069, 5.778201, 5.778205, 5.778218, 
    5.778208, 5.778226, 5.778216, 5.77821, 5.778186, 5.778181, 5.778176, 
    5.778167, 5.778155, 5.778133, 5.778115, 5.778098, 5.778099, 5.778099, 
    5.778095, 5.778104, 5.778093, 5.778092, 5.778097, 5.778069, 5.778077, 
    5.778069, 5.778074, 5.778203, 5.778197, 5.778201, 5.778194, 5.778199, 
    5.778178, 5.778172, 5.778143, 5.778155, 5.778136, 5.778153, 5.77815, 
    5.778136, 5.778152, 5.778116, 5.778141, 5.778095, 5.77812, 5.778093, 
    5.778098, 5.77809, 5.778083, 5.778074, 5.778058, 5.778062, 5.778049, 
    5.778187, 5.778179, 5.77818, 5.778171, 5.778165, 5.778151, 5.778128, 
    5.778137, 5.778121, 5.778118, 5.778141, 5.778127, 5.778173, 5.778166, 
    5.778171, 5.778187, 5.778135, 5.778162, 5.778112, 5.778127, 5.778084, 
    5.778105, 5.778064, 5.778046, 5.77803, 5.77801, 5.778174, 5.77818, 
    5.77817, 5.778156, 5.778143, 5.778126, 5.778124, 5.778121, 5.778112, 
    5.778105, 5.77812, 5.778103, 5.778164, 5.778132, 5.778183, 5.778167, 
    5.778157, 5.778162, 5.778138, 5.778132, 5.778109, 5.778121, 5.778051, 
    5.778082, 5.777996, 5.778019, 5.778182, 5.778174, 5.778148, 5.778161, 
    5.778124, 5.778116, 5.778109, 5.778099, 5.778098, 5.778093, 5.778101, 
    5.778093, 5.778126, 5.778111, 5.778151, 5.778141, 5.778146, 5.778151, 
    5.778136, 5.77812, 5.778119, 5.778114, 5.778099, 5.778124, 5.778047, 
    5.778095, 5.778166, 5.778152, 5.77815, 5.778155, 5.778117, 5.778131, 
    5.778093, 5.778103, 5.778086, 5.778095, 5.778096, 5.778106, 5.778113, 
    5.77813, 5.778143, 5.778154, 5.778152, 5.77814, 5.778119, 5.778098, 
    5.778102, 5.778088, 5.778127, 5.778111, 5.778117, 5.7781, 5.778137, 
    5.778106, 5.778145, 5.778141, 5.778131, 5.77811, 5.778105, 5.7781, 
    5.778103, 5.778118, 5.778121, 5.778131, 5.778134, 5.778142, 5.778149, 
    5.778143, 5.778136, 5.778118, 5.778101, 5.778083, 5.778079, 5.778058, 
    5.778075, 5.778047, 5.77807, 5.778029, 5.778104, 5.778071, 5.778131, 
    5.778124, 5.778112, 5.778086, 5.7781, 5.778084, 5.778121, 5.77814, 
    5.778144, 5.778154, 5.778144, 5.778145, 5.778136, 5.778139, 5.778117, 
    5.778129, 5.778096, 5.778084, 5.778049, 5.778029, 5.778008, 5.777998, 
    5.777995, 5.777994 ;

 SOIL1C_TO_SOIL2C =
  3.109261e-08, 3.122964e-08, 3.1203e-08, 3.131352e-08, 3.125221e-08, 
    3.132458e-08, 3.112039e-08, 3.123507e-08, 3.116186e-08, 3.110495e-08, 
    3.152799e-08, 3.131845e-08, 3.17457e-08, 3.161205e-08, 3.194781e-08, 
    3.172489e-08, 3.199276e-08, 3.194139e-08, 3.209603e-08, 3.205173e-08, 
    3.224952e-08, 3.211647e-08, 3.235206e-08, 3.221775e-08, 3.223876e-08, 
    3.211208e-08, 3.136062e-08, 3.15019e-08, 3.135225e-08, 3.13724e-08, 
    3.136336e-08, 3.125347e-08, 3.11981e-08, 3.108214e-08, 3.110319e-08, 
    3.118836e-08, 3.138146e-08, 3.131591e-08, 3.148111e-08, 3.147738e-08, 
    3.16613e-08, 3.157838e-08, 3.188752e-08, 3.179966e-08, 3.205357e-08, 
    3.198971e-08, 3.205057e-08, 3.203212e-08, 3.205081e-08, 3.195716e-08, 
    3.199728e-08, 3.191488e-08, 3.159391e-08, 3.168823e-08, 3.140691e-08, 
    3.123775e-08, 3.112542e-08, 3.10457e-08, 3.105697e-08, 3.107846e-08, 
    3.118886e-08, 3.129267e-08, 3.137178e-08, 3.14247e-08, 3.147685e-08, 
    3.163467e-08, 3.171822e-08, 3.190529e-08, 3.187153e-08, 3.192872e-08, 
    3.198336e-08, 3.207509e-08, 3.206e-08, 3.210041e-08, 3.192721e-08, 
    3.204232e-08, 3.185231e-08, 3.190427e-08, 3.1491e-08, 3.13336e-08, 
    3.126668e-08, 3.120812e-08, 3.106564e-08, 3.116403e-08, 3.112524e-08, 
    3.121752e-08, 3.127616e-08, 3.124716e-08, 3.142615e-08, 3.135656e-08, 
    3.172317e-08, 3.156526e-08, 3.197699e-08, 3.187846e-08, 3.200061e-08, 
    3.193828e-08, 3.204507e-08, 3.194896e-08, 3.211546e-08, 3.215172e-08, 
    3.212693e-08, 3.222211e-08, 3.194363e-08, 3.205057e-08, 3.124635e-08, 
    3.125108e-08, 3.127311e-08, 3.117625e-08, 3.117032e-08, 3.108156e-08, 
    3.116055e-08, 3.119418e-08, 3.127956e-08, 3.133006e-08, 3.137808e-08, 
    3.148364e-08, 3.160153e-08, 3.176639e-08, 3.188485e-08, 3.196425e-08, 
    3.191556e-08, 3.195855e-08, 3.19105e-08, 3.188797e-08, 3.213813e-08, 
    3.199766e-08, 3.220843e-08, 3.219677e-08, 3.210137e-08, 3.219808e-08, 
    3.12544e-08, 3.122718e-08, 3.113268e-08, 3.120664e-08, 3.10719e-08, 
    3.114732e-08, 3.119068e-08, 3.135801e-08, 3.139478e-08, 3.142888e-08, 
    3.149621e-08, 3.158262e-08, 3.173421e-08, 3.186612e-08, 3.198654e-08, 
    3.197772e-08, 3.198083e-08, 3.200772e-08, 3.194109e-08, 3.201867e-08, 
    3.203168e-08, 3.199764e-08, 3.21952e-08, 3.213876e-08, 3.219652e-08, 
    3.215977e-08, 3.123603e-08, 3.128183e-08, 3.125708e-08, 3.130361e-08, 
    3.127083e-08, 3.141661e-08, 3.146032e-08, 3.166486e-08, 3.158092e-08, 
    3.171451e-08, 3.159449e-08, 3.161576e-08, 3.171886e-08, 3.160098e-08, 
    3.185884e-08, 3.168401e-08, 3.200877e-08, 3.183417e-08, 3.201971e-08, 
    3.198602e-08, 3.20418e-08, 3.209176e-08, 3.215463e-08, 3.22706e-08, 
    3.224374e-08, 3.234073e-08, 3.13501e-08, 3.140951e-08, 3.140428e-08, 
    3.146645e-08, 3.151242e-08, 3.161208e-08, 3.177192e-08, 3.171181e-08, 
    3.182216e-08, 3.184432e-08, 3.167667e-08, 3.17796e-08, 3.144926e-08, 
    3.150263e-08, 3.147086e-08, 3.135479e-08, 3.172566e-08, 3.153532e-08, 
    3.18868e-08, 3.178369e-08, 3.208464e-08, 3.193496e-08, 3.222896e-08, 
    3.235462e-08, 3.247292e-08, 3.261115e-08, 3.144193e-08, 3.140157e-08, 
    3.147384e-08, 3.157383e-08, 3.166662e-08, 3.178998e-08, 3.18026e-08, 
    3.182571e-08, 3.188557e-08, 3.19359e-08, 3.183301e-08, 3.194852e-08, 
    3.151499e-08, 3.174218e-08, 3.13863e-08, 3.149346e-08, 3.156794e-08, 
    3.153527e-08, 3.170495e-08, 3.174494e-08, 3.190744e-08, 3.182344e-08, 
    3.232361e-08, 3.210231e-08, 3.271641e-08, 3.254479e-08, 3.138747e-08, 
    3.144179e-08, 3.163088e-08, 3.154091e-08, 3.179821e-08, 3.186155e-08, 
    3.191304e-08, 3.197886e-08, 3.198597e-08, 3.202496e-08, 3.196106e-08, 
    3.202244e-08, 3.179024e-08, 3.1894e-08, 3.160927e-08, 3.167857e-08, 
    3.164669e-08, 3.161172e-08, 3.171965e-08, 3.183463e-08, 3.183709e-08, 
    3.187396e-08, 3.197784e-08, 3.179926e-08, 3.235215e-08, 3.201067e-08, 
    3.150103e-08, 3.160568e-08, 3.162063e-08, 3.158009e-08, 3.18552e-08, 
    3.175552e-08, 3.202401e-08, 3.195145e-08, 3.207035e-08, 3.201126e-08, 
    3.200257e-08, 3.192669e-08, 3.187944e-08, 3.176008e-08, 3.166297e-08, 
    3.158598e-08, 3.160388e-08, 3.168847e-08, 3.184167e-08, 3.198661e-08, 
    3.195485e-08, 3.206131e-08, 3.177956e-08, 3.18977e-08, 3.185203e-08, 
    3.19711e-08, 3.171021e-08, 3.193235e-08, 3.165344e-08, 3.167789e-08, 
    3.175354e-08, 3.19057e-08, 3.193938e-08, 3.197533e-08, 3.195315e-08, 
    3.184556e-08, 3.182793e-08, 3.17517e-08, 3.173065e-08, 3.167257e-08, 
    3.162448e-08, 3.166841e-08, 3.171455e-08, 3.18456e-08, 3.19637e-08, 
    3.209247e-08, 3.212399e-08, 3.227443e-08, 3.215196e-08, 3.235405e-08, 
    3.218222e-08, 3.247968e-08, 3.194523e-08, 3.217718e-08, 3.175698e-08, 
    3.180225e-08, 3.188412e-08, 3.207192e-08, 3.197054e-08, 3.20891e-08, 
    3.182724e-08, 3.169138e-08, 3.165623e-08, 3.159066e-08, 3.165773e-08, 
    3.165228e-08, 3.171647e-08, 3.169584e-08, 3.184995e-08, 3.176717e-08, 
    3.200235e-08, 3.208817e-08, 3.233056e-08, 3.247915e-08, 3.263042e-08, 
    3.26972e-08, 3.271753e-08, 3.272602e-08 ;

 SOIL1C_TO_SOIL3C =
  3.687849e-10, 3.704106e-10, 3.700946e-10, 3.714059e-10, 3.706785e-10, 
    3.715372e-10, 3.691145e-10, 3.704752e-10, 3.696066e-10, 3.689313e-10, 
    3.739507e-10, 3.714644e-10, 3.765339e-10, 3.74948e-10, 3.78932e-10, 
    3.762871e-10, 3.794654e-10, 3.788558e-10, 3.806907e-10, 3.801651e-10, 
    3.82512e-10, 3.809334e-10, 3.837288e-10, 3.821351e-10, 3.823844e-10, 
    3.808813e-10, 3.719648e-10, 3.736411e-10, 3.718655e-10, 3.721045e-10, 
    3.719973e-10, 3.706935e-10, 3.700365e-10, 3.686607e-10, 3.689105e-10, 
    3.69921e-10, 3.72212e-10, 3.714344e-10, 3.733945e-10, 3.733502e-10, 
    3.755325e-10, 3.745486e-10, 3.782167e-10, 3.771741e-10, 3.80187e-10, 
    3.794293e-10, 3.801514e-10, 3.799324e-10, 3.801542e-10, 3.79043e-10, 
    3.795191e-10, 3.785412e-10, 3.747328e-10, 3.75852e-10, 3.72514e-10, 
    3.70507e-10, 3.691742e-10, 3.682284e-10, 3.683621e-10, 3.686169e-10, 
    3.699269e-10, 3.711586e-10, 3.720973e-10, 3.727252e-10, 3.733439e-10, 
    3.752164e-10, 3.762078e-10, 3.784275e-10, 3.780269e-10, 3.787055e-10, 
    3.793539e-10, 3.804423e-10, 3.802632e-10, 3.807427e-10, 3.786877e-10, 
    3.800534e-10, 3.777988e-10, 3.784154e-10, 3.735118e-10, 3.716442e-10, 
    3.708502e-10, 3.701554e-10, 3.684649e-10, 3.696323e-10, 3.691721e-10, 
    3.70267e-10, 3.709627e-10, 3.706186e-10, 3.727423e-10, 3.719167e-10, 
    3.762665e-10, 3.743929e-10, 3.792782e-10, 3.781092e-10, 3.795585e-10, 
    3.788189e-10, 3.800861e-10, 3.789457e-10, 3.809213e-10, 3.813515e-10, 
    3.810575e-10, 3.821869e-10, 3.788825e-10, 3.801514e-10, 3.70609e-10, 
    3.706651e-10, 3.709265e-10, 3.697772e-10, 3.697069e-10, 3.686538e-10, 
    3.695909e-10, 3.6999e-10, 3.710031e-10, 3.716023e-10, 3.721719e-10, 
    3.734244e-10, 3.748232e-10, 3.767794e-10, 3.78185e-10, 3.791271e-10, 
    3.785494e-10, 3.790594e-10, 3.784893e-10, 3.78222e-10, 3.811903e-10, 
    3.795235e-10, 3.820245e-10, 3.818861e-10, 3.807542e-10, 3.819017e-10, 
    3.707045e-10, 3.703816e-10, 3.692603e-10, 3.701378e-10, 3.685391e-10, 
    3.694339e-10, 3.699484e-10, 3.719339e-10, 3.723702e-10, 3.727746e-10, 
    3.735736e-10, 3.745989e-10, 3.763976e-10, 3.779627e-10, 3.793916e-10, 
    3.792869e-10, 3.793238e-10, 3.79643e-10, 3.788523e-10, 3.797728e-10, 
    3.799272e-10, 3.795233e-10, 3.818675e-10, 3.811979e-10, 3.818831e-10, 
    3.814471e-10, 3.704865e-10, 3.710299e-10, 3.707363e-10, 3.712884e-10, 
    3.708994e-10, 3.726291e-10, 3.731478e-10, 3.755747e-10, 3.745787e-10, 
    3.761639e-10, 3.747397e-10, 3.749921e-10, 3.762154e-10, 3.748167e-10, 
    3.778764e-10, 3.758019e-10, 3.796554e-10, 3.775835e-10, 3.797852e-10, 
    3.793854e-10, 3.800473e-10, 3.806401e-10, 3.813861e-10, 3.827621e-10, 
    3.824435e-10, 3.835944e-10, 3.7184e-10, 3.725448e-10, 3.724829e-10, 
    3.732205e-10, 3.73766e-10, 3.749485e-10, 3.76845e-10, 3.761318e-10, 
    3.774412e-10, 3.77704e-10, 3.757148e-10, 3.769361e-10, 3.730166e-10, 
    3.736498e-10, 3.732728e-10, 3.718956e-10, 3.762961e-10, 3.740377e-10, 
    3.782082e-10, 3.769846e-10, 3.805556e-10, 3.787796e-10, 3.822681e-10, 
    3.837592e-10, 3.85163e-10, 3.868032e-10, 3.729295e-10, 3.724507e-10, 
    3.733082e-10, 3.744946e-10, 3.755956e-10, 3.770592e-10, 3.77209e-10, 
    3.774832e-10, 3.781935e-10, 3.787907e-10, 3.775699e-10, 3.789405e-10, 
    3.737965e-10, 3.764921e-10, 3.722695e-10, 3.735409e-10, 3.744247e-10, 
    3.740371e-10, 3.760503e-10, 3.765248e-10, 3.78453e-10, 3.774563e-10, 
    3.833912e-10, 3.807653e-10, 3.880523e-10, 3.860157e-10, 3.722833e-10, 
    3.729279e-10, 3.751714e-10, 3.74104e-10, 3.77157e-10, 3.779085e-10, 
    3.785195e-10, 3.793004e-10, 3.793848e-10, 3.798475e-10, 3.790892e-10, 
    3.798176e-10, 3.770624e-10, 3.782936e-10, 3.749151e-10, 3.757373e-10, 
    3.753591e-10, 3.749441e-10, 3.762248e-10, 3.775891e-10, 3.776183e-10, 
    3.780558e-10, 3.792884e-10, 3.771694e-10, 3.837299e-10, 3.79678e-10, 
    3.736309e-10, 3.748724e-10, 3.750499e-10, 3.745689e-10, 3.778332e-10, 
    3.766503e-10, 3.798362e-10, 3.789752e-10, 3.80386e-10, 3.79685e-10, 
    3.795818e-10, 3.786814e-10, 3.781208e-10, 3.767046e-10, 3.755523e-10, 
    3.746387e-10, 3.748511e-10, 3.758548e-10, 3.776726e-10, 3.793924e-10, 
    3.790156e-10, 3.802788e-10, 3.769356e-10, 3.783374e-10, 3.777956e-10, 
    3.792084e-10, 3.761129e-10, 3.787486e-10, 3.754391e-10, 3.757293e-10, 
    3.766269e-10, 3.784324e-10, 3.78832e-10, 3.792585e-10, 3.789954e-10, 
    3.777187e-10, 3.775096e-10, 3.766051e-10, 3.763553e-10, 3.756661e-10, 
    3.750955e-10, 3.756168e-10, 3.761643e-10, 3.777193e-10, 3.791206e-10, 
    3.806485e-10, 3.810225e-10, 3.828077e-10, 3.813544e-10, 3.837524e-10, 
    3.817135e-10, 3.852432e-10, 3.789015e-10, 3.816537e-10, 3.766678e-10, 
    3.772049e-10, 3.781763e-10, 3.804047e-10, 3.792018e-10, 3.806086e-10, 
    3.775014e-10, 3.758893e-10, 3.754723e-10, 3.746942e-10, 3.754901e-10, 
    3.754254e-10, 3.761871e-10, 3.759423e-10, 3.777709e-10, 3.767887e-10, 
    3.795792e-10, 3.805975e-10, 3.834737e-10, 3.852369e-10, 3.870319e-10, 
    3.878243e-10, 3.880655e-10, 3.881664e-10 ;

 SOIL1C_vr =
  19.98093, 19.98088, 19.98089, 19.98085, 19.98087, 19.98085, 19.98092, 
    19.98088, 19.98091, 19.98093, 19.98077, 19.98085, 19.98069, 19.98074, 
    19.98061, 19.98069, 19.98059, 19.98061, 19.98055, 19.98057, 19.9805, 
    19.98055, 19.98046, 19.98051, 19.9805, 19.98055, 19.98083, 19.98078, 
    19.98083, 19.98083, 19.98083, 19.98087, 19.98089, 19.98094, 19.98093, 
    19.9809, 19.98082, 19.98085, 19.98079, 19.98079, 19.98072, 19.98075, 
    19.98063, 19.98067, 19.98057, 19.98059, 19.98057, 19.98058, 19.98057, 
    19.98061, 19.98059, 19.98062, 19.98074, 19.98071, 19.98081, 19.98088, 
    19.98092, 19.98095, 19.98095, 19.98094, 19.9809, 19.98086, 19.98083, 
    19.98081, 19.98079, 19.98073, 19.9807, 19.98063, 19.98064, 19.98062, 
    19.9806, 19.98056, 19.98057, 19.98055, 19.98062, 19.98057, 19.98065, 
    19.98063, 19.98078, 19.98084, 19.98087, 19.98089, 19.98094, 19.98091, 
    19.98092, 19.98089, 19.98086, 19.98088, 19.98081, 19.98083, 19.98069, 
    19.98075, 19.9806, 19.98064, 19.98059, 19.98061, 19.98057, 19.98061, 
    19.98055, 19.98053, 19.98054, 19.98051, 19.98061, 19.98057, 19.98088, 
    19.98087, 19.98087, 19.9809, 19.9809, 19.98094, 19.98091, 19.9809, 
    19.98086, 19.98084, 19.98083, 19.98079, 19.98074, 19.98068, 19.98063, 
    19.9806, 19.98062, 19.98061, 19.98062, 19.98063, 19.98054, 19.98059, 
    19.98051, 19.98052, 19.98055, 19.98051, 19.98087, 19.98088, 19.98092, 
    19.98089, 19.98094, 19.98091, 19.9809, 19.98083, 19.98082, 19.98081, 
    19.98078, 19.98075, 19.98069, 19.98064, 19.98059, 19.9806, 19.9806, 
    19.98059, 19.98061, 19.98058, 19.98058, 19.98059, 19.98052, 19.98054, 
    19.98052, 19.98053, 19.98088, 19.98086, 19.98087, 19.98085, 19.98087, 
    19.98081, 19.98079, 19.98072, 19.98075, 19.9807, 19.98074, 19.98074, 
    19.9807, 19.98074, 19.98064, 19.98071, 19.98059, 19.98065, 19.98058, 
    19.98059, 19.98057, 19.98055, 19.98053, 19.98049, 19.9805, 19.98046, 
    19.98083, 19.98081, 19.98082, 19.98079, 19.98077, 19.98074, 19.98068, 
    19.9807, 19.98066, 19.98065, 19.98071, 19.98067, 19.9808, 19.98078, 
    19.98079, 19.98083, 19.98069, 19.98077, 19.98063, 19.98067, 19.98056, 
    19.98061, 19.9805, 19.98046, 19.98041, 19.98036, 19.9808, 19.98082, 
    19.98079, 19.98075, 19.98072, 19.98067, 19.98067, 19.98066, 19.98063, 
    19.98061, 19.98065, 19.98061, 19.98077, 19.98069, 19.98082, 19.98078, 
    19.98075, 19.98077, 19.9807, 19.98069, 19.98063, 19.98066, 19.98047, 
    19.98055, 19.98032, 19.98038, 19.98082, 19.9808, 19.98073, 19.98076, 
    19.98067, 19.98064, 19.98062, 19.9806, 19.98059, 19.98058, 19.9806, 
    19.98058, 19.98067, 19.98063, 19.98074, 19.98071, 19.98072, 19.98074, 
    19.9807, 19.98065, 19.98065, 19.98064, 19.9806, 19.98067, 19.98046, 
    19.98059, 19.98078, 19.98074, 19.98073, 19.98075, 19.98064, 19.98068, 
    19.98058, 19.98061, 19.98056, 19.98059, 19.98059, 19.98062, 19.98063, 
    19.98068, 19.98072, 19.98075, 19.98074, 19.98071, 19.98065, 19.98059, 
    19.98061, 19.98057, 19.98067, 19.98063, 19.98065, 19.9806, 19.9807, 
    19.98062, 19.98072, 19.98071, 19.98068, 19.98063, 19.98061, 19.9806, 
    19.98061, 19.98065, 19.98066, 19.98068, 19.98069, 19.98071, 19.98073, 
    19.98071, 19.9807, 19.98065, 19.9806, 19.98055, 19.98054, 19.98049, 
    19.98053, 19.98046, 19.98052, 19.98041, 19.98061, 19.98052, 19.98068, 
    19.98067, 19.98063, 19.98056, 19.9806, 19.98056, 19.98066, 19.98071, 
    19.98072, 19.98075, 19.98072, 19.98072, 19.9807, 19.98071, 19.98065, 
    19.98068, 19.98059, 19.98056, 19.98046, 19.98041, 19.98035, 19.98033, 
    19.98032, 19.98032,
  19.98316, 19.98309, 19.9831, 19.98305, 19.98308, 19.98305, 19.98314, 
    19.98309, 19.98312, 19.98315, 19.98295, 19.98305, 19.98285, 19.98291, 
    19.98276, 19.98286, 19.98273, 19.98276, 19.98269, 19.98271, 19.98262, 
    19.98268, 19.98257, 19.98263, 19.98262, 19.98268, 19.98303, 19.98296, 
    19.98303, 19.98302, 19.98303, 19.98308, 19.98311, 19.98316, 19.98315, 
    19.98311, 19.98302, 19.98305, 19.98298, 19.98298, 19.98289, 19.98293, 
    19.98278, 19.98283, 19.98271, 19.98274, 19.98271, 19.98272, 19.98271, 
    19.98275, 19.98273, 19.98277, 19.98292, 19.98288, 19.98301, 19.98309, 
    19.98314, 19.98318, 19.98317, 19.98316, 19.98311, 19.98306, 19.98302, 
    19.983, 19.98298, 19.9829, 19.98286, 19.98278, 19.98279, 19.98277, 
    19.98274, 19.9827, 19.9827, 19.98269, 19.98277, 19.98271, 19.9828, 
    19.98278, 19.98297, 19.98304, 19.98307, 19.9831, 19.98317, 19.98312, 
    19.98314, 19.9831, 19.98307, 19.98308, 19.983, 19.98303, 19.98286, 
    19.98293, 19.98274, 19.98279, 19.98273, 19.98276, 19.98271, 19.98276, 
    19.98268, 19.98266, 19.98267, 19.98263, 19.98276, 19.98271, 19.98308, 
    19.98308, 19.98307, 19.98312, 19.98312, 19.98316, 19.98312, 19.98311, 
    19.98307, 19.98305, 19.98302, 19.98297, 19.98292, 19.98284, 19.98279, 
    19.98275, 19.98277, 19.98275, 19.98277, 19.98278, 19.98267, 19.98273, 
    19.98264, 19.98264, 19.98269, 19.98264, 19.98308, 19.98309, 19.98314, 
    19.9831, 19.98317, 19.98313, 19.98311, 19.98303, 19.98302, 19.983, 
    19.98297, 19.98293, 19.98286, 19.98279, 19.98274, 19.98274, 19.98274, 
    19.98273, 19.98276, 19.98272, 19.98272, 19.98273, 19.98264, 19.98267, 
    19.98264, 19.98266, 19.98309, 19.98307, 19.98308, 19.98306, 19.98307, 
    19.983, 19.98298, 19.98289, 19.98293, 19.98286, 19.98292, 19.98291, 
    19.98286, 19.98292, 19.9828, 19.98288, 19.98273, 19.98281, 19.98272, 
    19.98274, 19.98271, 19.98269, 19.98266, 19.9826, 19.98262, 19.98257, 
    19.98304, 19.98301, 19.98301, 19.98298, 19.98296, 19.98291, 19.98284, 
    19.98287, 19.98281, 19.98281, 19.98288, 19.98283, 19.98299, 19.98296, 
    19.98298, 19.98303, 19.98286, 19.98295, 19.98278, 19.98283, 19.98269, 
    19.98276, 19.98263, 19.98257, 19.98251, 19.98245, 19.98299, 19.98301, 
    19.98298, 19.98293, 19.98289, 19.98283, 19.98282, 19.98281, 19.98278, 
    19.98276, 19.98281, 19.98276, 19.98296, 19.98285, 19.98302, 19.98297, 
    19.98293, 19.98295, 19.98287, 19.98285, 19.98277, 19.98281, 19.98258, 
    19.98269, 19.9824, 19.98248, 19.98302, 19.98299, 19.9829, 19.98295, 
    19.98283, 19.9828, 19.98277, 19.98274, 19.98274, 19.98272, 19.98275, 
    19.98272, 19.98283, 19.98278, 19.98291, 19.98288, 19.9829, 19.98291, 
    19.98286, 19.98281, 19.98281, 19.98279, 19.98274, 19.98283, 19.98257, 
    19.98273, 19.98297, 19.98292, 19.98291, 19.98293, 19.9828, 19.98285, 
    19.98272, 19.98275, 19.9827, 19.98273, 19.98273, 19.98277, 19.98279, 
    19.98284, 19.98289, 19.98293, 19.98292, 19.98288, 19.98281, 19.98274, 
    19.98275, 19.9827, 19.98283, 19.98278, 19.9828, 19.98275, 19.98287, 
    19.98276, 19.98289, 19.98288, 19.98285, 19.98278, 19.98276, 19.98274, 
    19.98275, 19.9828, 19.98281, 19.98285, 19.98286, 19.98289, 19.98291, 
    19.98289, 19.98286, 19.9828, 19.98275, 19.98269, 19.98267, 19.9826, 
    19.98266, 19.98257, 19.98265, 19.98251, 19.98276, 19.98265, 19.98285, 
    19.98282, 19.98279, 19.9827, 19.98275, 19.98269, 19.98281, 19.98288, 
    19.98289, 19.98292, 19.98289, 19.98289, 19.98286, 19.98287, 19.9828, 
    19.98284, 19.98273, 19.98269, 19.98258, 19.98251, 19.98244, 19.98241, 
    19.9824, 19.98239,
  19.98417, 19.9841, 19.98411, 19.98406, 19.98409, 19.98405, 19.98416, 
    19.9841, 19.98413, 19.98417, 19.98395, 19.98405, 19.98384, 19.98391, 
    19.98373, 19.98385, 19.98371, 19.98374, 19.98366, 19.98368, 19.98358, 
    19.98365, 19.98353, 19.9836, 19.98359, 19.98365, 19.98403, 19.98396, 
    19.98404, 19.98403, 19.98403, 19.98409, 19.98412, 19.98418, 19.98417, 
    19.98412, 19.98402, 19.98406, 19.98397, 19.98397, 19.98388, 19.98392, 
    19.98376, 19.98381, 19.98368, 19.98371, 19.98368, 19.98369, 19.98368, 
    19.98373, 19.98371, 19.98375, 19.98392, 19.98387, 19.98401, 19.9841, 
    19.98415, 19.9842, 19.98419, 19.98418, 19.98412, 19.98407, 19.98403, 
    19.984, 19.98397, 19.98389, 19.98385, 19.98376, 19.98377, 19.98374, 
    19.98372, 19.98367, 19.98368, 19.98366, 19.98374, 19.98369, 19.98378, 
    19.98376, 19.98397, 19.98405, 19.98408, 19.98411, 19.98418, 19.98413, 
    19.98415, 19.98411, 19.98408, 19.98409, 19.984, 19.98404, 19.98385, 
    19.98393, 19.98372, 19.98377, 19.98371, 19.98374, 19.98368, 19.98373, 
    19.98365, 19.98363, 19.98364, 19.98359, 19.98374, 19.98368, 19.98409, 
    19.98409, 19.98408, 19.98413, 19.98413, 19.98418, 19.98414, 19.98412, 
    19.98408, 19.98405, 19.98402, 19.98397, 19.98391, 19.98383, 19.98377, 
    19.98372, 19.98375, 19.98373, 19.98375, 19.98376, 19.98364, 19.98371, 
    19.9836, 19.98361, 19.98366, 19.98361, 19.98409, 19.9841, 19.98415, 
    19.98411, 19.98418, 19.98414, 19.98412, 19.98404, 19.98402, 19.984, 
    19.98396, 19.98392, 19.98384, 19.98378, 19.98371, 19.98372, 19.98372, 
    19.9837, 19.98374, 19.9837, 19.98369, 19.98371, 19.98361, 19.98364, 
    19.98361, 19.98363, 19.9841, 19.98407, 19.98409, 19.98406, 19.98408, 
    19.984, 19.98398, 19.98388, 19.98392, 19.98385, 19.98391, 19.9839, 
    19.98385, 19.98391, 19.98378, 19.98387, 19.9837, 19.98379, 19.9837, 
    19.98372, 19.98369, 19.98366, 19.98363, 19.98357, 19.98358, 19.98353, 
    19.98404, 19.98401, 19.98401, 19.98398, 19.98396, 19.98391, 19.98382, 
    19.98385, 19.9838, 19.98379, 19.98387, 19.98382, 19.98399, 19.98396, 
    19.98398, 19.98404, 19.98385, 19.98394, 19.98376, 19.98382, 19.98366, 
    19.98374, 19.98359, 19.98353, 19.98347, 19.9834, 19.98399, 19.98401, 
    19.98398, 19.98392, 19.98388, 19.98381, 19.98381, 19.9838, 19.98376, 
    19.98374, 19.98379, 19.98373, 19.98396, 19.98384, 19.98402, 19.98397, 
    19.98393, 19.98394, 19.98386, 19.98384, 19.98376, 19.9838, 19.98354, 
    19.98366, 19.98334, 19.98343, 19.98402, 19.98399, 19.9839, 19.98394, 
    19.98381, 19.98378, 19.98375, 19.98372, 19.98372, 19.98369, 19.98373, 
    19.9837, 19.98381, 19.98376, 19.98391, 19.98387, 19.98389, 19.98391, 
    19.98385, 19.98379, 19.98379, 19.98377, 19.98372, 19.98381, 19.98353, 
    19.9837, 19.98396, 19.98391, 19.9839, 19.98392, 19.98378, 19.98383, 
    19.98369, 19.98373, 19.98367, 19.9837, 19.98371, 19.98374, 19.98377, 
    19.98383, 19.98388, 19.98392, 19.98391, 19.98387, 19.98379, 19.98371, 
    19.98373, 19.98368, 19.98382, 19.98376, 19.98378, 19.98372, 19.98385, 
    19.98374, 19.98388, 19.98387, 19.98383, 19.98376, 19.98374, 19.98372, 
    19.98373, 19.98379, 19.9838, 19.98383, 19.98384, 19.98388, 19.9839, 
    19.98388, 19.98385, 19.98379, 19.98373, 19.98366, 19.98364, 19.98357, 
    19.98363, 19.98353, 19.98361, 19.98346, 19.98374, 19.98362, 19.98383, 
    19.98381, 19.98377, 19.98367, 19.98372, 19.98366, 19.9838, 19.98386, 
    19.98388, 19.98392, 19.98388, 19.98388, 19.98385, 19.98386, 19.98378, 
    19.98383, 19.98371, 19.98366, 19.98354, 19.98346, 19.98339, 19.98335, 
    19.98334, 19.98334,
  19.98496, 19.98489, 19.9849, 19.98484, 19.98487, 19.98484, 19.98494, 
    19.98488, 19.98492, 19.98495, 19.98473, 19.98484, 19.98462, 19.98469, 
    19.98451, 19.98463, 19.98449, 19.98451, 19.98443, 19.98446, 19.98435, 
    19.98442, 19.9843, 19.98437, 19.98436, 19.98443, 19.98482, 19.98474, 
    19.98482, 19.98481, 19.98482, 19.98487, 19.9849, 19.98496, 19.98495, 
    19.98491, 19.98481, 19.98484, 19.98475, 19.98476, 19.98466, 19.9847, 
    19.98454, 19.98459, 19.98446, 19.98449, 19.98446, 19.98447, 19.98446, 
    19.98451, 19.98449, 19.98453, 19.9847, 19.98465, 19.98479, 19.98488, 
    19.98494, 19.98498, 19.98498, 19.98496, 19.98491, 19.98485, 19.98481, 
    19.98478, 19.98476, 19.98467, 19.98463, 19.98453, 19.98455, 19.98452, 
    19.98449, 19.98445, 19.98445, 19.98443, 19.98452, 19.98446, 19.98456, 
    19.98453, 19.98475, 19.98483, 19.98487, 19.9849, 19.98497, 19.98492, 
    19.98494, 19.98489, 19.98486, 19.98488, 19.98478, 19.98482, 19.98463, 
    19.98471, 19.9845, 19.98455, 19.98448, 19.98452, 19.98446, 19.98451, 
    19.98442, 19.98441, 19.98442, 19.98437, 19.98451, 19.98446, 19.98488, 
    19.98487, 19.98486, 19.98491, 19.98492, 19.98496, 19.98492, 19.9849, 
    19.98486, 19.98483, 19.98481, 19.98475, 19.98469, 19.98461, 19.98454, 
    19.9845, 19.98453, 19.98451, 19.98453, 19.98454, 19.98441, 19.98449, 
    19.98438, 19.98438, 19.98443, 19.98438, 19.98487, 19.98489, 19.98494, 
    19.9849, 19.98497, 19.98493, 19.98491, 19.98482, 19.9848, 19.98478, 
    19.98475, 19.9847, 19.98462, 19.98455, 19.98449, 19.9845, 19.98449, 
    19.98448, 19.98451, 19.98447, 19.98447, 19.98449, 19.98438, 19.98441, 
    19.98438, 19.9844, 19.98488, 19.98486, 19.98487, 19.98485, 19.98486, 
    19.98479, 19.98477, 19.98466, 19.9847, 19.98463, 19.9847, 19.98468, 
    19.98463, 19.98469, 19.98456, 19.98465, 19.98448, 19.98457, 19.98447, 
    19.98449, 19.98446, 19.98444, 19.9844, 19.98434, 19.98436, 19.98431, 
    19.98482, 19.98479, 19.98479, 19.98476, 19.98474, 19.98469, 19.9846, 
    19.98463, 19.98458, 19.98457, 19.98465, 19.9846, 19.98477, 19.98474, 
    19.98476, 19.98482, 19.98463, 19.98473, 19.98454, 19.9846, 19.98444, 
    19.98452, 19.98437, 19.9843, 19.98424, 19.98417, 19.98478, 19.9848, 
    19.98476, 19.98471, 19.98466, 19.98459, 19.98459, 19.98458, 19.98454, 
    19.98452, 19.98457, 19.98451, 19.98474, 19.98462, 19.9848, 19.98475, 
    19.98471, 19.98473, 19.98464, 19.98462, 19.98453, 19.98458, 19.98432, 
    19.98443, 19.98411, 19.9842, 19.9848, 19.98478, 19.98468, 19.98472, 
    19.98459, 19.98456, 19.98453, 19.9845, 19.98449, 19.98447, 19.9845, 
    19.98447, 19.98459, 19.98454, 19.98469, 19.98465, 19.98467, 19.98469, 
    19.98463, 19.98457, 19.98457, 19.98455, 19.9845, 19.98459, 19.9843, 
    19.98448, 19.98474, 19.98469, 19.98468, 19.9847, 19.98456, 19.98461, 
    19.98447, 19.98451, 19.98445, 19.98448, 19.98448, 19.98452, 19.98455, 
    19.98461, 19.98466, 19.9847, 19.98469, 19.98465, 19.98457, 19.98449, 
    19.98451, 19.98445, 19.9846, 19.98454, 19.98456, 19.9845, 19.98463, 
    19.98452, 19.98466, 19.98465, 19.98461, 19.98453, 19.98452, 19.9845, 
    19.98451, 19.98456, 19.98457, 19.98461, 19.98462, 19.98466, 19.98468, 
    19.98466, 19.98463, 19.98456, 19.9845, 19.98444, 19.98442, 19.98434, 
    19.98441, 19.9843, 19.98439, 19.98423, 19.98451, 19.98439, 19.98461, 
    19.98459, 19.98454, 19.98445, 19.9845, 19.98444, 19.98457, 19.98464, 
    19.98466, 19.9847, 19.98466, 19.98466, 19.98463, 19.98464, 19.98456, 
    19.98461, 19.98448, 19.98444, 19.98431, 19.98424, 19.98416, 19.98412, 
    19.98411, 19.98411,
  19.98606, 19.986, 19.98601, 19.98596, 19.98599, 19.98595, 19.98605, 19.986, 
    19.98603, 19.98606, 19.98586, 19.98596, 19.98576, 19.98582, 19.98566, 
    19.98577, 19.98564, 19.98566, 19.98559, 19.98561, 19.98552, 19.98558, 
    19.98547, 19.98553, 19.98552, 19.98558, 19.98594, 19.98587, 19.98594, 
    19.98593, 19.98594, 19.98599, 19.98602, 19.98607, 19.98606, 19.98602, 
    19.98593, 19.98596, 19.98588, 19.98588, 19.9858, 19.98583, 19.98569, 
    19.98573, 19.98561, 19.98564, 19.98561, 19.98562, 19.98561, 19.98565, 
    19.98564, 19.98568, 19.98583, 19.98578, 19.98592, 19.986, 19.98605, 
    19.98609, 19.98608, 19.98607, 19.98602, 19.98597, 19.98593, 19.98591, 
    19.98588, 19.98581, 19.98577, 19.98568, 19.98569, 19.98567, 19.98564, 
    19.9856, 19.98561, 19.98559, 19.98567, 19.98561, 19.9857, 19.98568, 
    19.98588, 19.98595, 19.98598, 19.98601, 19.98608, 19.98603, 19.98605, 
    19.98601, 19.98598, 19.98599, 19.98591, 19.98594, 19.98577, 19.98584, 
    19.98565, 19.98569, 19.98563, 19.98566, 19.98561, 19.98566, 19.98558, 
    19.98556, 19.98557, 19.98553, 19.98566, 19.98561, 19.98599, 19.98599, 
    19.98598, 19.98602, 19.98603, 19.98607, 19.98603, 19.98602, 19.98598, 
    19.98595, 19.98593, 19.98588, 19.98582, 19.98575, 19.98569, 19.98565, 
    19.98567, 19.98565, 19.98568, 19.98569, 19.98557, 19.98564, 19.98553, 
    19.98554, 19.98559, 19.98554, 19.98599, 19.986, 19.98605, 19.98601, 
    19.98607, 19.98604, 19.98602, 19.98594, 19.98592, 19.98591, 19.98587, 
    19.98583, 19.98576, 19.9857, 19.98564, 19.98565, 19.98564, 19.98563, 
    19.98566, 19.98563, 19.98562, 19.98564, 19.98554, 19.98557, 19.98554, 
    19.98556, 19.986, 19.98598, 19.98599, 19.98597, 19.98598, 19.98591, 
    19.98589, 19.98579, 19.98583, 19.98577, 19.98583, 19.98582, 19.98577, 
    19.98582, 19.9857, 19.98578, 19.98563, 19.98571, 19.98562, 19.98564, 
    19.98561, 19.98559, 19.98556, 19.98551, 19.98552, 19.98547, 19.98594, 
    19.98591, 19.98592, 19.98589, 19.98587, 19.98582, 19.98574, 19.98577, 
    19.98572, 19.98571, 19.98579, 19.98574, 19.9859, 19.98587, 19.98589, 
    19.98594, 19.98577, 19.98586, 19.98569, 19.98574, 19.98559, 19.98567, 
    19.98553, 19.98547, 19.98541, 19.98534, 19.9859, 19.98592, 19.98588, 
    19.98584, 19.98579, 19.98573, 19.98573, 19.98572, 19.98569, 19.98566, 
    19.98571, 19.98566, 19.98586, 19.98576, 19.98593, 19.98587, 19.98584, 
    19.98586, 19.98577, 19.98576, 19.98568, 19.98572, 19.98548, 19.98559, 
    19.98529, 19.98537, 19.98593, 19.9859, 19.98581, 19.98585, 19.98573, 
    19.9857, 19.98568, 19.98565, 19.98564, 19.98562, 19.98565, 19.98562, 
    19.98573, 19.98569, 19.98582, 19.98579, 19.9858, 19.98582, 19.98577, 
    19.98571, 19.98571, 19.98569, 19.98565, 19.98573, 19.98547, 19.98563, 
    19.98587, 19.98582, 19.98582, 19.98583, 19.9857, 19.98575, 19.98562, 
    19.98566, 19.9856, 19.98563, 19.98563, 19.98567, 19.98569, 19.98575, 
    19.98579, 19.98583, 19.98582, 19.98578, 19.98571, 19.98564, 19.98566, 
    19.98561, 19.98574, 19.98568, 19.9857, 19.98565, 19.98577, 19.98567, 
    19.9858, 19.98579, 19.98575, 19.98568, 19.98566, 19.98565, 19.98566, 
    19.98571, 19.98572, 19.98575, 19.98576, 19.98579, 19.98581, 19.98579, 
    19.98577, 19.98571, 19.98565, 19.98559, 19.98557, 19.9855, 19.98556, 
    19.98547, 19.98555, 19.9854, 19.98566, 19.98555, 19.98575, 19.98573, 
    19.98569, 19.9856, 19.98565, 19.98559, 19.98572, 19.98578, 19.9858, 
    19.98583, 19.9858, 19.9858, 19.98577, 19.98578, 19.98571, 19.98574, 
    19.98563, 19.98559, 19.98548, 19.98541, 19.98533, 19.9853, 19.98529, 
    19.98529,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222779, 0.7222756, 0.722276, 0.7222741, 0.7222751, 0.7222739, 0.7222775, 
    0.7222754, 0.7222767, 0.7222778, 0.7222703, 0.722274, 0.7222665, 
    0.7222688, 0.7222629, 0.7222669, 0.7222621, 0.722263, 0.7222604, 
    0.7222611, 0.7222576, 0.72226, 0.7222558, 0.7222582, 0.7222579, 
    0.7222601, 0.7222732, 0.7222708, 0.7222734, 0.7222731, 0.7222732, 
    0.7222751, 0.7222761, 0.7222781, 0.7222778, 0.7222763, 0.7222729, 
    0.722274, 0.7222711, 0.7222712, 0.722268, 0.7222694, 0.722264, 0.7222655, 
    0.7222611, 0.7222622, 0.7222611, 0.7222614, 0.7222611, 0.7222628, 
    0.7222621, 0.7222635, 0.7222692, 0.7222675, 0.7222725, 0.7222754, 
    0.7222774, 0.7222788, 0.7222786, 0.7222782, 0.7222763, 0.7222744, 
    0.7222731, 0.7222721, 0.7222712, 0.7222685, 0.722267, 0.7222637, 
    0.7222643, 0.7222633, 0.7222623, 0.7222607, 0.722261, 0.7222602, 
    0.7222633, 0.7222613, 0.7222646, 0.7222637, 0.722271, 0.7222737, 
    0.7222749, 0.7222759, 0.7222784, 0.7222767, 0.7222774, 0.7222757, 
    0.7222747, 0.7222753, 0.7222721, 0.7222733, 0.7222669, 0.7222697, 
    0.7222624, 0.7222642, 0.722262, 0.7222631, 0.7222613, 0.7222629, 0.72226, 
    0.7222593, 0.7222598, 0.7222581, 0.722263, 0.7222611, 0.7222753, 
    0.7222752, 0.7222748, 0.7222765, 0.7222766, 0.7222782, 0.7222767, 
    0.7222762, 0.7222747, 0.7222738, 0.7222729, 0.7222711, 0.722269, 
    0.7222661, 0.7222641, 0.7222626, 0.7222635, 0.7222627, 0.7222636, 
    0.722264, 0.7222596, 0.7222621, 0.7222583, 0.7222586, 0.7222602, 
    0.7222586, 0.7222751, 0.7222756, 0.7222772, 0.722276, 0.7222783, 
    0.722277, 0.7222762, 0.7222733, 0.7222726, 0.722272, 0.7222708, 
    0.7222694, 0.7222667, 0.7222643, 0.7222623, 0.7222624, 0.7222624, 
    0.7222619, 0.722263, 0.7222617, 0.7222615, 0.7222621, 0.7222586, 
    0.7222596, 0.7222586, 0.7222592, 0.7222754, 0.7222747, 0.7222751, 
    0.7222742, 0.7222748, 0.7222723, 0.7222715, 0.7222679, 0.7222694, 
    0.722267, 0.7222691, 0.7222688, 0.722267, 0.722269, 0.7222645, 0.7222676, 
    0.7222618, 0.7222649, 0.7222617, 0.7222623, 0.7222613, 0.7222604, 
    0.7222593, 0.7222573, 0.7222577, 0.7222561, 0.7222734, 0.7222724, 
    0.7222725, 0.7222714, 0.7222706, 0.7222688, 0.722266, 0.7222671, 
    0.7222651, 0.7222648, 0.7222677, 0.7222659, 0.7222717, 0.7222707, 
    0.7222713, 0.7222733, 0.7222669, 0.7222702, 0.722264, 0.7222658, 
    0.7222605, 0.7222632, 0.722258, 0.7222558, 0.7222537, 0.7222513, 
    0.7222718, 0.7222725, 0.7222713, 0.7222695, 0.7222679, 0.7222657, 
    0.7222655, 0.7222651, 0.7222641, 0.7222632, 0.7222649, 0.7222629, 
    0.7222705, 0.7222666, 0.7222728, 0.7222709, 0.7222696, 0.7222702, 
    0.7222672, 0.7222665, 0.7222636, 0.7222651, 0.7222564, 0.7222602, 
    0.7222494, 0.7222524, 0.7222728, 0.7222718, 0.7222685, 0.7222701, 
    0.7222655, 0.7222645, 0.7222636, 0.7222624, 0.7222623, 0.7222616, 
    0.7222627, 0.7222616, 0.7222657, 0.7222639, 0.7222689, 0.7222677, 
    0.7222682, 0.7222688, 0.722267, 0.7222649, 0.7222649, 0.7222642, 
    0.7222624, 0.7222655, 0.7222558, 0.7222618, 0.7222708, 0.7222689, 
    0.7222687, 0.7222694, 0.7222646, 0.7222663, 0.7222616, 0.7222629, 
    0.7222608, 0.7222618, 0.722262, 0.7222633, 0.7222641, 0.7222663, 
    0.7222679, 0.7222693, 0.722269, 0.7222675, 0.7222648, 0.7222623, 
    0.7222628, 0.722261, 0.7222659, 0.7222638, 0.7222646, 0.7222625, 
    0.7222671, 0.7222632, 0.7222681, 0.7222677, 0.7222664, 0.7222637, 
    0.7222631, 0.7222624, 0.7222629, 0.7222647, 0.7222651, 0.7222664, 
    0.7222667, 0.7222677, 0.7222686, 0.7222679, 0.722267, 0.7222647, 
    0.7222627, 0.7222604, 0.7222598, 0.7222572, 0.7222593, 0.7222558, 
    0.7222588, 0.7222536, 0.722263, 0.7222589, 0.7222663, 0.7222655, 
    0.7222641, 0.7222608, 0.7222626, 0.7222605, 0.7222651, 0.7222674, 
    0.722268, 0.7222692, 0.722268, 0.7222681, 0.722267, 0.7222674, 0.7222646, 
    0.7222661, 0.722262, 0.7222605, 0.7222562, 0.7222536, 0.7222509, 
    0.7222497, 0.7222494, 0.7222493 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  -1.027984e-20, 2.055969e-20, 2.006177e-36, -1.541976e-20, 0, 3.083953e-20, 
    0, 0, -5.139921e-21, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, 0, -3.083953e-20, 
    2.055969e-20, 6.167906e-20, 2.055969e-20, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, -4.111937e-20, -5.139921e-21, 
    -2.055969e-20, 2.569961e-20, 1.541976e-20, -5.139921e-21, 2.055969e-20, 
    -2.055969e-20, -2.055969e-20, 1.541976e-20, 0, 3.083953e-20, 
    -3.083953e-20, -1.027984e-20, 1.027984e-20, -1.027984e-20, 1.027984e-20, 
    -3.083953e-20, -1.027984e-20, 5.139921e-21, -5.139921e-21, -2.006177e-36, 
    1.027984e-20, 1.027984e-20, 2.055969e-20, -5.139921e-21, -2.569961e-20, 
    5.139921e-21, 2.055969e-20, -3.083953e-20, -1.027984e-20, 2.055969e-20, 
    -2.569961e-20, -4.111937e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -4.625929e-20, -1.541976e-20, -2.006177e-36, 
    1.027984e-20, -2.055969e-20, 1.027984e-20, 0, -2.569961e-20, 
    -1.027984e-20, 1.541976e-20, -2.569961e-20, 5.139921e-21, -5.139921e-21, 
    2.569961e-20, 1.541976e-20, -2.569961e-20, 5.139921e-21, -5.139921e-21, 
    -3.083953e-20, 2.055969e-20, -1.541976e-20, -1.027984e-20, -1.541976e-20, 
    5.653913e-20, -1.027984e-20, 1.027984e-20, -3.083953e-20, 0, 
    -2.055969e-20, 0, 1.027984e-20, -1.027984e-20, -1.541976e-20, 
    1.541976e-20, 1.541976e-20, -2.006177e-36, 2.055969e-20, 2.055969e-20, 
    5.139921e-21, 0, 2.055969e-20, -3.083953e-20, -2.569961e-20, 
    -2.006177e-36, 1.541976e-20, 2.569961e-20, -2.055969e-20, 3.083953e-20, 
    1.027984e-20, -5.139921e-21, -2.055969e-20, 5.139921e-21, -5.139921e-21, 
    -4.625929e-20, 1.027984e-20, 1.541976e-20, -2.006177e-36, -2.006177e-36, 
    -1.541976e-20, -3.597945e-20, 0, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, 2.569961e-20, -2.569961e-20, -1.541976e-20, -1.541976e-20, 
    0, -1.027984e-20, -1.027984e-20, -3.597945e-20, 1.541976e-20, 
    1.027984e-20, 0, -1.541976e-20, 0, 2.569961e-20, -1.541976e-20, 
    3.597945e-20, 1.027984e-20, 1.541976e-20, 2.569961e-20, -5.139921e-21, 
    3.597945e-20, 3.597945e-20, -1.541976e-20, 5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 4.111937e-20, -1.541976e-20, 5.139921e-21, -1.541976e-20, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, -2.055969e-20, -1.027984e-20, 
    1.541976e-20, 6.167906e-20, -1.027984e-20, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 0, -1.541976e-20, 3.083953e-20, -5.139921e-21, 
    -3.083953e-20, 5.139921e-21, -3.083953e-20, -2.569961e-20, -1.541976e-20, 
    -1.541976e-20, -1.027984e-20, 1.027984e-20, -4.111937e-20, 1.541976e-20, 
    -1.027984e-20, 2.569961e-20, 3.597945e-20, 2.569961e-20, 2.006177e-36, 
    -2.055969e-20, -5.139921e-21, 0, -5.139921e-21, -2.055969e-20, 
    1.027984e-20, -3.083953e-20, -1.541976e-20, 2.569961e-20, 0, 
    2.569961e-20, 5.139921e-21, 2.006177e-36, -2.569961e-20, 5.139921e-21, 
    -1.027984e-20, 3.597945e-20, -1.027984e-20, -1.541976e-20, -1.027984e-20, 
    2.055969e-20, 5.139921e-21, 1.541976e-20, 2.569961e-20, -5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 1.027984e-20, 2.569961e-20, 0, 0, 
    3.083953e-20, 2.055969e-20, 5.139921e-21, -3.597945e-20, 1.027984e-20, 
    5.139921e-21, 5.139921e-21, -3.597945e-20, 1.541976e-20, -2.055969e-20, 
    -5.139921e-21, 3.597945e-20, 0, 5.139921e-21, 3.597945e-20, 
    -5.139921e-21, 2.569961e-20, 2.569961e-20, 5.139921e-21, 0, 
    -3.083953e-20, -2.569961e-20, -2.055969e-20, -1.541976e-20, 
    -3.597945e-20, -2.006177e-36, 0, 5.139921e-21, -1.027984e-20, 
    1.027984e-20, -3.083953e-20, -3.597945e-20, -5.139921e-21, -2.055969e-20, 
    5.139921e-21, -1.027984e-20, -1.541976e-20, -5.139921e-21, 3.597945e-20, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 0, -2.569961e-20, -5.139921e-21, 
    2.055969e-20, 1.541976e-20, 0, -1.541976e-20, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    0, -2.569961e-20, 1.027984e-20, 1.541976e-20, 1.541976e-20, 
    -3.597945e-20, -1.027984e-20, -1.027984e-20, -2.055969e-20, 2.569961e-20, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, -2.055969e-20, 3.597945e-20, 
    -2.055969e-20, -1.027984e-20, 1.027984e-20, 2.055969e-20, 5.653913e-20, 
    1.541976e-20, -2.055969e-20, 3.083953e-20, 1.541976e-20, 5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, -2.055969e-20, 
    1.027984e-20, 1.541976e-20, -2.055969e-20, 0, -5.139921e-21, 
    5.139921e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 2.569961e-20, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, -1.027984e-20, 0, 
    3.083953e-20, 1.027984e-20, -5.139921e-21, 1.541976e-20, 2.569961e-20, 0, 
    2.569961e-20, 5.139921e-21, 2.569961e-20, 1.541976e-20, -3.083953e-20, 
    5.139921e-21, 1.541976e-20, -2.006177e-36, -5.139921e-21, 1.541976e-20,
  0, 3.597945e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, 0, 
    -2.006177e-36, -1.541976e-20, 5.139921e-21, -5.139921e-21, 2.569961e-20, 
    0, 1.027984e-20, 1.027984e-20, 5.139921e-21, 0, -5.139921e-21, 
    1.027984e-20, 2.569961e-20, 5.139921e-21, -1.027984e-20, -4.111937e-20, 
    1.027984e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, -1.027984e-20, 
    1.027984e-20, 2.055969e-20, 5.139921e-21, 0, 1.541976e-20, -5.139921e-21, 
    0, -5.139921e-21, 1.027984e-20, 0, -2.055969e-20, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 1.541976e-20, 1.541976e-20, -3.083953e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -2.055969e-20, -5.139921e-21, 
    -1.541976e-20, 2.569961e-20, -5.139921e-21, 0, 1.541976e-20, 
    -5.139921e-21, 1.027984e-20, -1.541976e-20, -3.083953e-20, -3.083953e-20, 
    -2.569961e-20, -2.569961e-20, 2.055969e-20, 1.027984e-20, -2.569961e-20, 
    2.006177e-36, -1.541976e-20, 0, 1.027984e-20, 5.139921e-21, 1.541976e-20, 
    3.083953e-20, -2.569961e-20, 5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, -1.027984e-20, 1.027984e-20, 0, 1.541976e-20, 
    -1.027984e-20, 2.569961e-20, -5.139921e-21, -1.541976e-20, 5.139921e-21, 
    2.569961e-20, 5.139921e-21, 2.569961e-20, -2.055969e-20, -5.139921e-21, 
    2.055969e-20, 1.027984e-20, 1.541976e-20, 1.541976e-20, 2.569961e-20, 
    2.055969e-20, 1.027984e-20, 1.027984e-20, 1.027984e-20, -2.569961e-20, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, 1.027984e-20, 5.139921e-21, 0, 
    0, -3.083953e-20, -5.139921e-21, 3.083953e-20, -1.541976e-20, 
    5.139921e-21, 2.055969e-20, 1.027984e-20, 2.055969e-20, 1.541976e-20, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, 2.055969e-20, 
    5.139921e-21, -1.541976e-20, 0, 2.569961e-20, -1.027984e-20, 
    -1.541976e-20, 5.139921e-21, -2.055969e-20, -1.541976e-20, -1.541976e-20, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, 1.027984e-20, 1.541976e-20, 3.083953e-20, 1.541976e-20, 
    3.083953e-20, -5.139921e-21, 5.139921e-21, -2.055969e-20, -4.625929e-20, 
    -1.027984e-20, -5.139921e-21, 1.027984e-20, 2.055969e-20, 1.027984e-20, 
    0, -5.139921e-21, -2.055969e-20, 1.541976e-20, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, 0, -5.139921e-21, 3.083953e-20, 
    -1.027984e-20, 1.541976e-20, 5.139921e-21, 0, -1.027984e-20, 
    -2.055969e-20, 1.027984e-20, 1.541976e-20, -3.083953e-20, 2.055969e-20, 
    1.541976e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    4.111937e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, 2.006177e-36, -3.597945e-20, -2.006177e-36, 
    -2.055969e-20, -2.006177e-36, 2.006177e-36, -1.541976e-20, 5.139921e-21, 
    5.139921e-21, -1.541976e-20, 0, 0, 2.055969e-20, 3.083953e-20, 
    5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    0, -2.569961e-20, 2.055969e-20, -2.006177e-36, 1.027984e-20, 
    1.027984e-20, -1.541976e-20, 5.139921e-21, 0, 1.541976e-20, 
    -2.055969e-20, 0, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    1.027984e-20, 1.027984e-20, -1.027984e-20, 1.027984e-20, 0, 0, 
    5.139921e-21, -1.027984e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    1.541976e-20, -1.541976e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, 0, 
    -1.541976e-20, -3.597945e-20, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 3.083953e-20, -2.055969e-20, -1.541976e-20, 1.027984e-20, 
    2.006177e-36, 5.139921e-21, 2.569961e-20, -5.139921e-21, -1.027984e-20, 
    -1.541976e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, -2.055969e-20, -2.006177e-36, -1.541976e-20, 
    2.055969e-20, 0, -2.055969e-20, 1.027984e-20, -1.027984e-20, 0, 
    2.569961e-20, -2.055969e-20, 0, -2.006177e-36, 1.541976e-20, 
    5.139921e-21, 0, -2.569961e-20, -1.027984e-20, 2.055969e-20, 
    5.139921e-21, 0, -1.541976e-20, 0, -1.027984e-20, 2.569961e-20, 
    -1.541976e-20, -2.055969e-20, -1.541976e-20, -2.055969e-20, 0, 
    1.541976e-20, 2.569961e-20, -4.111937e-20, -2.569961e-20, -1.541976e-20, 
    1.541976e-20, -1.541976e-20, 5.139921e-21, 0, -1.541976e-20, 
    2.055969e-20, 0, -1.027984e-20, 0, 5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 1.027984e-20, 0, 1.541976e-20, 2.006177e-36, 
    -1.541976e-20, 0, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    2.055969e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, 0, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, 0, -2.055969e-20, 
    -2.055969e-20, 1.027984e-20, -1.027984e-20, -2.055969e-20, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    0, -5.139921e-21, 5.139921e-21, 3.083953e-20,
  3.083953e-20, -5.139921e-21, -5.139921e-21, 1.541976e-20, 1.541976e-20, 
    2.055969e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 2.055969e-20, -1.541976e-20, -1.027984e-20, 0, 
    2.569961e-20, 1.541976e-20, -1.027984e-20, -1.541976e-20, 2.055969e-20, 
    -2.569961e-20, -2.055969e-20, -2.569961e-20, -1.541976e-20, 5.139921e-21, 
    0, -1.027984e-20, -5.139921e-21, -2.055969e-20, -1.541976e-20, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    2.006177e-36, -2.055969e-20, 1.027984e-20, -1.027984e-20, -1.027984e-20, 
    5.139921e-21, -2.569961e-20, 5.139921e-21, 3.597945e-20, 2.055969e-20, 
    1.027984e-20, -1.027984e-20, 0, -1.027984e-20, -2.006177e-36, 
    2.006177e-36, 3.083953e-20, 2.569961e-20, 1.541976e-20, 0, 2.055969e-20, 
    -5.139921e-21, -2.055969e-20, 0, -3.597945e-20, -1.027984e-20, 
    2.055969e-20, 1.541976e-20, -3.597945e-20, 0, 2.055969e-20, 5.139921e-21, 
    -1.541976e-20, 1.027984e-20, 0, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, -2.055969e-20, 0, 2.569961e-20, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -2.569961e-20, -3.083953e-20, -2.569961e-20, 
    -2.006177e-36, -1.027984e-20, 5.139921e-21, -2.006177e-36, 5.139921e-21, 
    -2.055969e-20, 0, 5.139921e-21, -2.569961e-20, 1.027984e-20, 
    1.541976e-20, -3.597945e-20, -5.139921e-21, 3.083953e-20, -5.139921e-21, 
    1.541976e-20, 1.541976e-20, 0, -2.055969e-20, 1.541976e-20, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 2.569961e-20, 3.083953e-20, 2.569961e-20, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, -1.027984e-20, -2.055969e-20, 
    0, -5.139921e-21, 1.027984e-20, -1.027984e-20, 2.006177e-36, 
    -1.541976e-20, -1.541976e-20, -2.055969e-20, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, 0, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, -2.569961e-20, 1.027984e-20, -5.139921e-21, -2.006177e-36, 
    5.139921e-21, 2.006177e-36, -5.139921e-21, -2.006177e-36, 0, 
    -5.139921e-21, -2.006177e-36, -1.027984e-20, -1.027984e-20, 1.541976e-20, 
    -1.541976e-20, -5.139921e-21, 0, 0, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, 2.055969e-20, -5.139921e-21, 2.006177e-36, 
    3.597945e-20, 0, 5.139921e-21, 5.139921e-21, 3.083953e-20, -1.541976e-20, 
    1.027984e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, 
    1.541976e-20, -3.083953e-20, 1.541976e-20, 2.055969e-20, 2.055969e-20, 
    2.055969e-20, -3.597945e-20, -1.541976e-20, 5.139921e-21, 5.139921e-21, 
    3.597945e-20, -1.027984e-20, 1.541976e-20, -1.027984e-20, -2.006177e-36, 
    -1.027984e-20, 0, 3.083953e-20, -5.139921e-21, 2.569961e-20, 
    -1.027984e-20, 5.139921e-21, -1.541976e-20, 1.541976e-20, 1.027984e-20, 
    0, -1.541976e-20, 5.139921e-21, -5.139921e-21, 0, -5.139921e-21, 
    -2.055969e-20, 0, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    1.541976e-20, -2.006177e-36, -1.541976e-20, -1.027984e-20, 2.006177e-36, 
    3.083953e-20, 3.083953e-20, -1.027984e-20, 1.541976e-20, -1.027984e-20, 
    1.027984e-20, -1.541976e-20, -5.139921e-21, 0, 0, -4.111937e-20, 
    5.139921e-21, -2.006177e-36, -1.541976e-20, 0, -5.139921e-21, 
    1.541976e-20, 3.083953e-20, 5.139921e-21, 5.139921e-21, -1.541976e-20, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 1.027984e-20, 0, -2.055969e-20, 1.027984e-20, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, 
    -2.569961e-20, -1.027984e-20, -1.027984e-20, -1.541976e-20, 2.055969e-20, 
    1.541976e-20, -5.139921e-21, 5.139921e-21, -1.541976e-20, -1.541976e-20, 
    1.541976e-20, 1.541976e-20, 5.139921e-21, 0, -1.541976e-20, 2.006177e-36, 
    -5.139921e-21, 1.541976e-20, -3.083953e-20, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, -1.541976e-20, -5.139921e-20, 4.111937e-20, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -3.083953e-20, 2.569961e-20, -2.055969e-20, 
    5.139921e-21, -2.006177e-36, -1.541976e-20, 2.055969e-20, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, -1.027984e-20, -2.006177e-36, 2.569961e-20, 
    1.027984e-20, -5.139921e-21, -2.055969e-20, -2.055969e-20, -2.055969e-20, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, 1.027984e-20, 1.027984e-20, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, -2.569961e-20, 3.597945e-20, 
    0, 0, 2.006177e-36, 5.139921e-21, -1.541976e-20, -1.541976e-20, 
    -3.597945e-20, -2.006177e-36, 2.055969e-20, 5.139921e-21, -1.027984e-20, 
    -2.055969e-20, 1.541976e-20, -5.139921e-21, 2.569961e-20, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, 3.083953e-20, -1.027984e-20, -1.541976e-20, 
    -2.055969e-20, 4.111937e-20, -2.055969e-20, -3.083953e-20, 1.027984e-20, 
    -2.055969e-20, 4.625929e-20, 2.055969e-20, -2.006177e-36, -1.027984e-20, 
    -5.139921e-21, 2.569961e-20, 2.055969e-20, 1.541976e-20, 2.569961e-20, 
    -5.139921e-21, 1.541976e-20, 2.006177e-36, 1.541976e-20,
  1.027984e-20, 3.083953e-20, 2.006177e-36, 0, 0, -1.027984e-20, 
    -2.569961e-20, -2.569961e-20, 0, 0, 1.027984e-20, 1.027984e-20, 0, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, -1.027984e-20, -1.027984e-20, 
    2.055969e-20, -1.027984e-20, 1.027984e-20, -3.597945e-20, -1.027984e-20, 
    1.541976e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, 2.055969e-20, 
    2.569961e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 2.569961e-20, 
    2.569961e-20, -5.139921e-21, 5.139921e-21, -4.625929e-20, 3.597945e-20, 
    5.139921e-21, 0, 1.541976e-20, 1.027984e-20, -1.541976e-20, 
    -1.541976e-20, 0, 2.006177e-36, -3.083953e-20, 5.139921e-21, 
    -2.569961e-20, -5.139921e-21, -1.541976e-20, 1.027984e-20, 5.139921e-21, 
    1.027984e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, 3.597945e-20, 
    1.541976e-20, -2.055969e-20, 0, 5.139921e-21, 0, -5.139921e-21, 
    -2.055969e-20, -3.597945e-20, -5.139921e-21, -2.006177e-36, 1.541976e-20, 
    1.027984e-20, -1.027984e-20, -2.006177e-36, 1.541976e-20, -1.027984e-20, 
    -5.139921e-21, -2.569961e-20, 1.027984e-20, 3.597945e-20, -1.541976e-20, 
    2.055969e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 0, 
    -3.597945e-20, 2.055969e-20, -2.569961e-20, -1.541976e-20, -2.055969e-20, 
    1.027984e-20, -1.541976e-20, -1.027984e-20, 5.139921e-21, 0, 
    2.569961e-20, 1.541976e-20, 3.597945e-20, 1.027984e-20, 1.027984e-20, 
    -1.541976e-20, 2.006177e-36, 2.569961e-20, 3.597945e-20, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, -5.139921e-21, 1.541976e-20, -1.541976e-20, 
    -5.139921e-21, -2.569961e-20, 5.139921e-21, -2.055969e-20, -1.027984e-20, 
    -2.055969e-20, 4.111937e-20, -2.569961e-20, 2.569961e-20, -2.006177e-36, 
    0, 2.569961e-20, -1.027984e-20, -2.569961e-20, 5.139921e-21, 
    1.541976e-20, 5.139921e-21, -2.569961e-20, 2.055969e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 2.055969e-20, 2.569961e-20, -2.006177e-36, 
    -5.139921e-21, 2.055969e-20, -2.055969e-20, -2.569961e-20, 1.541976e-20, 
    -5.139921e-21, 2.055969e-20, -1.027984e-20, 1.027984e-20, -3.083953e-20, 
    5.139921e-21, 3.083953e-20, -5.139921e-21, -2.569961e-20, 3.083953e-20, 
    0, -1.027984e-20, -2.006177e-36, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, -2.055969e-20, -5.139921e-21, 2.569961e-20, 0, 
    -2.569961e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -1.541976e-20, -1.027984e-20, 5.139921e-21, -3.597945e-20, -1.027984e-20, 
    2.006177e-36, -1.027984e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 1.541976e-20, -1.541976e-20, 5.139921e-21, 2.055969e-20, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 2.006177e-36, 
    1.027984e-20, -3.083953e-20, -1.027984e-20, -1.541976e-20, 1.541976e-20, 
    -2.055969e-20, 2.006177e-36, -1.541976e-20, 1.541976e-20, -1.027984e-20, 
    0, 5.139921e-21, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    -5.653913e-20, 1.027984e-20, -2.569961e-20, -5.139921e-21, -5.139921e-21, 
    4.111937e-20, -1.027984e-20, -1.027984e-20, -1.027984e-20, 2.006177e-36, 
    -1.027984e-20, -2.055969e-20, -1.541976e-20, 0, -5.139921e-21, 
    1.027984e-20, 2.055969e-20, -1.541976e-20, -2.006177e-36, 1.027984e-20, 
    1.541976e-20, 1.541976e-20, 3.597945e-20, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, 2.055969e-20, -5.139921e-21, 2.569961e-20, 3.597945e-20, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, 0, 1.027984e-20, 0, 
    1.541976e-20, -5.139921e-21, -2.006177e-36, 1.027984e-20, -1.027984e-20, 
    -2.006177e-36, 5.139921e-21, 1.027984e-20, 5.139921e-21, 2.006177e-36, 
    -2.006177e-36, 0, -5.139921e-21, 2.006177e-36, 2.055969e-20, 0, 
    -1.541976e-20, -2.055969e-20, 1.027984e-20, -2.055969e-20, 2.055969e-20, 
    -1.541976e-20, -5.653913e-20, 2.006177e-36, -2.055969e-20, -3.597945e-20, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, -3.597945e-20, -2.569961e-20, -1.027984e-20, -3.597945e-20, 
    -5.139921e-21, 3.597945e-20, 5.139921e-21, 0, 5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 5.139921e-21, -1.027984e-20, -1.541976e-20, -5.139921e-21, 
    5.139921e-21, 3.083953e-20, -5.139921e-21, -2.569961e-20, 0, 
    2.006177e-36, 0, 1.027984e-20, 3.083953e-20, 2.569961e-20, 5.139921e-21, 
    0, 5.139921e-21, 2.006177e-36, -5.139921e-21, 3.597945e-20, 1.027984e-20, 
    -2.569961e-20, 2.569961e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    1.541976e-20, -2.569961e-20, 2.006177e-36, -5.653913e-20, 0, 
    1.027984e-20, 3.083953e-20, -4.111937e-20, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 2.569961e-20, 0, -1.541976e-20, -2.055969e-20, 
    4.625929e-20, -5.139921e-21, 2.055969e-20, 0, -2.569961e-20, 
    -1.541976e-20, 2.569961e-20, -2.006177e-36, -2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 1.541976e-20, 1.541976e-20, 4.111937e-20, -4.111937e-20, 
    2.569961e-20, 2.055969e-20, 5.139921e-21, -1.027984e-20,
  2.569961e-20, -1.027984e-20, 2.055969e-20, 4.111937e-20, -5.139921e-21, 
    -1.541976e-20, -2.055969e-20, 2.006177e-36, 1.027984e-20, -5.139921e-21, 
    1.541976e-20, 4.111937e-20, 5.139921e-21, -3.597945e-20, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -2.569961e-20, 0, -1.027984e-20, 
    -2.006177e-36, 1.027984e-20, 2.055969e-20, -2.055969e-20, 5.139921e-21, 
    1.541976e-20, 3.083953e-20, -1.541976e-20, -2.055969e-20, -1.027984e-20, 
    -1.027984e-20, 1.541976e-20, 1.027984e-20, 2.055969e-20, 4.111937e-20, 0, 
    1.027984e-20, 1.541976e-20, -2.569961e-20, 1.541976e-20, -1.541976e-20, 
    5.139921e-21, 5.139921e-21, 0, -1.027984e-20, -3.083953e-20, 
    2.055969e-20, 0, 1.541976e-20, -5.139921e-21, 3.597945e-20, 5.139921e-21, 
    2.569961e-20, -2.569961e-20, -1.541976e-20, 5.139921e-21, -2.569961e-20, 
    -2.006177e-36, -1.027984e-20, -5.139921e-21, 1.027984e-20, 4.111937e-20, 
    1.027984e-20, -1.541976e-20, -2.055969e-20, -4.625929e-20, 1.541976e-20, 
    0, -1.027984e-20, 2.569961e-20, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, 1.027984e-20, -1.541976e-20, -2.006177e-36, 
    1.541976e-20, -2.055969e-20, -1.027984e-20, 0, 1.541976e-20, 
    5.139921e-21, 2.055969e-20, -1.541976e-20, -1.541976e-20, -2.006177e-36, 
    1.027984e-20, 0, -1.541976e-20, 2.006177e-36, -1.027984e-20, 
    5.139921e-21, -2.055969e-20, -1.027984e-20, -2.569961e-20, -1.027984e-20, 
    1.027984e-20, -2.055969e-20, 2.569961e-20, -1.541976e-20, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 5.139921e-21, 2.055969e-20, -2.569961e-20, 
    -2.006177e-36, 5.139921e-21, -3.597945e-20, -1.541976e-20, 0, 
    5.139921e-21, -5.139921e-21, -3.597945e-20, 2.006177e-36, -1.541976e-20, 
    -2.569961e-20, -5.139921e-21, 1.027984e-20, 2.055969e-20, 0, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, 3.083953e-20, -1.027984e-20, 
    -5.139921e-21, -2.055969e-20, -2.055969e-20, -2.006177e-36, 1.027984e-20, 
    -5.139921e-21, -2.055969e-20, -5.139921e-21, 2.006177e-36, 2.569961e-20, 
    2.055969e-20, -5.139921e-21, -3.597945e-20, -2.569961e-20, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, 2.055969e-20, 4.111937e-20, 
    3.083953e-20, -1.027984e-20, 5.139921e-21, 2.006177e-36, 5.139921e-21, 
    -1.027984e-20, -5.139921e-21, -1.541976e-20, 2.006177e-36, -2.055969e-20, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 1.027984e-20, 
    -1.027984e-20, 2.055969e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    -2.055969e-20, -2.569961e-20, -1.541976e-20, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 2.055969e-20, -3.083953e-20, 2.055969e-20, 5.139921e-21, 
    5.139921e-21, 0, -1.541976e-20, 1.027984e-20, -5.139921e-21, 0, 
    -1.027984e-20, -1.027984e-20, 3.083953e-20, -1.541976e-20, -5.139921e-21, 
    0, -5.139921e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    1.027984e-20, -1.541976e-20, 2.006177e-36, -5.139921e-21, -1.541976e-20, 
    2.569961e-20, -2.055969e-20, 1.027984e-20, -2.569961e-20, 1.541976e-20, 
    -1.541976e-20, -3.083953e-20, -1.541976e-20, 3.083953e-20, 3.597945e-20, 
    1.541976e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 0, -1.541976e-20, 
    0, -1.027984e-20, -1.541976e-20, 2.569961e-20, -5.139921e-21, 
    -1.541976e-20, 2.569961e-20, 1.541976e-20, -5.139921e-21, -3.597945e-20, 
    -3.597945e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, -1.027984e-20, 
    2.569961e-20, 5.139921e-21, 5.139921e-21, 3.597945e-20, -4.111937e-20, 
    -2.006177e-36, 2.569961e-20, -1.027984e-20, 3.597945e-20, -3.083953e-20, 
    -4.111937e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, -2.569961e-20, 
    3.083953e-20, -1.541976e-20, 0, 3.083953e-20, -2.055969e-20, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 0, 
    -1.027984e-20, -2.006177e-36, -1.541976e-20, 1.027984e-20, 5.139921e-21, 
    1.027984e-20, 2.569961e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, 
    2.569961e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -2.006177e-36, -5.139921e-21, 5.139921e-21, -5.139921e-21, -1.541976e-20, 
    5.139921e-21, 3.597945e-20, 5.139921e-21, -2.055969e-20, 2.055969e-20, 
    -1.541976e-20, -2.006177e-36, 2.055969e-20, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, 1.027984e-20, 0, -2.055969e-20, -5.139921e-21, 0, 
    1.027984e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, -2.006177e-36, 
    5.139921e-21, -2.569961e-20, 1.541976e-20, -5.139921e-21, -2.055969e-20, 
    -5.139921e-21, 0, 1.541976e-20, 2.569961e-20, 1.027984e-20, 0, 
    -2.569961e-20, -5.139921e-21, -2.569961e-20, 3.083953e-20, 5.139921e-21, 
    -1.027984e-20, -2.006177e-36, -1.541976e-20, 1.541976e-20, 1.541976e-20, 
    -2.055969e-20, 1.541976e-20, -4.111937e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.541976e-20, 3.083953e-20, 5.139921e-21, 
    -2.569961e-20, -1.027984e-20, 0, 1.027984e-20, 1.541976e-20, 
    -1.541976e-20, 1.541976e-20, 5.139921e-21, 2.055969e-20, -5.139921e-21, 
    1.027984e-20, -2.055969e-20,
  8.598819e-29, 8.59879e-29, 8.598796e-29, 8.598773e-29, 8.598786e-29, 
    8.598771e-29, 8.598813e-29, 8.598789e-29, 8.598804e-29, 8.598816e-29, 
    8.59873e-29, 8.598772e-29, 8.598685e-29, 8.598713e-29, 8.598643e-29, 
    8.598689e-29, 8.598634e-29, 8.598645e-29, 8.598613e-29, 8.598622e-29, 
    8.598582e-29, 8.598609e-29, 8.598561e-29, 8.598589e-29, 8.598584e-29, 
    8.59861e-29, 8.598764e-29, 8.598735e-29, 8.598766e-29, 8.598761e-29, 
    8.598763e-29, 8.598785e-29, 8.598797e-29, 8.59882e-29, 8.598816e-29, 
    8.598799e-29, 8.59876e-29, 8.598773e-29, 8.598739e-29, 8.59874e-29, 
    8.598702e-29, 8.598719e-29, 8.598656e-29, 8.598674e-29, 8.598622e-29, 
    8.598635e-29, 8.598622e-29, 8.598627e-29, 8.598622e-29, 8.598642e-29, 
    8.598634e-29, 8.598651e-29, 8.598716e-29, 8.598697e-29, 8.598754e-29, 
    8.598788e-29, 8.598812e-29, 8.598828e-29, 8.598826e-29, 8.598821e-29, 
    8.598799e-29, 8.598778e-29, 8.598761e-29, 8.598751e-29, 8.59874e-29, 
    8.598708e-29, 8.59869e-29, 8.598652e-29, 8.598659e-29, 8.598648e-29, 
    8.598636e-29, 8.598618e-29, 8.598621e-29, 8.598613e-29, 8.598648e-29, 
    8.598624e-29, 8.598663e-29, 8.598652e-29, 8.598737e-29, 8.598769e-29, 
    8.598783e-29, 8.598795e-29, 8.598824e-29, 8.598804e-29, 8.598812e-29, 
    8.598793e-29, 8.598781e-29, 8.598787e-29, 8.598751e-29, 8.598764e-29, 
    8.59869e-29, 8.598722e-29, 8.598638e-29, 8.598658e-29, 8.598633e-29, 
    8.598646e-29, 8.598624e-29, 8.598643e-29, 8.598609e-29, 8.598602e-29, 
    8.598607e-29, 8.598587e-29, 8.598645e-29, 8.598622e-29, 8.598787e-29, 
    8.598786e-29, 8.598781e-29, 8.598801e-29, 8.598802e-29, 8.59882e-29, 
    8.598805e-29, 8.598798e-29, 8.59878e-29, 8.59877e-29, 8.59876e-29, 
    8.598739e-29, 8.598714e-29, 8.598681e-29, 8.598657e-29, 8.59864e-29, 
    8.59865e-29, 8.598642e-29, 8.598651e-29, 8.598656e-29, 8.598605e-29, 
    8.598633e-29, 8.59859e-29, 8.598593e-29, 8.598612e-29, 8.598592e-29, 
    8.598785e-29, 8.598791e-29, 8.59881e-29, 8.598795e-29, 8.598823e-29, 
    8.598807e-29, 8.598798e-29, 8.598764e-29, 8.598757e-29, 8.59875e-29, 
    8.598736e-29, 8.598719e-29, 8.598687e-29, 8.59866e-29, 8.598636e-29, 
    8.598637e-29, 8.598637e-29, 8.598631e-29, 8.598645e-29, 8.598629e-29, 
    8.598627e-29, 8.598633e-29, 8.598593e-29, 8.598604e-29, 8.598593e-29, 
    8.5986e-29, 8.598789e-29, 8.59878e-29, 8.598785e-29, 8.598775e-29, 
    8.598782e-29, 8.598752e-29, 8.598743e-29, 8.598702e-29, 8.598719e-29, 
    8.598692e-29, 8.598716e-29, 8.598711e-29, 8.59869e-29, 8.598714e-29, 
    8.598662e-29, 8.598698e-29, 8.598631e-29, 8.598667e-29, 8.598629e-29, 
    8.598636e-29, 8.598624e-29, 8.598614e-29, 8.598601e-29, 8.598578e-29, 
    8.598583e-29, 8.598563e-29, 8.598766e-29, 8.598754e-29, 8.598755e-29, 
    8.598742e-29, 8.598733e-29, 8.598713e-29, 8.59868e-29, 8.598692e-29, 
    8.598669e-29, 8.598665e-29, 8.598699e-29, 8.598678e-29, 8.598746e-29, 
    8.598735e-29, 8.598741e-29, 8.598765e-29, 8.598689e-29, 8.598728e-29, 
    8.598656e-29, 8.598677e-29, 8.598616e-29, 8.598646e-29, 8.598586e-29, 
    8.59856e-29, 8.598536e-29, 8.598507e-29, 8.598747e-29, 8.598755e-29, 
    8.59874e-29, 8.59872e-29, 8.598701e-29, 8.598676e-29, 8.598674e-29, 
    8.598669e-29, 8.598657e-29, 8.598646e-29, 8.598667e-29, 8.598643e-29, 
    8.598732e-29, 8.598686e-29, 8.598758e-29, 8.598737e-29, 8.598721e-29, 
    8.598728e-29, 8.598693e-29, 8.598685e-29, 8.598652e-29, 8.598669e-29, 
    8.598567e-29, 8.598612e-29, 8.598486e-29, 8.598521e-29, 8.598758e-29, 
    8.598747e-29, 8.598708e-29, 8.598727e-29, 8.598674e-29, 8.598662e-29, 
    8.598651e-29, 8.598637e-29, 8.598636e-29, 8.598628e-29, 8.598641e-29, 
    8.598628e-29, 8.598676e-29, 8.598655e-29, 8.598713e-29, 8.598699e-29, 
    8.598705e-29, 8.598713e-29, 8.59869e-29, 8.598667e-29, 8.598666e-29, 
    8.598659e-29, 8.598637e-29, 8.598674e-29, 8.598561e-29, 8.598631e-29, 
    8.598735e-29, 8.598714e-29, 8.598711e-29, 8.598719e-29, 8.598663e-29, 
    8.598683e-29, 8.598628e-29, 8.598643e-29, 8.598619e-29, 8.598631e-29, 
    8.598633e-29, 8.598648e-29, 8.598658e-29, 8.598682e-29, 8.598702e-29, 
    8.598717e-29, 8.598714e-29, 8.598697e-29, 8.598666e-29, 8.598636e-29, 
    8.598642e-29, 8.598621e-29, 8.598678e-29, 8.598654e-29, 8.598663e-29, 
    8.598639e-29, 8.598692e-29, 8.598647e-29, 8.598704e-29, 8.598699e-29, 
    8.598683e-29, 8.598652e-29, 8.598645e-29, 8.598638e-29, 8.598643e-29, 
    8.598665e-29, 8.598668e-29, 8.598684e-29, 8.598688e-29, 8.5987e-29, 
    8.59871e-29, 8.598701e-29, 8.598692e-29, 8.598665e-29, 8.59864e-29, 
    8.598614e-29, 8.598608e-29, 8.598577e-29, 8.598602e-29, 8.59856e-29, 
    8.598596e-29, 8.598535e-29, 8.598644e-29, 8.598597e-29, 8.598683e-29, 
    8.598674e-29, 8.598657e-29, 8.598618e-29, 8.598639e-29, 8.598615e-29, 
    8.598668e-29, 8.598696e-29, 8.598704e-29, 8.598717e-29, 8.598703e-29, 
    8.598704e-29, 8.598691e-29, 8.598695e-29, 8.598664e-29, 8.598681e-29, 
    8.598633e-29, 8.598615e-29, 8.598565e-29, 8.598535e-29, 8.598504e-29, 
    8.59849e-29, 8.598486e-29, 8.598484e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.138939e-08, 1.14396e-08, 1.142984e-08, 1.147034e-08, 1.144787e-08, 
    1.147439e-08, 1.139957e-08, 1.144159e-08, 1.141477e-08, 1.139391e-08, 
    1.154893e-08, 1.147214e-08, 1.162871e-08, 1.157973e-08, 1.170277e-08, 
    1.162108e-08, 1.171924e-08, 1.170041e-08, 1.175708e-08, 1.174085e-08, 
    1.181333e-08, 1.176458e-08, 1.185091e-08, 1.180169e-08, 1.180939e-08, 
    1.176297e-08, 1.14876e-08, 1.153937e-08, 1.148453e-08, 1.149191e-08, 
    1.14886e-08, 1.144834e-08, 1.142804e-08, 1.138555e-08, 1.139327e-08, 
    1.142448e-08, 1.149523e-08, 1.147122e-08, 1.153175e-08, 1.153038e-08, 
    1.159778e-08, 1.156739e-08, 1.168068e-08, 1.164848e-08, 1.174153e-08, 
    1.171813e-08, 1.174043e-08, 1.173366e-08, 1.174052e-08, 1.170619e-08, 
    1.17209e-08, 1.16907e-08, 1.157308e-08, 1.160765e-08, 1.150456e-08, 
    1.144257e-08, 1.140141e-08, 1.13722e-08, 1.137633e-08, 1.13842e-08, 
    1.142466e-08, 1.14627e-08, 1.149169e-08, 1.151108e-08, 1.153019e-08, 
    1.158802e-08, 1.161863e-08, 1.168719e-08, 1.167482e-08, 1.169577e-08, 
    1.17158e-08, 1.174941e-08, 1.174388e-08, 1.175869e-08, 1.169522e-08, 
    1.17374e-08, 1.166777e-08, 1.168682e-08, 1.153537e-08, 1.14777e-08, 
    1.145317e-08, 1.143172e-08, 1.137951e-08, 1.141556e-08, 1.140135e-08, 
    1.143516e-08, 1.145665e-08, 1.144602e-08, 1.151161e-08, 1.148611e-08, 
    1.162045e-08, 1.156258e-08, 1.171346e-08, 1.167736e-08, 1.172212e-08, 
    1.169928e-08, 1.173841e-08, 1.170319e-08, 1.17642e-08, 1.177749e-08, 
    1.176841e-08, 1.180329e-08, 1.170124e-08, 1.174043e-08, 1.144572e-08, 
    1.144746e-08, 1.145553e-08, 1.142004e-08, 1.141787e-08, 1.138534e-08, 
    1.141428e-08, 1.142661e-08, 1.14579e-08, 1.14764e-08, 1.149399e-08, 
    1.153267e-08, 1.157588e-08, 1.163629e-08, 1.16797e-08, 1.170879e-08, 
    1.169095e-08, 1.17067e-08, 1.16891e-08, 1.168084e-08, 1.177251e-08, 
    1.172104e-08, 1.179827e-08, 1.1794e-08, 1.175904e-08, 1.179448e-08, 
    1.144867e-08, 1.14387e-08, 1.140407e-08, 1.143117e-08, 1.13818e-08, 
    1.140944e-08, 1.142532e-08, 1.148664e-08, 1.150012e-08, 1.151261e-08, 
    1.153728e-08, 1.156895e-08, 1.16245e-08, 1.167283e-08, 1.171696e-08, 
    1.171373e-08, 1.171487e-08, 1.172472e-08, 1.170031e-08, 1.172873e-08, 
    1.17335e-08, 1.172103e-08, 1.179343e-08, 1.177275e-08, 1.179391e-08, 
    1.178044e-08, 1.144194e-08, 1.145872e-08, 1.144966e-08, 1.146671e-08, 
    1.145469e-08, 1.150811e-08, 1.152413e-08, 1.159908e-08, 1.156832e-08, 
    1.161728e-08, 1.15733e-08, 1.158109e-08, 1.161887e-08, 1.157567e-08, 
    1.167017e-08, 1.16061e-08, 1.172511e-08, 1.166112e-08, 1.172912e-08, 
    1.171677e-08, 1.173721e-08, 1.175552e-08, 1.177856e-08, 1.182106e-08, 
    1.181122e-08, 1.184676e-08, 1.148374e-08, 1.150551e-08, 1.15036e-08, 
    1.152638e-08, 1.154322e-08, 1.157974e-08, 1.163831e-08, 1.161629e-08, 
    1.165673e-08, 1.166484e-08, 1.160341e-08, 1.164113e-08, 1.152008e-08, 
    1.153963e-08, 1.152799e-08, 1.148546e-08, 1.162136e-08, 1.155161e-08, 
    1.168041e-08, 1.164263e-08, 1.175291e-08, 1.169806e-08, 1.18058e-08, 
    1.185185e-08, 1.18952e-08, 1.194586e-08, 1.151739e-08, 1.15026e-08, 
    1.152909e-08, 1.156573e-08, 1.159973e-08, 1.164493e-08, 1.164956e-08, 
    1.165802e-08, 1.167996e-08, 1.169841e-08, 1.16607e-08, 1.170303e-08, 
    1.154417e-08, 1.162742e-08, 1.149701e-08, 1.153627e-08, 1.156357e-08, 
    1.15516e-08, 1.161377e-08, 1.162843e-08, 1.168798e-08, 1.165719e-08, 
    1.184048e-08, 1.175938e-08, 1.198443e-08, 1.192154e-08, 1.149743e-08, 
    1.151734e-08, 1.158663e-08, 1.155366e-08, 1.164795e-08, 1.167116e-08, 
    1.169003e-08, 1.171415e-08, 1.171675e-08, 1.173104e-08, 1.170762e-08, 
    1.173012e-08, 1.164503e-08, 1.168305e-08, 1.157871e-08, 1.160411e-08, 
    1.159242e-08, 1.157961e-08, 1.161916e-08, 1.166129e-08, 1.16622e-08, 
    1.167571e-08, 1.171377e-08, 1.164833e-08, 1.185094e-08, 1.172581e-08, 
    1.153905e-08, 1.15774e-08, 1.158288e-08, 1.156802e-08, 1.166883e-08, 
    1.16323e-08, 1.173069e-08, 1.17041e-08, 1.174767e-08, 1.172602e-08, 
    1.172284e-08, 1.169503e-08, 1.167772e-08, 1.163398e-08, 1.159839e-08, 
    1.157018e-08, 1.157674e-08, 1.160773e-08, 1.166387e-08, 1.171699e-08, 
    1.170535e-08, 1.174436e-08, 1.164111e-08, 1.16844e-08, 1.166767e-08, 
    1.17113e-08, 1.16157e-08, 1.16971e-08, 1.15949e-08, 1.160386e-08, 
    1.163158e-08, 1.168734e-08, 1.169968e-08, 1.171285e-08, 1.170472e-08, 
    1.16653e-08, 1.165884e-08, 1.163091e-08, 1.162319e-08, 1.160191e-08, 
    1.158428e-08, 1.160038e-08, 1.161729e-08, 1.166531e-08, 1.170859e-08, 
    1.175578e-08, 1.176733e-08, 1.182246e-08, 1.177758e-08, 1.185164e-08, 
    1.178867e-08, 1.189768e-08, 1.170183e-08, 1.178682e-08, 1.163284e-08, 
    1.164943e-08, 1.167943e-08, 1.174825e-08, 1.17111e-08, 1.175455e-08, 
    1.165859e-08, 1.16088e-08, 1.159592e-08, 1.157189e-08, 1.159647e-08, 
    1.159447e-08, 1.161799e-08, 1.161044e-08, 1.166691e-08, 1.163657e-08, 
    1.172276e-08, 1.17542e-08, 1.184303e-08, 1.189748e-08, 1.195292e-08, 
    1.197739e-08, 1.198484e-08, 1.198796e-08 ;

 SOIL1N_TO_SOIL3N =
  1.351374e-10, 1.357334e-10, 1.356176e-10, 1.360982e-10, 1.358316e-10, 
    1.361463e-10, 1.352583e-10, 1.35757e-10, 1.354386e-10, 1.351911e-10, 
    1.370311e-10, 1.361197e-10, 1.37978e-10, 1.373967e-10, 1.388572e-10, 
    1.378875e-10, 1.390527e-10, 1.388292e-10, 1.395019e-10, 1.393092e-10, 
    1.401696e-10, 1.395909e-10, 1.406157e-10, 1.400314e-10, 1.401228e-10, 
    1.395718e-10, 1.363031e-10, 1.369176e-10, 1.362667e-10, 1.363543e-10, 
    1.36315e-10, 1.358371e-10, 1.355962e-10, 1.350919e-10, 1.351835e-10, 
    1.355539e-10, 1.363937e-10, 1.361087e-10, 1.368272e-10, 1.36811e-10, 
    1.37611e-10, 1.372503e-10, 1.385949e-10, 1.382127e-10, 1.393172e-10, 
    1.390395e-10, 1.393042e-10, 1.392239e-10, 1.393052e-10, 1.388978e-10, 
    1.390724e-10, 1.387139e-10, 1.373178e-10, 1.377281e-10, 1.365044e-10, 
    1.357687e-10, 1.352801e-10, 1.349334e-10, 1.349825e-10, 1.350759e-10, 
    1.355561e-10, 1.360076e-10, 1.363517e-10, 1.365818e-10, 1.368086e-10, 
    1.374951e-10, 1.378585e-10, 1.386722e-10, 1.385254e-10, 1.387741e-10, 
    1.390118e-10, 1.394108e-10, 1.393452e-10, 1.39521e-10, 1.387676e-10, 
    1.392683e-10, 1.384417e-10, 1.386678e-10, 1.368702e-10, 1.361856e-10, 
    1.358945e-10, 1.356398e-10, 1.350201e-10, 1.354481e-10, 1.352794e-10, 
    1.356807e-10, 1.359358e-10, 1.358096e-10, 1.365881e-10, 1.362855e-10, 
    1.3788e-10, 1.371932e-10, 1.389841e-10, 1.385555e-10, 1.390868e-10, 
    1.388157e-10, 1.392802e-10, 1.388622e-10, 1.395864e-10, 1.397441e-10, 
    1.396363e-10, 1.400504e-10, 1.38839e-10, 1.393042e-10, 1.358061e-10, 
    1.358267e-10, 1.359225e-10, 1.355012e-10, 1.354754e-10, 1.350894e-10, 
    1.354329e-10, 1.355792e-10, 1.359506e-10, 1.361702e-10, 1.36379e-10, 
    1.368382e-10, 1.37351e-10, 1.380681e-10, 1.385833e-10, 1.389287e-10, 
    1.387169e-10, 1.389039e-10, 1.386949e-10, 1.385969e-10, 1.396851e-10, 
    1.39074e-10, 1.399908e-10, 1.399401e-10, 1.395252e-10, 1.399458e-10, 
    1.358411e-10, 1.357227e-10, 1.353117e-10, 1.356334e-10, 1.350474e-10, 
    1.353754e-10, 1.35564e-10, 1.362918e-10, 1.364517e-10, 1.366e-10, 
    1.368928e-10, 1.372687e-10, 1.379281e-10, 1.385018e-10, 1.390257e-10, 
    1.389873e-10, 1.390008e-10, 1.391178e-10, 1.388279e-10, 1.391654e-10, 
    1.39222e-10, 1.390739e-10, 1.399333e-10, 1.396878e-10, 1.39939e-10, 
    1.397792e-10, 1.357612e-10, 1.359604e-10, 1.358528e-10, 1.360552e-10, 
    1.359126e-10, 1.365466e-10, 1.367367e-10, 1.376264e-10, 1.372613e-10, 
    1.378424e-10, 1.373203e-10, 1.374128e-10, 1.378613e-10, 1.373486e-10, 
    1.384702e-10, 1.377097e-10, 1.391223e-10, 1.383628e-10, 1.391699e-10, 
    1.390234e-10, 1.39266e-10, 1.394833e-10, 1.397568e-10, 1.402613e-10, 
    1.401445e-10, 1.405664e-10, 1.362574e-10, 1.365157e-10, 1.36493e-10, 
    1.367634e-10, 1.369634e-10, 1.373968e-10, 1.380921e-10, 1.378306e-10, 
    1.383106e-10, 1.38407e-10, 1.376778e-10, 1.381255e-10, 1.366887e-10, 
    1.369208e-10, 1.367826e-10, 1.362777e-10, 1.378909e-10, 1.37063e-10, 
    1.385918e-10, 1.381433e-10, 1.394524e-10, 1.388013e-10, 1.400802e-10, 
    1.406268e-10, 1.411414e-10, 1.417428e-10, 1.366568e-10, 1.364812e-10, 
    1.367956e-10, 1.372305e-10, 1.376341e-10, 1.381706e-10, 1.382255e-10, 
    1.383261e-10, 1.385864e-10, 1.388054e-10, 1.383578e-10, 1.388603e-10, 
    1.369746e-10, 1.379627e-10, 1.364148e-10, 1.368809e-10, 1.372048e-10, 
    1.370628e-10, 1.378008e-10, 1.379747e-10, 1.386816e-10, 1.383162e-10, 
    1.404919e-10, 1.395292e-10, 1.422007e-10, 1.414541e-10, 1.364199e-10, 
    1.366562e-10, 1.374786e-10, 1.370873e-10, 1.382065e-10, 1.384819e-10, 
    1.387059e-10, 1.389922e-10, 1.390231e-10, 1.391928e-10, 1.389148e-10, 
    1.391818e-10, 1.381718e-10, 1.386231e-10, 1.373846e-10, 1.37686e-10, 
    1.375474e-10, 1.373953e-10, 1.378647e-10, 1.383649e-10, 1.383756e-10, 
    1.385359e-10, 1.389878e-10, 1.38211e-10, 1.406161e-10, 1.391306e-10, 
    1.369138e-10, 1.37369e-10, 1.37434e-10, 1.372577e-10, 1.384543e-10, 
    1.380207e-10, 1.391886e-10, 1.38873e-10, 1.393902e-10, 1.391332e-10, 
    1.390954e-10, 1.387653e-10, 1.385598e-10, 1.380406e-10, 1.376182e-10, 
    1.372833e-10, 1.373612e-10, 1.377291e-10, 1.383955e-10, 1.390259e-10, 
    1.388878e-10, 1.393509e-10, 1.381253e-10, 1.386392e-10, 1.384406e-10, 
    1.389585e-10, 1.378237e-10, 1.387899e-10, 1.375767e-10, 1.376831e-10, 
    1.380121e-10, 1.38674e-10, 1.388205e-10, 1.389769e-10, 1.388804e-10, 
    1.384124e-10, 1.383357e-10, 1.380041e-10, 1.379126e-10, 1.376599e-10, 
    1.374508e-10, 1.376419e-10, 1.378426e-10, 1.384126e-10, 1.389263e-10, 
    1.394864e-10, 1.396235e-10, 1.40278e-10, 1.397452e-10, 1.406243e-10, 
    1.398769e-10, 1.411708e-10, 1.38846e-10, 1.398549e-10, 1.380271e-10, 
    1.38224e-10, 1.385801e-10, 1.39397e-10, 1.38956e-10, 1.394718e-10, 
    1.383327e-10, 1.377418e-10, 1.375889e-10, 1.373037e-10, 1.375954e-10, 
    1.375717e-10, 1.378509e-10, 1.377612e-10, 1.384315e-10, 1.380714e-10, 
    1.390944e-10, 1.394677e-10, 1.405221e-10, 1.411685e-10, 1.418266e-10, 
    1.421171e-10, 1.422055e-10, 1.422425e-10 ;

 SOIL1N_vr =
  2.497617, 2.49761, 2.497612, 2.497606, 2.497609, 2.497606, 2.497615, 
    2.49761, 2.497613, 2.497616, 2.497596, 2.497606, 2.497586, 2.497592, 
    2.497576, 2.497587, 2.497574, 2.497576, 2.497569, 2.497571, 2.497562, 
    2.497568, 2.497557, 2.497563, 2.497562, 2.497568, 2.497604, 2.497597, 
    2.497604, 2.497603, 2.497604, 2.497609, 2.497612, 2.497617, 2.497616, 
    2.497612, 2.497603, 2.497606, 2.497598, 2.497598, 2.49759, 2.497594, 
    2.497579, 2.497583, 2.497571, 2.497574, 2.497571, 2.497572, 2.497571, 
    2.497576, 2.497574, 2.497578, 2.497593, 2.497588, 2.497602, 2.49761, 
    2.497615, 2.497619, 2.497618, 2.497617, 2.497612, 2.497607, 2.497603, 
    2.497601, 2.497598, 2.497591, 2.497587, 2.497578, 2.49758, 2.497577, 
    2.497575, 2.49757, 2.497571, 2.497569, 2.497577, 2.497572, 2.497581, 
    2.497578, 2.497598, 2.497605, 2.497608, 2.497611, 2.497618, 2.497613, 
    2.497615, 2.497611, 2.497608, 2.497609, 2.497601, 2.497604, 2.497587, 
    2.497594, 2.497575, 2.49758, 2.497574, 2.497577, 2.497572, 2.497576, 
    2.497568, 2.497566, 2.497568, 2.497563, 2.497576, 2.497571, 2.497609, 
    2.497609, 2.497608, 2.497613, 2.497613, 2.497617, 2.497613, 2.497612, 
    2.497608, 2.497605, 2.497603, 2.497598, 2.497593, 2.497585, 2.497579, 
    2.497576, 2.497578, 2.497576, 2.497578, 2.497579, 2.497567, 2.497574, 
    2.497564, 2.497565, 2.497569, 2.497564, 2.497609, 2.49761, 2.497615, 
    2.497611, 2.497618, 2.497614, 2.497612, 2.497604, 2.497602, 2.497601, 
    2.497597, 2.497593, 2.497586, 2.49758, 2.497574, 2.497575, 2.497575, 
    2.497573, 2.497576, 2.497573, 2.497572, 2.497574, 2.497565, 2.497567, 
    2.497565, 2.497566, 2.49761, 2.497608, 2.497609, 2.497607, 2.497608, 
    2.497601, 2.497599, 2.49759, 2.497594, 2.497587, 2.497593, 2.497592, 
    2.497587, 2.497593, 2.49758, 2.497589, 2.497573, 2.497581, 2.497573, 
    2.497574, 2.497572, 2.497569, 2.497566, 2.497561, 2.497562, 2.497558, 
    2.497604, 2.497602, 2.497602, 2.497599, 2.497597, 2.497592, 2.497585, 
    2.497587, 2.497582, 2.497581, 2.497589, 2.497584, 2.4976, 2.497597, 
    2.497599, 2.497604, 2.497587, 2.497596, 2.497579, 2.497584, 2.49757, 
    2.497577, 2.497563, 2.497557, 2.497551, 2.497545, 2.4976, 2.497602, 
    2.497599, 2.497594, 2.49759, 2.497584, 2.497583, 2.497582, 2.497579, 
    2.497577, 2.497582, 2.497576, 2.497597, 2.497586, 2.497603, 2.497598, 
    2.497594, 2.497596, 2.497588, 2.497586, 2.497578, 2.497582, 2.497558, 
    2.497569, 2.49754, 2.497548, 2.497603, 2.4976, 2.497591, 2.497596, 
    2.497583, 2.49758, 2.497578, 2.497575, 2.497574, 2.497573, 2.497576, 
    2.497573, 2.497584, 2.497579, 2.497592, 2.497589, 2.497591, 2.497592, 
    2.497587, 2.497581, 2.497581, 2.49758, 2.497575, 2.497583, 2.497557, 
    2.497573, 2.497597, 2.497592, 2.497592, 2.497594, 2.497581, 2.497585, 
    2.497573, 2.497576, 2.497571, 2.497573, 2.497574, 2.497577, 2.497579, 
    2.497585, 2.49759, 2.497593, 2.497592, 2.497588, 2.497581, 2.497574, 
    2.497576, 2.497571, 2.497584, 2.497579, 2.497581, 2.497575, 2.497587, 
    2.497577, 2.49759, 2.497589, 2.497585, 2.497578, 2.497576, 2.497575, 
    2.497576, 2.497581, 2.497582, 2.497586, 2.497586, 2.497589, 2.497591, 
    2.497589, 2.497587, 2.497581, 2.497576, 2.497569, 2.497568, 2.497561, 
    2.497566, 2.497557, 2.497565, 2.497551, 2.497576, 2.497565, 2.497585, 
    2.497583, 2.497579, 2.49757, 2.497575, 2.49757, 2.497582, 2.497588, 
    2.49759, 2.497593, 2.49759, 2.49759, 2.497587, 2.497588, 2.497581, 
    2.497585, 2.497574, 2.49757, 2.497558, 2.497551, 2.497544, 2.497541, 
    2.49754, 2.49754,
  2.497895, 2.497886, 2.497888, 2.497882, 2.497885, 2.497881, 2.497893, 
    2.497886, 2.49789, 2.497894, 2.497869, 2.497881, 2.497856, 2.497864, 
    2.497844, 2.497858, 2.497842, 2.497845, 2.497836, 2.497838, 2.497827, 
    2.497835, 2.497821, 2.497829, 2.497828, 2.497835, 2.497879, 2.49787, 
    2.497879, 2.497878, 2.497879, 2.497885, 2.497888, 2.497895, 2.497894, 
    2.497889, 2.497878, 2.497881, 2.497872, 2.497872, 2.497861, 2.497866, 
    2.497848, 2.497853, 2.497838, 2.497842, 2.497838, 2.49784, 2.497838, 
    2.497844, 2.497842, 2.497846, 2.497865, 2.49786, 2.497876, 2.497886, 
    2.497893, 2.497897, 2.497897, 2.497895, 2.497889, 2.497883, 2.497878, 
    2.497875, 2.497872, 2.497863, 2.497858, 2.497847, 2.497849, 2.497846, 
    2.497843, 2.497837, 2.497838, 2.497836, 2.497846, 2.497839, 2.49785, 
    2.497847, 2.497871, 2.49788, 2.497884, 2.497888, 2.497896, 2.49789, 
    2.497893, 2.497887, 2.497884, 2.497885, 2.497875, 2.497879, 2.497858, 
    2.497867, 2.497843, 2.497849, 2.497841, 2.497845, 2.497839, 2.497844, 
    2.497835, 2.497833, 2.497834, 2.497828, 2.497845, 2.497838, 2.497885, 
    2.497885, 2.497884, 2.49789, 2.49789, 2.497895, 2.49789, 2.497889, 
    2.497884, 2.497881, 2.497878, 2.497872, 2.497865, 2.497855, 2.497848, 
    2.497844, 2.497846, 2.497844, 2.497847, 2.497848, 2.497833, 2.497842, 
    2.497829, 2.49783, 2.497836, 2.49783, 2.497885, 2.497887, 2.497892, 
    2.497888, 2.497896, 2.497891, 2.497889, 2.497879, 2.497877, 2.497875, 
    2.497871, 2.497866, 2.497857, 2.497849, 2.497842, 2.497843, 2.497843, 
    2.497841, 2.497845, 2.49784, 2.49784, 2.497842, 2.49783, 2.497833, 
    2.49783, 2.497832, 2.497886, 2.497884, 2.497885, 2.497882, 2.497884, 
    2.497875, 2.497873, 2.497861, 2.497866, 2.497858, 2.497865, 2.497864, 
    2.497858, 2.497865, 2.49785, 2.49786, 2.497841, 2.497851, 2.49784, 
    2.497842, 2.497839, 2.497836, 2.497833, 2.497826, 2.497827, 2.497822, 
    2.49788, 2.497876, 2.497876, 2.497873, 2.49787, 2.497864, 2.497855, 
    2.497858, 2.497852, 2.497851, 2.49786, 2.497854, 2.497874, 2.49787, 
    2.497872, 2.497879, 2.497858, 2.497869, 2.497848, 2.497854, 2.497837, 
    2.497845, 2.497828, 2.497821, 2.497814, 2.497806, 2.497874, 2.497876, 
    2.497872, 2.497866, 2.497861, 2.497854, 2.497853, 2.497852, 2.497848, 
    2.497845, 2.497851, 2.497844, 2.49787, 2.497857, 2.497877, 2.497871, 
    2.497867, 2.497869, 2.497859, 2.497856, 2.497847, 2.497852, 2.497823, 
    2.497836, 2.4978, 2.49781, 2.497877, 2.497874, 2.497863, 2.497868, 
    2.497853, 2.497849, 2.497847, 2.497843, 2.497842, 2.49784, 2.497844, 
    2.49784, 2.497854, 2.497848, 2.497864, 2.49786, 2.497862, 2.497864, 
    2.497858, 2.497851, 2.497851, 2.497849, 2.497843, 2.497853, 2.497821, 
    2.497841, 2.497871, 2.497864, 2.497864, 2.497866, 2.49785, 2.497856, 
    2.49784, 2.497844, 2.497837, 2.497841, 2.497841, 2.497846, 2.497849, 
    2.497855, 2.497861, 2.497866, 2.497864, 2.49786, 2.497851, 2.497842, 
    2.497844, 2.497838, 2.497854, 2.497848, 2.49785, 2.497843, 2.497858, 
    2.497845, 2.497862, 2.49786, 2.497856, 2.497847, 2.497845, 2.497843, 
    2.497844, 2.49785, 2.497852, 2.497856, 2.497857, 2.497861, 2.497863, 
    2.497861, 2.497858, 2.49785, 2.497844, 2.497836, 2.497834, 2.497825, 
    2.497833, 2.497821, 2.497831, 2.497813, 2.497845, 2.497831, 2.497856, 
    2.497853, 2.497848, 2.497837, 2.497843, 2.497836, 2.497852, 2.497859, 
    2.497862, 2.497865, 2.497861, 2.497862, 2.497858, 2.497859, 2.49785, 
    2.497855, 2.497841, 2.497836, 2.497822, 2.497814, 2.497805, 2.497801, 
    2.4978, 2.497799,
  2.498021, 2.498013, 2.498014, 2.498007, 2.498011, 2.498007, 2.49802, 
    2.498012, 2.498017, 2.498021, 2.497993, 2.498007, 2.49798, 2.497988, 
    2.497967, 2.497981, 2.497964, 2.497967, 2.497957, 2.49796, 2.497947, 
    2.497956, 2.497941, 2.49795, 2.497948, 2.497956, 2.498004, 2.497995, 
    2.498005, 2.498003, 2.498004, 2.498011, 2.498015, 2.498022, 2.498021, 
    2.498015, 2.498003, 2.498007, 2.497997, 2.497997, 2.497985, 2.49799, 
    2.497971, 2.497976, 2.49796, 2.497964, 2.49796, 2.497961, 2.49796, 
    2.497966, 2.497964, 2.497969, 2.497989, 2.497983, 2.498001, 2.498012, 
    2.498019, 2.498024, 2.498024, 2.498022, 2.498015, 2.498008, 2.498003, 
    2.498, 2.497997, 2.497987, 2.497981, 2.497969, 2.497972, 2.497968, 
    2.497964, 2.497959, 2.49796, 2.497957, 2.497968, 2.497961, 2.497973, 
    2.497969, 2.497996, 2.498006, 2.49801, 2.498014, 2.498023, 2.498017, 
    2.498019, 2.498013, 2.49801, 2.498012, 2.498, 2.498004, 2.497981, 
    2.497991, 2.497965, 2.497971, 2.497963, 2.497967, 2.497961, 2.497967, 
    2.497956, 2.497954, 2.497955, 2.497949, 2.497967, 2.49796, 2.498012, 
    2.498011, 2.49801, 2.498016, 2.498016, 2.498022, 2.498017, 2.498015, 
    2.498009, 2.498006, 2.498003, 2.497996, 2.497989, 2.497978, 2.497971, 
    2.497966, 2.497969, 2.497966, 2.497969, 2.497971, 2.497955, 2.497964, 
    2.49795, 2.497951, 2.497957, 2.497951, 2.498011, 2.498013, 2.498019, 
    2.498014, 2.498023, 2.498018, 2.498015, 2.498004, 2.498002, 2.498, 
    2.497996, 2.49799, 2.49798, 2.497972, 2.497964, 2.497965, 2.497965, 
    2.497963, 2.497967, 2.497962, 2.497961, 2.497964, 2.497951, 2.497955, 
    2.497951, 2.497953, 2.498012, 2.498009, 2.498011, 2.498008, 2.49801, 
    2.498001, 2.497998, 2.497985, 2.49799, 2.497982, 2.497989, 2.497988, 
    2.497981, 2.497989, 2.497972, 2.497983, 2.497963, 2.497974, 2.497962, 
    2.497964, 2.497961, 2.497957, 2.497954, 2.497946, 2.497948, 2.497942, 
    2.498005, 2.498001, 2.498001, 2.497998, 2.497994, 2.497988, 2.497978, 
    2.497982, 2.497975, 2.497973, 2.497984, 2.497977, 2.497998, 2.497995, 
    2.497997, 2.498005, 2.497981, 2.497993, 2.497971, 2.497977, 2.497958, 
    2.497967, 2.497949, 2.497941, 2.497933, 2.497925, 2.497999, 2.498002, 
    2.497997, 2.497991, 2.497985, 2.497977, 2.497976, 2.497975, 2.497971, 
    2.497967, 2.497974, 2.497967, 2.497994, 2.49798, 2.498003, 2.497996, 
    2.497991, 2.497993, 2.497982, 2.49798, 2.497969, 2.497975, 2.497943, 
    2.497957, 2.497918, 2.497929, 2.498003, 2.497999, 2.497987, 2.497993, 
    2.497976, 2.497972, 2.497969, 2.497965, 2.497964, 2.497962, 2.497966, 
    2.497962, 2.497977, 2.49797, 2.497988, 2.497984, 2.497986, 2.497988, 
    2.497981, 2.497974, 2.497974, 2.497972, 2.497965, 2.497976, 2.497941, 
    2.497963, 2.497995, 2.497988, 2.497988, 2.49799, 2.497973, 2.497979, 
    2.497962, 2.497967, 2.497959, 2.497963, 2.497963, 2.497968, 2.497971, 
    2.497979, 2.497985, 2.49799, 2.497989, 2.497983, 2.497973, 2.497964, 
    2.497966, 2.497959, 2.497977, 2.49797, 2.497973, 2.497965, 2.497982, 
    2.497968, 2.497986, 2.497984, 2.497979, 2.497969, 2.497967, 2.497965, 
    2.497966, 2.497973, 2.497974, 2.497979, 2.497981, 2.497984, 2.497987, 
    2.497985, 2.497982, 2.497973, 2.497966, 2.497957, 2.497956, 2.497946, 
    2.497954, 2.497941, 2.497952, 2.497933, 2.497967, 2.497952, 2.497979, 
    2.497976, 2.497971, 2.497959, 2.497965, 2.497958, 2.497974, 2.497983, 
    2.497985, 2.497989, 2.497985, 2.497986, 2.497982, 2.497983, 2.497973, 
    2.497978, 2.497963, 2.497958, 2.497942, 2.497933, 2.497923, 2.497919, 
    2.497918, 2.497917,
  2.49812, 2.498111, 2.498112, 2.498105, 2.498109, 2.498105, 2.498118, 
    2.49811, 2.498115, 2.498119, 2.498091, 2.498105, 2.498077, 2.498086, 
    2.498064, 2.498078, 2.498061, 2.498064, 2.498054, 2.498057, 2.498044, 
    2.498053, 2.498038, 2.498046, 2.498045, 2.498053, 2.498102, 2.498093, 
    2.498103, 2.498101, 2.498102, 2.498109, 2.498113, 2.49812, 2.498119, 
    2.498113, 2.498101, 2.498105, 2.498094, 2.498095, 2.498083, 2.498088, 
    2.498068, 2.498074, 2.498057, 2.498061, 2.498057, 2.498058, 2.498057, 
    2.498063, 2.498061, 2.498066, 2.498087, 2.498081, 2.498099, 2.49811, 
    2.498117, 2.498123, 2.498122, 2.498121, 2.498113, 2.498106, 2.498101, 
    2.498098, 2.498095, 2.498084, 2.498079, 2.498067, 2.498069, 2.498065, 
    2.498062, 2.498056, 2.498057, 2.498054, 2.498065, 2.498058, 2.49807, 
    2.498067, 2.498094, 2.498104, 2.498108, 2.498112, 2.498121, 2.498115, 
    2.498117, 2.498111, 2.498108, 2.49811, 2.498098, 2.498102, 2.498079, 
    2.498089, 2.498062, 2.498068, 2.49806, 2.498065, 2.498058, 2.498064, 
    2.498053, 2.498051, 2.498052, 2.498046, 2.498064, 2.498057, 2.49811, 
    2.498109, 2.498108, 2.498114, 2.498115, 2.49812, 2.498115, 2.498113, 
    2.498107, 2.498104, 2.498101, 2.498094, 2.498086, 2.498076, 2.498068, 
    2.498063, 2.498066, 2.498063, 2.498066, 2.498068, 2.498052, 2.498061, 
    2.498047, 2.498048, 2.498054, 2.498048, 2.498109, 2.498111, 2.498117, 
    2.498112, 2.498121, 2.498116, 2.498113, 2.498102, 2.4981, 2.498098, 
    2.498093, 2.498088, 2.498078, 2.498069, 2.498061, 2.498062, 2.498062, 
    2.49806, 2.498064, 2.498059, 2.498059, 2.498061, 2.498048, 2.498051, 
    2.498048, 2.49805, 2.49811, 2.498107, 2.498109, 2.498106, 2.498108, 
    2.498098, 2.498096, 2.498082, 2.498088, 2.498079, 2.498087, 2.498085, 
    2.498079, 2.498086, 2.49807, 2.498081, 2.49806, 2.498071, 2.498059, 
    2.498061, 2.498058, 2.498055, 2.49805, 2.498043, 2.498045, 2.498038, 
    2.498103, 2.498099, 2.498099, 2.498095, 2.498092, 2.498086, 2.498075, 
    2.498079, 2.498072, 2.498071, 2.498081, 2.498075, 2.498096, 2.498093, 
    2.498095, 2.498102, 2.498078, 2.498091, 2.498068, 2.498075, 2.498055, 
    2.498065, 2.498046, 2.498037, 2.49803, 2.498021, 2.498097, 2.4981, 
    2.498095, 2.498088, 2.498082, 2.498074, 2.498073, 2.498072, 2.498068, 
    2.498065, 2.498071, 2.498064, 2.498092, 2.498077, 2.498101, 2.498093, 
    2.498089, 2.498091, 2.49808, 2.498077, 2.498066, 2.498072, 2.498039, 
    2.498054, 2.498014, 2.498025, 2.4981, 2.498097, 2.498085, 2.498091, 
    2.498074, 2.49807, 2.498066, 2.498062, 2.498061, 2.498059, 2.498063, 
    2.498059, 2.498074, 2.498067, 2.498086, 2.498081, 2.498084, 2.498086, 
    2.498079, 2.498071, 2.498071, 2.498069, 2.498062, 2.498074, 2.498038, 
    2.49806, 2.498093, 2.498086, 2.498085, 2.498088, 2.49807, 2.498076, 
    2.498059, 2.498064, 2.498056, 2.49806, 2.49806, 2.498065, 2.498068, 
    2.498076, 2.498082, 2.498087, 2.498086, 2.498081, 2.498071, 2.498061, 
    2.498064, 2.498056, 2.498075, 2.498067, 2.49807, 2.498062, 2.498079, 
    2.498065, 2.498083, 2.498081, 2.498076, 2.498067, 2.498065, 2.498062, 
    2.498064, 2.49807, 2.498072, 2.498077, 2.498078, 2.498082, 2.498085, 
    2.498082, 2.498079, 2.49807, 2.498063, 2.498055, 2.498052, 2.498043, 
    2.498051, 2.498038, 2.498049, 2.498029, 2.498064, 2.498049, 2.498076, 
    2.498073, 2.498068, 2.498056, 2.498062, 2.498055, 2.498072, 2.49808, 
    2.498083, 2.498087, 2.498083, 2.498083, 2.498079, 2.49808, 2.49807, 
    2.498076, 2.49806, 2.498055, 2.498039, 2.498029, 2.498019, 2.498015, 
    2.498014, 2.498013,
  2.498258, 2.49825, 2.498252, 2.498245, 2.498249, 2.498244, 2.498256, 
    2.49825, 2.498254, 2.498257, 2.498232, 2.498245, 2.498219, 2.498227, 
    2.498207, 2.498221, 2.498205, 2.498208, 2.498199, 2.498201, 2.498189, 
    2.498197, 2.498183, 2.498191, 2.49819, 2.498198, 2.498242, 2.498234, 
    2.498243, 2.498242, 2.498242, 2.498249, 2.498252, 2.498259, 2.498258, 
    2.498252, 2.498241, 2.498245, 2.498235, 2.498235, 2.498224, 2.498229, 
    2.498211, 2.498216, 2.498201, 2.498205, 2.498201, 2.498202, 2.498201, 
    2.498207, 2.498204, 2.498209, 2.498228, 2.498223, 2.49824, 2.49825, 
    2.498256, 2.498261, 2.49826, 2.498259, 2.498252, 2.498246, 2.498242, 
    2.498239, 2.498235, 2.498226, 2.498221, 2.49821, 2.498212, 2.498209, 
    2.498205, 2.4982, 2.498201, 2.498198, 2.498209, 2.498202, 2.498213, 
    2.49821, 2.498235, 2.498244, 2.498248, 2.498251, 2.49826, 2.498254, 
    2.498256, 2.498251, 2.498247, 2.498249, 2.498238, 2.498243, 2.498221, 
    2.49823, 2.498206, 2.498212, 2.498204, 2.498208, 2.498202, 2.498207, 
    2.498197, 2.498195, 2.498197, 2.498191, 2.498208, 2.498201, 2.498249, 
    2.498249, 2.498247, 2.498253, 2.498254, 2.498259, 2.498254, 2.498252, 
    2.498247, 2.498244, 2.498241, 2.498235, 2.498228, 2.498218, 2.498211, 
    2.498206, 2.498209, 2.498207, 2.49821, 2.498211, 2.498196, 2.498204, 
    2.498192, 2.498193, 2.498198, 2.498193, 2.498249, 2.49825, 2.498256, 
    2.498251, 2.498259, 2.498255, 2.498252, 2.498242, 2.49824, 2.498238, 
    2.498234, 2.498229, 2.49822, 2.498212, 2.498205, 2.498206, 2.498205, 
    2.498204, 2.498208, 2.498203, 2.498202, 2.498204, 2.498193, 2.498196, 
    2.498193, 2.498195, 2.49825, 2.498247, 2.498248, 2.498246, 2.498248, 
    2.498239, 2.498236, 2.498224, 2.498229, 2.498221, 2.498228, 2.498227, 
    2.498221, 2.498228, 2.498213, 2.498223, 2.498204, 2.498214, 2.498203, 
    2.498205, 2.498202, 2.498199, 2.498195, 2.498188, 2.49819, 2.498184, 
    2.498243, 2.498239, 2.49824, 2.498236, 2.498233, 2.498227, 2.498218, 
    2.498221, 2.498215, 2.498214, 2.498224, 2.498217, 2.498237, 2.498234, 
    2.498236, 2.498243, 2.498221, 2.498232, 2.498211, 2.498217, 2.498199, 
    2.498208, 2.498191, 2.498183, 2.498176, 2.498168, 2.498237, 2.49824, 
    2.498235, 2.49823, 2.498224, 2.498217, 2.498216, 2.498215, 2.498211, 
    2.498208, 2.498214, 2.498207, 2.498233, 2.49822, 2.498241, 2.498234, 
    2.49823, 2.498232, 2.498222, 2.498219, 2.49821, 2.498215, 2.498185, 
    2.498198, 2.498162, 2.498172, 2.498241, 2.498237, 2.498226, 2.498232, 
    2.498216, 2.498213, 2.498209, 2.498206, 2.498205, 2.498203, 2.498207, 
    2.498203, 2.498217, 2.498211, 2.498228, 2.498223, 2.498225, 2.498227, 
    2.498221, 2.498214, 2.498214, 2.498212, 2.498206, 2.498216, 2.498183, 
    2.498204, 2.498234, 2.498228, 2.498227, 2.498229, 2.498213, 2.498219, 
    2.498203, 2.498207, 2.4982, 2.498204, 2.498204, 2.498209, 2.498211, 
    2.498219, 2.498224, 2.498229, 2.498228, 2.498223, 2.498214, 2.498205, 
    2.498207, 2.498201, 2.498217, 2.49821, 2.498213, 2.498206, 2.498222, 
    2.498208, 2.498225, 2.498224, 2.498219, 2.49821, 2.498208, 2.498206, 
    2.498207, 2.498214, 2.498214, 2.498219, 2.49822, 2.498224, 2.498227, 
    2.498224, 2.498221, 2.498214, 2.498206, 2.498199, 2.498197, 2.498188, 
    2.498195, 2.498183, 2.498194, 2.498176, 2.498208, 2.498194, 2.498219, 
    2.498216, 2.498211, 2.4982, 2.498206, 2.498199, 2.498214, 2.498223, 
    2.498225, 2.498229, 2.498225, 2.498225, 2.498221, 2.498222, 2.498213, 
    2.498218, 2.498204, 2.498199, 2.498185, 2.498176, 2.498167, 2.498163, 
    2.498162, 2.498161,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  6.002251e-08, 6.028716e-08, 6.023572e-08, 6.044917e-08, 6.033077e-08, 
    6.047054e-08, 6.007617e-08, 6.029767e-08, 6.015627e-08, 6.004634e-08, 
    6.086344e-08, 6.04587e-08, 6.128394e-08, 6.102579e-08, 6.167433e-08, 
    6.124377e-08, 6.176116e-08, 6.166193e-08, 6.196064e-08, 6.187506e-08, 
    6.225714e-08, 6.200014e-08, 6.245521e-08, 6.219577e-08, 6.223635e-08, 
    6.199166e-08, 6.054017e-08, 6.081304e-08, 6.052399e-08, 6.05629e-08, 
    6.054545e-08, 6.033321e-08, 6.022625e-08, 6.000229e-08, 6.004295e-08, 
    6.020745e-08, 6.05804e-08, 6.045381e-08, 6.077289e-08, 6.076569e-08, 
    6.112093e-08, 6.096076e-08, 6.155789e-08, 6.138817e-08, 6.187864e-08, 
    6.175529e-08, 6.187284e-08, 6.18372e-08, 6.187331e-08, 6.16924e-08, 
    6.17699e-08, 6.161072e-08, 6.099075e-08, 6.117294e-08, 6.062957e-08, 
    6.030285e-08, 6.008588e-08, 5.993191e-08, 5.995368e-08, 5.999517e-08, 
    6.020841e-08, 6.040892e-08, 6.056172e-08, 6.066394e-08, 6.076465e-08, 
    6.106949e-08, 6.123086e-08, 6.15922e-08, 6.1527e-08, 6.163746e-08, 
    6.174302e-08, 6.19202e-08, 6.189104e-08, 6.196911e-08, 6.163456e-08, 
    6.185689e-08, 6.148986e-08, 6.159024e-08, 6.079198e-08, 6.048796e-08, 
    6.035871e-08, 6.02456e-08, 5.997042e-08, 6.016045e-08, 6.008553e-08, 
    6.026377e-08, 6.037703e-08, 6.032101e-08, 6.066673e-08, 6.053232e-08, 
    6.124043e-08, 6.093541e-08, 6.17307e-08, 6.154038e-08, 6.177632e-08, 
    6.165593e-08, 6.186221e-08, 6.167656e-08, 6.199816e-08, 6.206822e-08, 
    6.202034e-08, 6.22042e-08, 6.166627e-08, 6.187283e-08, 6.031944e-08, 
    6.032858e-08, 6.037114e-08, 6.018405e-08, 6.01726e-08, 6.000118e-08, 
    6.015372e-08, 6.021867e-08, 6.03836e-08, 6.048114e-08, 6.057387e-08, 
    6.077776e-08, 6.100547e-08, 6.132392e-08, 6.155273e-08, 6.17061e-08, 
    6.161205e-08, 6.169508e-08, 6.160226e-08, 6.155877e-08, 6.204197e-08, 
    6.177063e-08, 6.217776e-08, 6.215524e-08, 6.197097e-08, 6.215777e-08, 
    6.0335e-08, 6.028242e-08, 6.009991e-08, 6.024274e-08, 5.99825e-08, 
    6.012817e-08, 6.021192e-08, 6.053512e-08, 6.060615e-08, 6.067199e-08, 
    6.080204e-08, 6.096895e-08, 6.126176e-08, 6.151654e-08, 6.174916e-08, 
    6.173212e-08, 6.173811e-08, 6.179008e-08, 6.166136e-08, 6.181121e-08, 
    6.183635e-08, 6.17706e-08, 6.215222e-08, 6.20432e-08, 6.215475e-08, 
    6.208377e-08, 6.029951e-08, 6.038797e-08, 6.034017e-08, 6.043005e-08, 
    6.036673e-08, 6.06483e-08, 6.073272e-08, 6.112779e-08, 6.096567e-08, 
    6.122371e-08, 6.099188e-08, 6.103296e-08, 6.123211e-08, 6.100441e-08, 
    6.150249e-08, 6.116479e-08, 6.179209e-08, 6.145482e-08, 6.181322e-08, 
    6.174815e-08, 6.18559e-08, 6.19524e-08, 6.207384e-08, 6.229785e-08, 
    6.224597e-08, 6.243333e-08, 6.051985e-08, 6.063458e-08, 6.062449e-08, 
    6.074456e-08, 6.083337e-08, 6.102586e-08, 6.133459e-08, 6.121849e-08, 
    6.143164e-08, 6.147443e-08, 6.115062e-08, 6.134942e-08, 6.071137e-08, 
    6.081444e-08, 6.075308e-08, 6.052889e-08, 6.124524e-08, 6.087759e-08, 
    6.15565e-08, 6.135733e-08, 6.193864e-08, 6.164952e-08, 6.221742e-08, 
    6.246017e-08, 6.268869e-08, 6.295571e-08, 6.06972e-08, 6.061924e-08, 
    6.075884e-08, 6.095198e-08, 6.11312e-08, 6.136947e-08, 6.139386e-08, 
    6.143849e-08, 6.155413e-08, 6.165134e-08, 6.14526e-08, 6.167571e-08, 
    6.083833e-08, 6.127715e-08, 6.058976e-08, 6.079673e-08, 6.094059e-08, 
    6.08775e-08, 6.120523e-08, 6.128247e-08, 6.159637e-08, 6.143411e-08, 
    6.240025e-08, 6.197277e-08, 6.315906e-08, 6.282752e-08, 6.059201e-08, 
    6.069694e-08, 6.106216e-08, 6.088839e-08, 6.138538e-08, 6.150772e-08, 
    6.160718e-08, 6.173431e-08, 6.174804e-08, 6.182337e-08, 6.169994e-08, 
    6.18185e-08, 6.136998e-08, 6.157041e-08, 6.102042e-08, 6.115427e-08, 
    6.10927e-08, 6.102515e-08, 6.123363e-08, 6.145572e-08, 6.146048e-08, 
    6.153169e-08, 6.173236e-08, 6.13874e-08, 6.245539e-08, 6.179577e-08, 
    6.081137e-08, 6.101348e-08, 6.104237e-08, 6.096408e-08, 6.149546e-08, 
    6.130291e-08, 6.182153e-08, 6.168137e-08, 6.191103e-08, 6.17969e-08, 
    6.178011e-08, 6.163354e-08, 6.154228e-08, 6.131173e-08, 6.112416e-08, 
    6.097543e-08, 6.101001e-08, 6.11734e-08, 6.146931e-08, 6.174928e-08, 
    6.168795e-08, 6.189358e-08, 6.134935e-08, 6.157754e-08, 6.148934e-08, 
    6.171933e-08, 6.121541e-08, 6.164448e-08, 6.110573e-08, 6.115297e-08, 
    6.129908e-08, 6.159301e-08, 6.165806e-08, 6.172749e-08, 6.168465e-08, 
    6.147683e-08, 6.144278e-08, 6.129554e-08, 6.125487e-08, 6.114269e-08, 
    6.10498e-08, 6.113466e-08, 6.122379e-08, 6.147692e-08, 6.170504e-08, 
    6.195377e-08, 6.201465e-08, 6.230526e-08, 6.206869e-08, 6.245907e-08, 
    6.212714e-08, 6.270175e-08, 6.166937e-08, 6.211741e-08, 6.130574e-08, 
    6.139318e-08, 6.155132e-08, 6.191407e-08, 6.171825e-08, 6.194727e-08, 
    6.144145e-08, 6.117902e-08, 6.111114e-08, 6.098447e-08, 6.111404e-08, 
    6.11035e-08, 6.122748e-08, 6.118764e-08, 6.148532e-08, 6.132542e-08, 
    6.177969e-08, 6.194546e-08, 6.241369e-08, 6.270072e-08, 6.299293e-08, 
    6.312194e-08, 6.316121e-08, 6.317762e-08 ;

 SOIL1_HR_S3 =
  7.123147e-10, 7.154565e-10, 7.148458e-10, 7.1738e-10, 7.159743e-10, 
    7.176336e-10, 7.129517e-10, 7.155812e-10, 7.139026e-10, 7.125976e-10, 
    7.222981e-10, 7.174931e-10, 7.272904e-10, 7.242255e-10, 7.319253e-10, 
    7.268134e-10, 7.329562e-10, 7.31778e-10, 7.353245e-10, 7.343085e-10, 
    7.388447e-10, 7.357934e-10, 7.411965e-10, 7.381162e-10, 7.38598e-10, 
    7.356927e-10, 7.184602e-10, 7.216998e-10, 7.182682e-10, 7.187301e-10, 
    7.185229e-10, 7.160033e-10, 7.147334e-10, 7.120746e-10, 7.125573e-10, 
    7.145102e-10, 7.189379e-10, 7.174349e-10, 7.212231e-10, 7.211375e-10, 
    7.253551e-10, 7.234535e-10, 7.305428e-10, 7.285278e-10, 7.343509e-10, 
    7.328864e-10, 7.342821e-10, 7.338589e-10, 7.342876e-10, 7.321397e-10, 
    7.330599e-10, 7.311701e-10, 7.238096e-10, 7.259726e-10, 7.195216e-10, 
    7.156428e-10, 7.13067e-10, 7.112391e-10, 7.114975e-10, 7.119901e-10, 
    7.145217e-10, 7.16902e-10, 7.187161e-10, 7.199296e-10, 7.211253e-10, 
    7.247443e-10, 7.266602e-10, 7.309502e-10, 7.301761e-10, 7.314875e-10, 
    7.327407e-10, 7.348444e-10, 7.344982e-10, 7.35425e-10, 7.314531e-10, 
    7.340927e-10, 7.297352e-10, 7.309269e-10, 7.214498e-10, 7.178405e-10, 
    7.163059e-10, 7.149632e-10, 7.116962e-10, 7.139522e-10, 7.130629e-10, 
    7.151789e-10, 7.165234e-10, 7.158585e-10, 7.199628e-10, 7.18367e-10, 
    7.267738e-10, 7.231525e-10, 7.325945e-10, 7.30335e-10, 7.331361e-10, 
    7.317068e-10, 7.341558e-10, 7.319517e-10, 7.3577e-10, 7.366017e-10, 
    7.360333e-10, 7.382162e-10, 7.318295e-10, 7.34282e-10, 7.158398e-10, 
    7.159482e-10, 7.164535e-10, 7.142324e-10, 7.140966e-10, 7.120614e-10, 
    7.138724e-10, 7.146435e-10, 7.166014e-10, 7.177594e-10, 7.188603e-10, 
    7.212809e-10, 7.239843e-10, 7.27765e-10, 7.304815e-10, 7.323023e-10, 
    7.311858e-10, 7.321715e-10, 7.310696e-10, 7.305532e-10, 7.362901e-10, 
    7.330685e-10, 7.379023e-10, 7.376348e-10, 7.35447e-10, 7.376649e-10, 
    7.160244e-10, 7.154004e-10, 7.132335e-10, 7.149292e-10, 7.118398e-10, 
    7.13569e-10, 7.145633e-10, 7.184003e-10, 7.192434e-10, 7.200252e-10, 
    7.215692e-10, 7.235508e-10, 7.27027e-10, 7.30052e-10, 7.328136e-10, 
    7.326112e-10, 7.326825e-10, 7.332994e-10, 7.317713e-10, 7.335503e-10, 
    7.338488e-10, 7.330682e-10, 7.37599e-10, 7.363046e-10, 7.376291e-10, 
    7.367864e-10, 7.156032e-10, 7.166533e-10, 7.160859e-10, 7.171529e-10, 
    7.164012e-10, 7.197439e-10, 7.207462e-10, 7.254365e-10, 7.235118e-10, 
    7.265753e-10, 7.238229e-10, 7.243106e-10, 7.26675e-10, 7.239717e-10, 
    7.29885e-10, 7.258757e-10, 7.333233e-10, 7.293192e-10, 7.335743e-10, 
    7.328017e-10, 7.34081e-10, 7.352267e-10, 7.366684e-10, 7.39328e-10, 
    7.387122e-10, 7.409366e-10, 7.182189e-10, 7.195811e-10, 7.194612e-10, 
    7.208867e-10, 7.219411e-10, 7.242263e-10, 7.278917e-10, 7.265134e-10, 
    7.290439e-10, 7.295519e-10, 7.257074e-10, 7.280678e-10, 7.204927e-10, 
    7.217164e-10, 7.209879e-10, 7.183263e-10, 7.268308e-10, 7.224661e-10, 
    7.305263e-10, 7.281616e-10, 7.350633e-10, 7.316308e-10, 7.383731e-10, 
    7.412553e-10, 7.439685e-10, 7.471388e-10, 7.203245e-10, 7.19399e-10, 
    7.210563e-10, 7.233492e-10, 7.25477e-10, 7.283058e-10, 7.285953e-10, 
    7.291253e-10, 7.304981e-10, 7.316523e-10, 7.292927e-10, 7.319417e-10, 
    7.22e-10, 7.272097e-10, 7.19049e-10, 7.215061e-10, 7.232141e-10, 
    7.224649e-10, 7.263559e-10, 7.272729e-10, 7.309996e-10, 7.290731e-10, 
    7.405438e-10, 7.354685e-10, 7.495532e-10, 7.456168e-10, 7.190756e-10, 
    7.203214e-10, 7.246573e-10, 7.225943e-10, 7.284947e-10, 7.299472e-10, 
    7.31128e-10, 7.326373e-10, 7.328004e-10, 7.336947e-10, 7.322292e-10, 
    7.336368e-10, 7.283119e-10, 7.306914e-10, 7.241618e-10, 7.257509e-10, 
    7.250199e-10, 7.24218e-10, 7.26693e-10, 7.293298e-10, 7.293863e-10, 
    7.302318e-10, 7.326141e-10, 7.285186e-10, 7.411986e-10, 7.333671e-10, 
    7.216799e-10, 7.240795e-10, 7.244224e-10, 7.234928e-10, 7.298015e-10, 
    7.275155e-10, 7.336729e-10, 7.320088e-10, 7.347355e-10, 7.333805e-10, 
    7.331812e-10, 7.31441e-10, 7.303575e-10, 7.276204e-10, 7.253934e-10, 
    7.236277e-10, 7.240383e-10, 7.259779e-10, 7.294911e-10, 7.328151e-10, 
    7.320869e-10, 7.345283e-10, 7.280669e-10, 7.307761e-10, 7.297289e-10, 
    7.324595e-10, 7.264767e-10, 7.315708e-10, 7.251746e-10, 7.257354e-10, 
    7.274702e-10, 7.309597e-10, 7.317321e-10, 7.325563e-10, 7.320478e-10, 
    7.295804e-10, 7.291762e-10, 7.274281e-10, 7.269453e-10, 7.256133e-10, 
    7.245106e-10, 7.255181e-10, 7.265762e-10, 7.295815e-10, 7.322899e-10, 
    7.352429e-10, 7.359657e-10, 7.394161e-10, 7.366073e-10, 7.412422e-10, 
    7.373013e-10, 7.441235e-10, 7.318663e-10, 7.371857e-10, 7.275492e-10, 
    7.285872e-10, 7.304648e-10, 7.347716e-10, 7.324467e-10, 7.351658e-10, 
    7.291604e-10, 7.260448e-10, 7.252389e-10, 7.23735e-10, 7.252732e-10, 
    7.251481e-10, 7.266201e-10, 7.261471e-10, 7.296813e-10, 7.277828e-10, 
    7.331761e-10, 7.351443e-10, 7.407034e-10, 7.441113e-10, 7.475808e-10, 
    7.491125e-10, 7.495788e-10, 7.497737e-10 ;

 SOIL2C =
  5.783962, 5.783968, 5.783967, 5.783972, 5.783969, 5.783972, 5.783963, 
    5.783968, 5.783965, 5.783962, 5.783981, 5.783972, 5.78399, 5.783985, 
    5.783999, 5.78399, 5.784001, 5.783999, 5.784006, 5.784004, 5.784013, 
    5.784007, 5.784017, 5.784011, 5.784012, 5.784007, 5.783974, 5.78398, 
    5.783973, 5.783974, 5.783974, 5.783969, 5.783967, 5.783961, 5.783962, 
    5.783966, 5.783975, 5.783972, 5.783979, 5.783979, 5.783987, 5.783983, 
    5.783997, 5.783993, 5.784004, 5.784001, 5.784004, 5.784003, 5.784004, 
    5.784, 5.784002, 5.783998, 5.783984, 5.783988, 5.783976, 5.783968, 
    5.783963, 5.78396, 5.78396, 5.783961, 5.783966, 5.783971, 5.783974, 
    5.783977, 5.783979, 5.783986, 5.783989, 5.783998, 5.783996, 5.783998, 
    5.784001, 5.784005, 5.784004, 5.784006, 5.783998, 5.784004, 5.783995, 
    5.783998, 5.783979, 5.783972, 5.783969, 5.783967, 5.783961, 5.783965, 
    5.783963, 5.783967, 5.78397, 5.783968, 5.783977, 5.783974, 5.783989, 
    5.783983, 5.784001, 5.783997, 5.784002, 5.783999, 5.784004, 5.783999, 
    5.784007, 5.784009, 5.784008, 5.784011, 5.783999, 5.784004, 5.783968, 
    5.783969, 5.78397, 5.783966, 5.783965, 5.783961, 5.783965, 5.783967, 
    5.78397, 5.783972, 5.783975, 5.783979, 5.783984, 5.783991, 5.783997, 
    5.784, 5.783998, 5.784, 5.783998, 5.783997, 5.784008, 5.784002, 5.784011, 
    5.78401, 5.784006, 5.78401, 5.783969, 5.783968, 5.783964, 5.783967, 
    5.783961, 5.783964, 5.783966, 5.783974, 5.783975, 5.783977, 5.783979, 
    5.783983, 5.78399, 5.783996, 5.784001, 5.784001, 5.784001, 5.784002, 
    5.783999, 5.784003, 5.784003, 5.784002, 5.78401, 5.784008, 5.78401, 
    5.784009, 5.783968, 5.78397, 5.783969, 5.783971, 5.78397, 5.783976, 
    5.783978, 5.783987, 5.783983, 5.783989, 5.783984, 5.783985, 5.783989, 
    5.783984, 5.783996, 5.783988, 5.784002, 5.783995, 5.784003, 5.784001, 
    5.784004, 5.784006, 5.784009, 5.784014, 5.784012, 5.784017, 5.783973, 
    5.783976, 5.783976, 5.783978, 5.78398, 5.783985, 5.783992, 5.783989, 
    5.783994, 5.783995, 5.783988, 5.783992, 5.783978, 5.78398, 5.783978, 
    5.783973, 5.78399, 5.783981, 5.783997, 5.783992, 5.784006, 5.783999, 
    5.784012, 5.784018, 5.784023, 5.784029, 5.783977, 5.783976, 5.783978, 
    5.783983, 5.783987, 5.783993, 5.783993, 5.783994, 5.783997, 5.783999, 
    5.783995, 5.783999, 5.78398, 5.78399, 5.783975, 5.783979, 5.783983, 
    5.783981, 5.783989, 5.78399, 5.783998, 5.783994, 5.784016, 5.784006, 
    5.784033, 5.784026, 5.783975, 5.783977, 5.783986, 5.783982, 5.783993, 
    5.783996, 5.783998, 5.784001, 5.784001, 5.784003, 5.784, 5.784003, 
    5.783993, 5.783997, 5.783985, 5.783988, 5.783986, 5.783985, 5.783989, 
    5.783995, 5.783995, 5.783996, 5.784001, 5.783993, 5.784017, 5.784002, 
    5.78398, 5.783985, 5.783985, 5.783983, 5.783996, 5.783991, 5.784003, 
    5.783999, 5.784005, 5.784002, 5.784002, 5.783998, 5.783997, 5.783991, 
    5.783987, 5.783984, 5.783984, 5.783988, 5.783995, 5.784001, 5.784, 
    5.784005, 5.783992, 5.783998, 5.783995, 5.784, 5.783989, 5.783999, 
    5.783987, 5.783988, 5.783991, 5.783998, 5.783999, 5.784001, 5.784, 
    5.783995, 5.783994, 5.783991, 5.78399, 5.783988, 5.783985, 5.783987, 
    5.783989, 5.783995, 5.784, 5.784006, 5.784007, 5.784014, 5.784009, 
    5.784018, 5.78401, 5.784023, 5.783999, 5.784009, 5.783991, 5.783993, 
    5.783997, 5.784005, 5.784, 5.784006, 5.783994, 5.783988, 5.783987, 
    5.783984, 5.783987, 5.783987, 5.783989, 5.783988, 5.783995, 5.783991, 
    5.784002, 5.784006, 5.784016, 5.784023, 5.784029, 5.784032, 5.784033, 
    5.784034 ;

 SOIL2C_TO_SOIL1C =
  1.06187e-09, 1.066555e-09, 1.065645e-09, 1.069424e-09, 1.067327e-09, 
    1.069802e-09, 1.06282e-09, 1.066741e-09, 1.064238e-09, 1.062292e-09, 
    1.076758e-09, 1.069592e-09, 1.084203e-09, 1.079632e-09, 1.091115e-09, 
    1.083491e-09, 1.092652e-09, 1.090895e-09, 1.096183e-09, 1.094668e-09, 
    1.101433e-09, 1.096883e-09, 1.10494e-09, 1.100346e-09, 1.101065e-09, 
    1.096733e-09, 1.071035e-09, 1.075866e-09, 1.070748e-09, 1.071437e-09, 
    1.071128e-09, 1.067371e-09, 1.065477e-09, 1.061512e-09, 1.062232e-09, 
    1.065144e-09, 1.071747e-09, 1.069506e-09, 1.075155e-09, 1.075027e-09, 
    1.081317e-09, 1.078481e-09, 1.089053e-09, 1.086048e-09, 1.094732e-09, 
    1.092548e-09, 1.094629e-09, 1.093998e-09, 1.094637e-09, 1.091434e-09, 
    1.092807e-09, 1.089988e-09, 1.079012e-09, 1.082238e-09, 1.072617e-09, 
    1.066833e-09, 1.062992e-09, 1.060266e-09, 1.060651e-09, 1.061386e-09, 
    1.065161e-09, 1.068711e-09, 1.071416e-09, 1.073226e-09, 1.075009e-09, 
    1.080406e-09, 1.083263e-09, 1.08966e-09, 1.088506e-09, 1.090462e-09, 
    1.09233e-09, 1.095468e-09, 1.094951e-09, 1.096333e-09, 1.09041e-09, 
    1.094347e-09, 1.087848e-09, 1.089626e-09, 1.075493e-09, 1.07011e-09, 
    1.067822e-09, 1.06582e-09, 1.060948e-09, 1.064312e-09, 1.062986e-09, 
    1.066141e-09, 1.068146e-09, 1.067155e-09, 1.073275e-09, 1.070896e-09, 
    1.083432e-09, 1.078032e-09, 1.092112e-09, 1.088743e-09, 1.09292e-09, 
    1.090789e-09, 1.094441e-09, 1.091154e-09, 1.096848e-09, 1.098088e-09, 
    1.09724e-09, 1.100496e-09, 1.090972e-09, 1.094629e-09, 1.067127e-09, 
    1.067289e-09, 1.068042e-09, 1.06473e-09, 1.064527e-09, 1.061492e-09, 
    1.064193e-09, 1.065343e-09, 1.068263e-09, 1.06999e-09, 1.071631e-09, 
    1.075241e-09, 1.079273e-09, 1.084911e-09, 1.088961e-09, 1.091677e-09, 
    1.090012e-09, 1.091482e-09, 1.089838e-09, 1.089068e-09, 1.097623e-09, 
    1.092819e-09, 1.100027e-09, 1.099629e-09, 1.096366e-09, 1.099674e-09, 
    1.067402e-09, 1.066472e-09, 1.06324e-09, 1.065769e-09, 1.061162e-09, 
    1.063741e-09, 1.065223e-09, 1.070945e-09, 1.072203e-09, 1.073369e-09, 
    1.075671e-09, 1.078626e-09, 1.08381e-09, 1.088321e-09, 1.092439e-09, 
    1.092137e-09, 1.092244e-09, 1.093164e-09, 1.090885e-09, 1.093538e-09, 
    1.093983e-09, 1.092819e-09, 1.099575e-09, 1.097645e-09, 1.09962e-09, 
    1.098363e-09, 1.066774e-09, 1.06834e-09, 1.067494e-09, 1.069085e-09, 
    1.067964e-09, 1.072949e-09, 1.074444e-09, 1.081438e-09, 1.078568e-09, 
    1.083136e-09, 1.079032e-09, 1.079759e-09, 1.083285e-09, 1.079254e-09, 
    1.088072e-09, 1.082093e-09, 1.093199e-09, 1.087228e-09, 1.093574e-09, 
    1.092421e-09, 1.094329e-09, 1.096037e-09, 1.098187e-09, 1.102154e-09, 
    1.101235e-09, 1.104552e-09, 1.070675e-09, 1.072706e-09, 1.072528e-09, 
    1.074653e-09, 1.076226e-09, 1.079633e-09, 1.085099e-09, 1.083044e-09, 
    1.086818e-09, 1.087575e-09, 1.081842e-09, 1.085362e-09, 1.074066e-09, 
    1.075891e-09, 1.074804e-09, 1.070835e-09, 1.083517e-09, 1.077009e-09, 
    1.089028e-09, 1.085502e-09, 1.095794e-09, 1.090675e-09, 1.10073e-09, 
    1.105027e-09, 1.109073e-09, 1.113801e-09, 1.073815e-09, 1.072435e-09, 
    1.074906e-09, 1.078326e-09, 1.081499e-09, 1.085717e-09, 1.086149e-09, 
    1.086939e-09, 1.088986e-09, 1.090707e-09, 1.087189e-09, 1.091139e-09, 
    1.076313e-09, 1.084083e-09, 1.071913e-09, 1.075577e-09, 1.078124e-09, 
    1.077007e-09, 1.082809e-09, 1.084177e-09, 1.089734e-09, 1.086861e-09, 
    1.103966e-09, 1.096398e-09, 1.117401e-09, 1.111531e-09, 1.071952e-09, 
    1.07381e-09, 1.080276e-09, 1.0772e-09, 1.085999e-09, 1.088165e-09, 
    1.089926e-09, 1.092176e-09, 1.092419e-09, 1.093753e-09, 1.091568e-09, 
    1.093667e-09, 1.085726e-09, 1.089275e-09, 1.079537e-09, 1.081907e-09, 
    1.080817e-09, 1.079621e-09, 1.083312e-09, 1.087244e-09, 1.087328e-09, 
    1.088589e-09, 1.092142e-09, 1.086034e-09, 1.104943e-09, 1.093265e-09, 
    1.075836e-09, 1.079414e-09, 1.079926e-09, 1.07854e-09, 1.087948e-09, 
    1.084539e-09, 1.093721e-09, 1.091239e-09, 1.095305e-09, 1.093285e-09, 
    1.092987e-09, 1.090392e-09, 1.088777e-09, 1.084695e-09, 1.081374e-09, 
    1.078741e-09, 1.079353e-09, 1.082246e-09, 1.087485e-09, 1.092441e-09, 
    1.091356e-09, 1.094996e-09, 1.085361e-09, 1.089401e-09, 1.087839e-09, 
    1.091911e-09, 1.082989e-09, 1.090586e-09, 1.081048e-09, 1.081884e-09, 
    1.084471e-09, 1.089675e-09, 1.090826e-09, 1.092056e-09, 1.091297e-09, 
    1.087618e-09, 1.087015e-09, 1.084408e-09, 1.083688e-09, 1.081702e-09, 
    1.080057e-09, 1.08156e-09, 1.083138e-09, 1.087619e-09, 1.091658e-09, 
    1.096062e-09, 1.09714e-09, 1.102285e-09, 1.098096e-09, 1.105008e-09, 
    1.099131e-09, 1.109305e-09, 1.091026e-09, 1.098959e-09, 1.084589e-09, 
    1.086137e-09, 1.088937e-09, 1.095359e-09, 1.091892e-09, 1.095947e-09, 
    1.086991e-09, 1.082345e-09, 1.081144e-09, 1.078901e-09, 1.081195e-09, 
    1.081008e-09, 1.083203e-09, 1.082498e-09, 1.087768e-09, 1.084937e-09, 
    1.09298e-09, 1.095915e-09, 1.104205e-09, 1.109286e-09, 1.11446e-09, 
    1.116744e-09, 1.117439e-09, 1.11773e-09 ;

 SOIL2C_TO_SOIL3C =
  7.584785e-11, 7.618253e-11, 7.611747e-11, 7.638741e-11, 7.623768e-11, 
    7.641443e-11, 7.591571e-11, 7.619581e-11, 7.601701e-11, 7.587799e-11, 
    7.691128e-11, 7.639946e-11, 7.744306e-11, 7.711659e-11, 7.793675e-11, 
    7.739225e-11, 7.804656e-11, 7.792107e-11, 7.829882e-11, 7.819059e-11, 
    7.867377e-11, 7.834876e-11, 7.892426e-11, 7.859617e-11, 7.864748e-11, 
    7.833804e-11, 7.650248e-11, 7.684756e-11, 7.648203e-11, 7.653123e-11, 
    7.650915e-11, 7.624076e-11, 7.61055e-11, 7.582229e-11, 7.58737e-11, 
    7.608172e-11, 7.655336e-11, 7.639327e-11, 7.679678e-11, 7.678767e-11, 
    7.723691e-11, 7.703436e-11, 7.778949e-11, 7.757486e-11, 7.819511e-11, 
    7.803912e-11, 7.818778e-11, 7.814271e-11, 7.818837e-11, 7.795959e-11, 
    7.805761e-11, 7.78563e-11, 7.707229e-11, 7.730269e-11, 7.661553e-11, 
    7.620236e-11, 7.592799e-11, 7.573329e-11, 7.576081e-11, 7.581329e-11, 
    7.608295e-11, 7.63365e-11, 7.652973e-11, 7.665899e-11, 7.678636e-11, 
    7.717185e-11, 7.737593e-11, 7.783289e-11, 7.775043e-11, 7.789012e-11, 
    7.80236e-11, 7.824768e-11, 7.821081e-11, 7.830953e-11, 7.788645e-11, 
    7.816762e-11, 7.770346e-11, 7.783041e-11, 7.682092e-11, 7.643646e-11, 
    7.6273e-11, 7.612998e-11, 7.578198e-11, 7.602229e-11, 7.592756e-11, 
    7.615295e-11, 7.629617e-11, 7.622535e-11, 7.666253e-11, 7.649256e-11, 
    7.738803e-11, 7.700231e-11, 7.800803e-11, 7.776736e-11, 7.806572e-11, 
    7.791347e-11, 7.817434e-11, 7.793956e-11, 7.834627e-11, 7.843486e-11, 
    7.837431e-11, 7.860683e-11, 7.792655e-11, 7.818778e-11, 7.622335e-11, 
    7.623491e-11, 7.628873e-11, 7.605214e-11, 7.603766e-11, 7.582087e-11, 
    7.601378e-11, 7.609592e-11, 7.630448e-11, 7.642784e-11, 7.65451e-11, 
    7.680294e-11, 7.70909e-11, 7.749361e-11, 7.778296e-11, 7.797692e-11, 
    7.785798e-11, 7.796298e-11, 7.78456e-11, 7.779059e-11, 7.840167e-11, 
    7.805852e-11, 7.857339e-11, 7.85449e-11, 7.831187e-11, 7.854811e-11, 
    7.624302e-11, 7.617654e-11, 7.594572e-11, 7.612636e-11, 7.579726e-11, 
    7.598146e-11, 7.608738e-11, 7.649609e-11, 7.658591e-11, 7.666918e-11, 
    7.683365e-11, 7.704472e-11, 7.7415e-11, 7.773721e-11, 7.803137e-11, 
    7.800981e-11, 7.801741e-11, 7.808312e-11, 7.792034e-11, 7.810984e-11, 
    7.814163e-11, 7.805848e-11, 7.854108e-11, 7.840322e-11, 7.85443e-11, 
    7.845453e-11, 7.619815e-11, 7.631001e-11, 7.624957e-11, 7.636323e-11, 
    7.628315e-11, 7.663922e-11, 7.674598e-11, 7.724559e-11, 7.704056e-11, 
    7.736689e-11, 7.707372e-11, 7.712566e-11, 7.737751e-11, 7.708956e-11, 
    7.771944e-11, 7.729237e-11, 7.808566e-11, 7.765915e-11, 7.811239e-11, 
    7.80301e-11, 7.816636e-11, 7.82884e-11, 7.844196e-11, 7.872526e-11, 
    7.865966e-11, 7.889658e-11, 7.647678e-11, 7.662187e-11, 7.660911e-11, 
    7.676095e-11, 7.687326e-11, 7.711668e-11, 7.75071e-11, 7.736029e-11, 
    7.762984e-11, 7.768395e-11, 7.727445e-11, 7.752586e-11, 7.671899e-11, 
    7.684933e-11, 7.677173e-11, 7.648822e-11, 7.739411e-11, 7.692918e-11, 
    7.778773e-11, 7.753585e-11, 7.827099e-11, 7.790538e-11, 7.862355e-11, 
    7.893053e-11, 7.921952e-11, 7.955719e-11, 7.670107e-11, 7.660248e-11, 
    7.677901e-11, 7.702325e-11, 7.72499e-11, 7.755122e-11, 7.758205e-11, 
    7.76385e-11, 7.778473e-11, 7.790767e-11, 7.765634e-11, 7.79385e-11, 
    7.687954e-11, 7.743447e-11, 7.65652e-11, 7.682693e-11, 7.700886e-11, 
    7.692906e-11, 7.734351e-11, 7.74412e-11, 7.783815e-11, 7.763296e-11, 
    7.885475e-11, 7.831416e-11, 7.981435e-11, 7.939508e-11, 7.656803e-11, 
    7.670074e-11, 7.716259e-11, 7.694283e-11, 7.757134e-11, 7.772605e-11, 
    7.785182e-11, 7.80126e-11, 7.802996e-11, 7.812522e-11, 7.796912e-11, 
    7.811906e-11, 7.755186e-11, 7.780532e-11, 7.71098e-11, 7.727908e-11, 
    7.720121e-11, 7.711579e-11, 7.737943e-11, 7.766029e-11, 7.766631e-11, 
    7.775637e-11, 7.801013e-11, 7.757388e-11, 7.892449e-11, 7.809033e-11, 
    7.684544e-11, 7.710103e-11, 7.713757e-11, 7.703855e-11, 7.771053e-11, 
    7.746704e-11, 7.81229e-11, 7.794564e-11, 7.823608e-11, 7.809176e-11, 
    7.807052e-11, 7.788516e-11, 7.776976e-11, 7.74782e-11, 7.724099e-11, 
    7.705291e-11, 7.709665e-11, 7.730325e-11, 7.767748e-11, 7.803153e-11, 
    7.795397e-11, 7.821401e-11, 7.752576e-11, 7.781434e-11, 7.77028e-11, 
    7.799365e-11, 7.735639e-11, 7.789899e-11, 7.721769e-11, 7.727743e-11, 
    7.746221e-11, 7.78339e-11, 7.791617e-11, 7.800397e-11, 7.794979e-11, 
    7.768698e-11, 7.764393e-11, 7.745772e-11, 7.74063e-11, 7.726442e-11, 
    7.714696e-11, 7.725428e-11, 7.736698e-11, 7.768709e-11, 7.797558e-11, 
    7.829013e-11, 7.836712e-11, 7.873463e-11, 7.843545e-11, 7.892913e-11, 
    7.850938e-11, 7.923603e-11, 7.793047e-11, 7.849706e-11, 7.747062e-11, 
    7.75812e-11, 7.778118e-11, 7.823992e-11, 7.799228e-11, 7.828191e-11, 
    7.764225e-11, 7.731037e-11, 7.722453e-11, 7.706434e-11, 7.72282e-11, 
    7.721487e-11, 7.737166e-11, 7.732127e-11, 7.769772e-11, 7.749551e-11, 
    7.806998e-11, 7.827963e-11, 7.887175e-11, 7.923473e-11, 7.960427e-11, 
    7.976741e-11, 7.981708e-11, 7.983784e-11 ;

 SOIL2C_vr =
  20.00596, 20.00598, 20.00598, 20.00599, 20.00598, 20.00599, 20.00597, 
    20.00598, 20.00597, 20.00596, 20.00601, 20.00599, 20.00604, 20.00602, 
    20.00606, 20.00604, 20.00607, 20.00606, 20.00608, 20.00607, 20.0061, 
    20.00608, 20.00611, 20.0061, 20.0061, 20.00608, 20.00599, 20.00601, 
    20.00599, 20.00599, 20.00599, 20.00598, 20.00597, 20.00596, 20.00596, 
    20.00597, 20.006, 20.00599, 20.00601, 20.00601, 20.00603, 20.00602, 
    20.00606, 20.00605, 20.00607, 20.00607, 20.00607, 20.00607, 20.00607, 
    20.00607, 20.00607, 20.00606, 20.00602, 20.00603, 20.006, 20.00598, 
    20.00597, 20.00596, 20.00596, 20.00596, 20.00597, 20.00599, 20.00599, 
    20.006, 20.00601, 20.00603, 20.00604, 20.00606, 20.00605, 20.00606, 
    20.00607, 20.00608, 20.00608, 20.00608, 20.00606, 20.00607, 20.00605, 
    20.00606, 20.00601, 20.00599, 20.00598, 20.00598, 20.00596, 20.00597, 
    20.00597, 20.00598, 20.00598, 20.00598, 20.006, 20.00599, 20.00604, 
    20.00602, 20.00607, 20.00606, 20.00607, 20.00606, 20.00607, 20.00606, 
    20.00608, 20.00609, 20.00608, 20.0061, 20.00606, 20.00607, 20.00598, 
    20.00598, 20.00598, 20.00597, 20.00597, 20.00596, 20.00597, 20.00597, 
    20.00598, 20.00599, 20.006, 20.00601, 20.00602, 20.00604, 20.00606, 
    20.00607, 20.00606, 20.00607, 20.00606, 20.00606, 20.00609, 20.00607, 
    20.00609, 20.00609, 20.00608, 20.00609, 20.00598, 20.00598, 20.00597, 
    20.00598, 20.00596, 20.00597, 20.00597, 20.00599, 20.006, 20.006, 
    20.00601, 20.00602, 20.00604, 20.00605, 20.00607, 20.00607, 20.00607, 
    20.00607, 20.00606, 20.00607, 20.00607, 20.00607, 20.00609, 20.00609, 
    20.00609, 20.00609, 20.00598, 20.00599, 20.00598, 20.00599, 20.00598, 
    20.006, 20.00601, 20.00603, 20.00602, 20.00603, 20.00602, 20.00602, 
    20.00604, 20.00602, 20.00605, 20.00603, 20.00607, 20.00605, 20.00607, 
    20.00607, 20.00607, 20.00608, 20.00609, 20.0061, 20.0061, 20.00611, 
    20.00599, 20.006, 20.006, 20.00601, 20.00601, 20.00602, 20.00604, 
    20.00603, 20.00605, 20.00605, 20.00603, 20.00604, 20.006, 20.00601, 
    20.00601, 20.00599, 20.00604, 20.00601, 20.00606, 20.00604, 20.00608, 
    20.00606, 20.0061, 20.00611, 20.00612, 20.00614, 20.006, 20.006, 
    20.00601, 20.00602, 20.00603, 20.00604, 20.00605, 20.00605, 20.00606, 
    20.00606, 20.00605, 20.00606, 20.00601, 20.00604, 20.006, 20.00601, 
    20.00602, 20.00601, 20.00603, 20.00604, 20.00606, 20.00605, 20.00611, 
    20.00608, 20.00615, 20.00613, 20.006, 20.006, 20.00603, 20.00602, 
    20.00605, 20.00605, 20.00606, 20.00607, 20.00607, 20.00607, 20.00607, 
    20.00607, 20.00604, 20.00606, 20.00602, 20.00603, 20.00603, 20.00602, 
    20.00604, 20.00605, 20.00605, 20.00605, 20.00607, 20.00605, 20.00611, 
    20.00607, 20.00601, 20.00602, 20.00603, 20.00602, 20.00605, 20.00604, 
    20.00607, 20.00606, 20.00608, 20.00607, 20.00607, 20.00606, 20.00606, 
    20.00604, 20.00603, 20.00602, 20.00602, 20.00603, 20.00605, 20.00607, 
    20.00606, 20.00608, 20.00604, 20.00606, 20.00605, 20.00607, 20.00603, 
    20.00606, 20.00603, 20.00603, 20.00604, 20.00606, 20.00606, 20.00607, 
    20.00606, 20.00605, 20.00605, 20.00604, 20.00604, 20.00603, 20.00603, 
    20.00603, 20.00603, 20.00605, 20.00607, 20.00608, 20.00608, 20.0061, 
    20.00609, 20.00611, 20.00609, 20.00613, 20.00606, 20.00609, 20.00604, 
    20.00605, 20.00606, 20.00608, 20.00607, 20.00608, 20.00605, 20.00603, 
    20.00603, 20.00602, 20.00603, 20.00603, 20.00604, 20.00603, 20.00605, 
    20.00604, 20.00607, 20.00608, 20.00611, 20.00613, 20.00614, 20.00615, 
    20.00615, 20.00616,
  20.00538, 20.0054, 20.0054, 20.00541, 20.00541, 20.00542, 20.00539, 
    20.0054, 20.00539, 20.00538, 20.00545, 20.00542, 20.00548, 20.00546, 
    20.00551, 20.00548, 20.00552, 20.00551, 20.00553, 20.00553, 20.00556, 
    20.00554, 20.00557, 20.00555, 20.00555, 20.00554, 20.00542, 20.00544, 
    20.00542, 20.00542, 20.00542, 20.00541, 20.0054, 20.00538, 20.00538, 
    20.0054, 20.00543, 20.00542, 20.00544, 20.00544, 20.00547, 20.00546, 
    20.0055, 20.00549, 20.00553, 20.00552, 20.00553, 20.00552, 20.00553, 
    20.00551, 20.00552, 20.0055, 20.00546, 20.00547, 20.00543, 20.0054, 
    20.00539, 20.00537, 20.00538, 20.00538, 20.0054, 20.00541, 20.00542, 
    20.00543, 20.00544, 20.00546, 20.00548, 20.0055, 20.0055, 20.00551, 
    20.00552, 20.00553, 20.00553, 20.00553, 20.00551, 20.00552, 20.0055, 
    20.0055, 20.00544, 20.00542, 20.00541, 20.0054, 20.00538, 20.00539, 
    20.00539, 20.0054, 20.00541, 20.00541, 20.00543, 20.00542, 20.00548, 
    20.00545, 20.00551, 20.0055, 20.00552, 20.00551, 20.00553, 20.00551, 
    20.00554, 20.00554, 20.00554, 20.00555, 20.00551, 20.00553, 20.00541, 
    20.00541, 20.00541, 20.0054, 20.00539, 20.00538, 20.00539, 20.0054, 
    20.00541, 20.00542, 20.00542, 20.00544, 20.00546, 20.00548, 20.0055, 
    20.00551, 20.0055, 20.00551, 20.0055, 20.0055, 20.00554, 20.00552, 
    20.00555, 20.00555, 20.00553, 20.00555, 20.00541, 20.0054, 20.00539, 
    20.0054, 20.00538, 20.00539, 20.0054, 20.00542, 20.00543, 20.00543, 
    20.00544, 20.00546, 20.00548, 20.0055, 20.00552, 20.00551, 20.00552, 
    20.00552, 20.00551, 20.00552, 20.00552, 20.00552, 20.00555, 20.00554, 
    20.00555, 20.00554, 20.0054, 20.00541, 20.00541, 20.00541, 20.00541, 
    20.00543, 20.00544, 20.00547, 20.00546, 20.00548, 20.00546, 20.00546, 
    20.00548, 20.00546, 20.0055, 20.00547, 20.00552, 20.00549, 20.00552, 
    20.00552, 20.00552, 20.00553, 20.00554, 20.00556, 20.00555, 20.00557, 
    20.00542, 20.00543, 20.00543, 20.00544, 20.00545, 20.00546, 20.00548, 
    20.00548, 20.00549, 20.0055, 20.00547, 20.00549, 20.00544, 20.00544, 
    20.00544, 20.00542, 20.00548, 20.00545, 20.0055, 20.00549, 20.00553, 
    20.00551, 20.00555, 20.00557, 20.00559, 20.00561, 20.00543, 20.00543, 
    20.00544, 20.00546, 20.00547, 20.00549, 20.00549, 20.00549, 20.0055, 
    20.00551, 20.00549, 20.00551, 20.00545, 20.00548, 20.00543, 20.00544, 
    20.00545, 20.00545, 20.00547, 20.00548, 20.0055, 20.00549, 20.00557, 
    20.00553, 20.00562, 20.0056, 20.00543, 20.00543, 20.00546, 20.00545, 
    20.00549, 20.0055, 20.0055, 20.00551, 20.00552, 20.00552, 20.00551, 
    20.00552, 20.00549, 20.0055, 20.00546, 20.00547, 20.00546, 20.00546, 
    20.00548, 20.00549, 20.00549, 20.0055, 20.00551, 20.00549, 20.00557, 
    20.00552, 20.00544, 20.00546, 20.00546, 20.00546, 20.0055, 20.00548, 
    20.00552, 20.00551, 20.00553, 20.00552, 20.00552, 20.00551, 20.0055, 
    20.00548, 20.00547, 20.00546, 20.00546, 20.00547, 20.0055, 20.00552, 
    20.00551, 20.00553, 20.00549, 20.0055, 20.0055, 20.00551, 20.00547, 
    20.00551, 20.00547, 20.00547, 20.00548, 20.0055, 20.00551, 20.00551, 
    20.00551, 20.0055, 20.00549, 20.00548, 20.00548, 20.00547, 20.00546, 
    20.00547, 20.00548, 20.0055, 20.00551, 20.00553, 20.00554, 20.00556, 
    20.00554, 20.00557, 20.00554, 20.00559, 20.00551, 20.00554, 20.00548, 
    20.00549, 20.0055, 20.00553, 20.00551, 20.00553, 20.00549, 20.00547, 
    20.00547, 20.00546, 20.00547, 20.00547, 20.00548, 20.00547, 20.0055, 
    20.00548, 20.00552, 20.00553, 20.00557, 20.00559, 20.00561, 20.00562, 
    20.00562, 20.00563,
  20.00506, 20.00508, 20.00508, 20.00509, 20.00508, 20.0051, 20.00506, 
    20.00508, 20.00507, 20.00506, 20.00513, 20.00509, 20.00517, 20.00514, 
    20.0052, 20.00516, 20.00521, 20.0052, 20.00522, 20.00521, 20.00525, 
    20.00523, 20.00526, 20.00524, 20.00525, 20.00522, 20.0051, 20.00513, 
    20.0051, 20.0051, 20.0051, 20.00508, 20.00508, 20.00506, 20.00506, 
    20.00507, 20.00511, 20.00509, 20.00512, 20.00512, 20.00515, 20.00514, 
    20.00519, 20.00517, 20.00521, 20.00521, 20.00521, 20.00521, 20.00521, 
    20.0052, 20.00521, 20.00519, 20.00514, 20.00516, 20.00511, 20.00508, 
    20.00506, 20.00505, 20.00505, 20.00506, 20.00507, 20.00509, 20.0051, 
    20.00511, 20.00512, 20.00515, 20.00516, 20.00519, 20.00519, 20.0052, 
    20.0052, 20.00522, 20.00522, 20.00522, 20.00519, 20.00521, 20.00518, 
    20.00519, 20.00512, 20.0051, 20.00509, 20.00508, 20.00505, 20.00507, 
    20.00506, 20.00508, 20.00509, 20.00508, 20.00511, 20.0051, 20.00516, 
    20.00513, 20.0052, 20.00519, 20.00521, 20.0052, 20.00521, 20.0052, 
    20.00523, 20.00523, 20.00523, 20.00524, 20.0052, 20.00521, 20.00508, 
    20.00508, 20.00509, 20.00507, 20.00507, 20.00506, 20.00507, 20.00508, 
    20.00509, 20.0051, 20.0051, 20.00512, 20.00514, 20.00517, 20.00519, 
    20.0052, 20.00519, 20.0052, 20.00519, 20.00519, 20.00523, 20.00521, 
    20.00524, 20.00524, 20.00522, 20.00524, 20.00508, 20.00508, 20.00506, 
    20.00508, 20.00505, 20.00507, 20.00507, 20.0051, 20.00511, 20.00511, 
    20.00513, 20.00514, 20.00516, 20.00518, 20.00521, 20.0052, 20.0052, 
    20.00521, 20.0052, 20.00521, 20.00521, 20.00521, 20.00524, 20.00523, 
    20.00524, 20.00523, 20.00508, 20.00509, 20.00508, 20.00509, 20.00509, 
    20.00511, 20.00512, 20.00515, 20.00514, 20.00516, 20.00514, 20.00514, 
    20.00516, 20.00514, 20.00518, 20.00516, 20.00521, 20.00518, 20.00521, 
    20.0052, 20.00521, 20.00522, 20.00523, 20.00525, 20.00525, 20.00526, 
    20.0051, 20.00511, 20.00511, 20.00512, 20.00513, 20.00514, 20.00517, 
    20.00516, 20.00518, 20.00518, 20.00515, 20.00517, 20.00512, 20.00513, 
    20.00512, 20.0051, 20.00516, 20.00513, 20.00519, 20.00517, 20.00522, 
    20.0052, 20.00524, 20.00526, 20.00528, 20.00531, 20.00512, 20.00511, 
    20.00512, 20.00514, 20.00515, 20.00517, 20.00517, 20.00518, 20.00519, 
    20.0052, 20.00518, 20.0052, 20.00513, 20.00517, 20.00511, 20.00512, 
    20.00514, 20.00513, 20.00516, 20.00517, 20.00519, 20.00518, 20.00526, 
    20.00522, 20.00532, 20.00529, 20.00511, 20.00512, 20.00515, 20.00513, 
    20.00517, 20.00518, 20.00519, 20.0052, 20.0052, 20.00521, 20.0052, 
    20.00521, 20.00517, 20.00519, 20.00514, 20.00515, 20.00515, 20.00514, 
    20.00516, 20.00518, 20.00518, 20.00519, 20.0052, 20.00517, 20.00526, 
    20.00521, 20.00513, 20.00514, 20.00514, 20.00514, 20.00518, 20.00517, 
    20.00521, 20.0052, 20.00522, 20.00521, 20.00521, 20.00519, 20.00519, 
    20.00517, 20.00515, 20.00514, 20.00514, 20.00516, 20.00518, 20.00521, 
    20.0052, 20.00522, 20.00517, 20.00519, 20.00518, 20.0052, 20.00516, 
    20.0052, 20.00515, 20.00515, 20.00517, 20.00519, 20.0052, 20.0052, 
    20.0052, 20.00518, 20.00518, 20.00517, 20.00516, 20.00515, 20.00515, 
    20.00515, 20.00516, 20.00518, 20.0052, 20.00522, 20.00523, 20.00525, 
    20.00523, 20.00526, 20.00524, 20.00529, 20.0052, 20.00524, 20.00517, 
    20.00517, 20.00519, 20.00522, 20.0052, 20.00522, 20.00518, 20.00516, 
    20.00515, 20.00514, 20.00515, 20.00515, 20.00516, 20.00516, 20.00518, 
    20.00517, 20.00521, 20.00522, 20.00526, 20.00529, 20.00531, 20.00532, 
    20.00532, 20.00533,
  20.00481, 20.00483, 20.00483, 20.00484, 20.00483, 20.00485, 20.00481, 
    20.00483, 20.00482, 20.00481, 20.00488, 20.00484, 20.00492, 20.00489, 
    20.00495, 20.00491, 20.00496, 20.00495, 20.00497, 20.00497, 20.005, 
    20.00498, 20.00502, 20.00499, 20.005, 20.00498, 20.00485, 20.00488, 
    20.00485, 20.00485, 20.00485, 20.00483, 20.00483, 20.0048, 20.00481, 
    20.00482, 20.00486, 20.00484, 20.00487, 20.00487, 20.0049, 20.00489, 
    20.00494, 20.00492, 20.00497, 20.00496, 20.00497, 20.00496, 20.00497, 
    20.00495, 20.00496, 20.00494, 20.00489, 20.00491, 20.00486, 20.00483, 
    20.00481, 20.0048, 20.0048, 20.0048, 20.00482, 20.00484, 20.00485, 
    20.00486, 20.00487, 20.0049, 20.00491, 20.00494, 20.00494, 20.00495, 
    20.00496, 20.00497, 20.00497, 20.00497, 20.00495, 20.00496, 20.00493, 
    20.00494, 20.00487, 20.00485, 20.00484, 20.00483, 20.0048, 20.00482, 
    20.00481, 20.00483, 20.00484, 20.00483, 20.00486, 20.00485, 20.00491, 
    20.00489, 20.00495, 20.00494, 20.00496, 20.00495, 20.00496, 20.00495, 
    20.00498, 20.00498, 20.00498, 20.005, 20.00495, 20.00497, 20.00483, 
    20.00483, 20.00484, 20.00482, 20.00482, 20.0048, 20.00482, 20.00482, 
    20.00484, 20.00485, 20.00485, 20.00487, 20.00489, 20.00492, 20.00494, 
    20.00495, 20.00494, 20.00495, 20.00494, 20.00494, 20.00498, 20.00496, 
    20.00499, 20.00499, 20.00497, 20.00499, 20.00483, 20.00483, 20.00481, 
    20.00483, 20.0048, 20.00482, 20.00482, 20.00485, 20.00486, 20.00486, 
    20.00488, 20.00489, 20.00491, 20.00494, 20.00496, 20.00496, 20.00496, 
    20.00496, 20.00495, 20.00496, 20.00496, 20.00496, 20.00499, 20.00498, 
    20.00499, 20.00498, 20.00483, 20.00484, 20.00484, 20.00484, 20.00484, 
    20.00486, 20.00487, 20.0049, 20.00489, 20.00491, 20.00489, 20.00489, 
    20.00491, 20.00489, 20.00493, 20.00491, 20.00496, 20.00493, 20.00496, 
    20.00496, 20.00496, 20.00497, 20.00498, 20.005, 20.005, 20.00501, 
    20.00485, 20.00486, 20.00486, 20.00487, 20.00488, 20.00489, 20.00492, 
    20.00491, 20.00493, 20.00493, 20.0049, 20.00492, 20.00487, 20.00488, 
    20.00487, 20.00485, 20.00491, 20.00488, 20.00494, 20.00492, 20.00497, 
    20.00495, 20.005, 20.00502, 20.00504, 20.00506, 20.00487, 20.00486, 
    20.00487, 20.00489, 20.0049, 20.00492, 20.00492, 20.00493, 20.00494, 
    20.00495, 20.00493, 20.00495, 20.00488, 20.00492, 20.00486, 20.00487, 
    20.00489, 20.00488, 20.00491, 20.00492, 20.00494, 20.00493, 20.00501, 
    20.00497, 20.00508, 20.00505, 20.00486, 20.00487, 20.0049, 20.00488, 
    20.00492, 20.00493, 20.00494, 20.00496, 20.00496, 20.00496, 20.00495, 
    20.00496, 20.00492, 20.00494, 20.00489, 20.0049, 20.0049, 20.00489, 
    20.00491, 20.00493, 20.00493, 20.00494, 20.00496, 20.00492, 20.00502, 
    20.00496, 20.00488, 20.00489, 20.00489, 20.00489, 20.00493, 20.00492, 
    20.00496, 20.00495, 20.00497, 20.00496, 20.00496, 20.00495, 20.00494, 
    20.00492, 20.0049, 20.00489, 20.00489, 20.00491, 20.00493, 20.00496, 
    20.00495, 20.00497, 20.00492, 20.00494, 20.00493, 20.00495, 20.00491, 
    20.00495, 20.0049, 20.0049, 20.00492, 20.00494, 20.00495, 20.00495, 
    20.00495, 20.00493, 20.00493, 20.00492, 20.00491, 20.0049, 20.0049, 
    20.0049, 20.00491, 20.00493, 20.00495, 20.00497, 20.00498, 20.005, 
    20.00498, 20.00502, 20.00499, 20.00504, 20.00495, 20.00499, 20.00492, 
    20.00492, 20.00494, 20.00497, 20.00495, 20.00497, 20.00493, 20.00491, 
    20.0049, 20.00489, 20.0049, 20.0049, 20.00491, 20.00491, 20.00493, 
    20.00492, 20.00496, 20.00497, 20.00501, 20.00504, 20.00506, 20.00507, 
    20.00508, 20.00508,
  20.00426, 20.00428, 20.00428, 20.00429, 20.00428, 20.0043, 20.00426, 
    20.00428, 20.00427, 20.00426, 20.00432, 20.00429, 20.00436, 20.00434, 
    20.00438, 20.00435, 20.00439, 20.00438, 20.00441, 20.0044, 20.00443, 
    20.00441, 20.00444, 20.00443, 20.00443, 20.00441, 20.0043, 20.00432, 
    20.0043, 20.0043, 20.0043, 20.00428, 20.00428, 20.00426, 20.00426, 
    20.00427, 20.0043, 20.00429, 20.00432, 20.00432, 20.00434, 20.00433, 
    20.00438, 20.00436, 20.0044, 20.00439, 20.0044, 20.0044, 20.0044, 
    20.00439, 20.00439, 20.00438, 20.00433, 20.00435, 20.00431, 20.00428, 
    20.00427, 20.00426, 20.00426, 20.00426, 20.00427, 20.00429, 20.0043, 
    20.00431, 20.00432, 20.00434, 20.00435, 20.00438, 20.00437, 20.00438, 
    20.00439, 20.0044, 20.0044, 20.00441, 20.00438, 20.0044, 20.00437, 
    20.00438, 20.00432, 20.0043, 20.00429, 20.00428, 20.00426, 20.00427, 
    20.00427, 20.00428, 20.00429, 20.00428, 20.00431, 20.0043, 20.00435, 
    20.00433, 20.00439, 20.00438, 20.00439, 20.00438, 20.0044, 20.00438, 
    20.00441, 20.00442, 20.00441, 20.00443, 20.00438, 20.0044, 20.00428, 
    20.00428, 20.00429, 20.00427, 20.00427, 20.00426, 20.00427, 20.00428, 
    20.00429, 20.0043, 20.0043, 20.00432, 20.00434, 20.00436, 20.00438, 
    20.00439, 20.00438, 20.00439, 20.00438, 20.00438, 20.00441, 20.00439, 
    20.00442, 20.00442, 20.00441, 20.00442, 20.00428, 20.00428, 20.00427, 
    20.00428, 20.00426, 20.00427, 20.00428, 20.0043, 20.0043, 20.00431, 
    20.00432, 20.00433, 20.00435, 20.00437, 20.00439, 20.00439, 20.00439, 
    20.00439, 20.00438, 20.0044, 20.0044, 20.00439, 20.00442, 20.00441, 
    20.00442, 20.00442, 20.00428, 20.00429, 20.00429, 20.00429, 20.00429, 
    20.00431, 20.00431, 20.00434, 20.00433, 20.00435, 20.00433, 20.00434, 
    20.00435, 20.00434, 20.00437, 20.00435, 20.00439, 20.00437, 20.0044, 
    20.00439, 20.0044, 20.00441, 20.00442, 20.00443, 20.00443, 20.00444, 
    20.0043, 20.00431, 20.00431, 20.00431, 20.00432, 20.00434, 20.00436, 
    20.00435, 20.00437, 20.00437, 20.00434, 20.00436, 20.00431, 20.00432, 
    20.00432, 20.0043, 20.00435, 20.00433, 20.00438, 20.00436, 20.00441, 
    20.00438, 20.00443, 20.00444, 20.00446, 20.00448, 20.00431, 20.00431, 
    20.00432, 20.00433, 20.00434, 20.00436, 20.00436, 20.00437, 20.00438, 
    20.00438, 20.00437, 20.00438, 20.00432, 20.00435, 20.0043, 20.00432, 
    20.00433, 20.00433, 20.00435, 20.00436, 20.00438, 20.00437, 20.00444, 
    20.00441, 20.0045, 20.00447, 20.0043, 20.00431, 20.00434, 20.00433, 
    20.00436, 20.00437, 20.00438, 20.00439, 20.00439, 20.0044, 20.00439, 
    20.0044, 20.00436, 20.00438, 20.00434, 20.00435, 20.00434, 20.00434, 
    20.00435, 20.00437, 20.00437, 20.00438, 20.00439, 20.00436, 20.00444, 
    20.00439, 20.00432, 20.00434, 20.00434, 20.00433, 20.00437, 20.00436, 
    20.0044, 20.00438, 20.0044, 20.00439, 20.00439, 20.00438, 20.00438, 
    20.00436, 20.00434, 20.00433, 20.00434, 20.00435, 20.00437, 20.00439, 
    20.00439, 20.0044, 20.00436, 20.00438, 20.00437, 20.00439, 20.00435, 
    20.00438, 20.00434, 20.00435, 20.00436, 20.00438, 20.00438, 20.00439, 
    20.00439, 20.00437, 20.00437, 20.00436, 20.00435, 20.00434, 20.00434, 
    20.00434, 20.00435, 20.00437, 20.00439, 20.00441, 20.00441, 20.00443, 
    20.00442, 20.00444, 20.00442, 20.00446, 20.00438, 20.00442, 20.00436, 
    20.00436, 20.00438, 20.0044, 20.00439, 20.00441, 20.00437, 20.00435, 
    20.00434, 20.00433, 20.00434, 20.00434, 20.00435, 20.00435, 20.00437, 
    20.00436, 20.00439, 20.00441, 20.00444, 20.00446, 20.00448, 20.00449, 
    20.0045, 20.0045,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258147, 0.5258152, 0.5258151, 0.5258156, 0.5258154, 0.5258157, 
    0.5258148, 0.5258153, 0.525815, 0.5258148, 0.5258164, 0.5258156, 
    0.5258173, 0.5258168, 0.5258181, 0.5258172, 0.5258183, 0.5258181, 
    0.5258187, 0.5258185, 0.5258194, 0.5258188, 0.5258198, 0.5258192, 
    0.5258193, 0.5258188, 0.5258158, 0.5258164, 0.5258157, 0.5258158, 
    0.5258158, 0.5258154, 0.5258151, 0.5258147, 0.5258148, 0.5258151, 
    0.5258158, 0.5258156, 0.5258163, 0.5258163, 0.525817, 0.5258167, 
    0.5258179, 0.5258176, 0.5258186, 0.5258183, 0.5258185, 0.5258185, 
    0.5258185, 0.5258182, 0.5258183, 0.525818, 0.5258167, 0.5258171, 
    0.525816, 0.5258153, 0.5258148, 0.5258145, 0.5258146, 0.5258147, 
    0.5258151, 0.5258155, 0.5258158, 0.525816, 0.5258163, 0.5258169, 
    0.5258172, 0.525818, 0.5258178, 0.525818, 0.5258183, 0.5258186, 
    0.5258186, 0.5258188, 0.525818, 0.5258185, 0.5258178, 0.525818, 
    0.5258163, 0.5258157, 0.5258154, 0.5258152, 0.5258146, 0.525815, 
    0.5258148, 0.5258152, 0.5258154, 0.5258153, 0.525816, 0.5258158, 
    0.5258172, 0.5258166, 0.5258182, 0.5258179, 0.5258183, 0.5258181, 
    0.5258185, 0.5258182, 0.5258188, 0.5258189, 0.5258188, 0.5258192, 
    0.5258181, 0.5258185, 0.5258153, 0.5258154, 0.5258154, 0.5258151, 
    0.525815, 0.5258147, 0.525815, 0.5258151, 0.5258155, 0.5258157, 
    0.5258158, 0.5258163, 0.5258167, 0.5258174, 0.5258179, 0.5258182, 
    0.525818, 0.5258182, 0.525818, 0.5258179, 0.5258189, 0.5258183, 
    0.5258192, 0.5258191, 0.5258188, 0.5258191, 0.5258154, 0.5258152, 
    0.5258149, 0.5258152, 0.5258147, 0.525815, 0.5258151, 0.5258158, 
    0.5258159, 0.5258161, 0.5258163, 0.5258167, 0.5258173, 0.5258178, 
    0.5258183, 0.5258182, 0.5258183, 0.5258183, 0.5258181, 0.5258184, 
    0.5258185, 0.5258183, 0.5258191, 0.5258189, 0.5258191, 0.525819, 
    0.5258153, 0.5258155, 0.5258154, 0.5258155, 0.5258154, 0.525816, 
    0.5258162, 0.525817, 0.5258167, 0.5258172, 0.5258167, 0.5258168, 
    0.5258172, 0.5258167, 0.5258178, 0.5258171, 0.5258184, 0.5258177, 
    0.5258184, 0.5258183, 0.5258185, 0.5258187, 0.5258189, 0.5258194, 
    0.5258193, 0.5258197, 0.5258157, 0.525816, 0.525816, 0.5258162, 
    0.5258164, 0.5258168, 0.5258175, 0.5258172, 0.5258176, 0.5258178, 
    0.525817, 0.5258175, 0.5258161, 0.5258164, 0.5258162, 0.5258158, 
    0.5258173, 0.5258165, 0.5258179, 0.5258175, 0.5258187, 0.5258181, 
    0.5258192, 0.5258198, 0.5258203, 0.5258208, 0.5258161, 0.525816, 
    0.5258163, 0.5258166, 0.525817, 0.5258175, 0.5258176, 0.5258176, 
    0.5258179, 0.5258181, 0.5258177, 0.5258182, 0.5258164, 0.5258173, 
    0.5258159, 0.5258163, 0.5258166, 0.5258165, 0.5258172, 0.5258173, 
    0.525818, 0.5258176, 0.5258197, 0.5258188, 0.5258212, 0.5258206, 
    0.5258159, 0.5258161, 0.5258169, 0.5258165, 0.5258175, 0.5258178, 
    0.525818, 0.5258183, 0.5258183, 0.5258185, 0.5258182, 0.5258184, 
    0.5258175, 0.5258179, 0.5258168, 0.525817, 0.5258169, 0.5258168, 
    0.5258172, 0.5258177, 0.5258177, 0.5258179, 0.5258182, 0.5258175, 
    0.5258198, 0.5258184, 0.5258163, 0.5258167, 0.5258168, 0.5258167, 
    0.5258178, 0.5258174, 0.5258185, 0.5258182, 0.5258186, 0.5258184, 
    0.5258183, 0.525818, 0.5258179, 0.5258174, 0.525817, 0.5258167, 
    0.5258167, 0.5258171, 0.5258177, 0.5258183, 0.5258182, 0.5258186, 
    0.5258175, 0.5258179, 0.5258178, 0.5258182, 0.5258172, 0.525818, 
    0.525817, 0.525817, 0.5258173, 0.525818, 0.5258181, 0.5258182, 0.5258182, 
    0.5258178, 0.5258176, 0.5258173, 0.5258173, 0.525817, 0.5258169, 
    0.525817, 0.5258172, 0.5258178, 0.5258182, 0.5258187, 0.5258188, 
    0.5258194, 0.5258189, 0.5258198, 0.5258191, 0.5258203, 0.5258181, 
    0.5258191, 0.5258174, 0.5258176, 0.5258179, 0.5258186, 0.5258182, 
    0.5258187, 0.5258176, 0.5258171, 0.525817, 0.5258167, 0.525817, 0.525817, 
    0.5258172, 0.5258172, 0.5258178, 0.5258174, 0.5258183, 0.5258187, 
    0.5258197, 0.5258203, 0.5258209, 0.5258211, 0.5258212, 0.5258213 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  7.709882e-21, -1.541976e-20, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, -1.003089e-36, 1.541976e-20, -1.027984e-20, 1.798972e-20, 
    1.541976e-20, 7.709882e-21, 2.569961e-21, -5.139921e-21, -1.003089e-36, 
    2.569961e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 0, 
    7.709882e-21, -1.798972e-20, -2.569961e-21, 2.569961e-21, 7.709882e-21, 
    1.28498e-20, -7.709882e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    -1.003089e-36, 1.003089e-36, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 1.027984e-20, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    1.28498e-20, -5.139921e-21, 5.139921e-21, -1.003089e-36, 7.709882e-21, 
    2.569961e-21, -1.28498e-20, 1.027984e-20, -5.139921e-21, -1.798972e-20, 
    -1.003089e-36, -2.569961e-21, 2.569961e-21, -2.569961e-21, 1.003089e-36, 
    0, -7.709882e-21, -2.569961e-20, 2.312965e-20, 1.28498e-20, 1.541976e-20, 
    1.027984e-20, -1.027984e-20, -2.569961e-21, -7.709882e-21, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, 1.28498e-20, -2.569961e-21, 
    1.027984e-20, 7.709882e-21, -2.569961e-21, 2.569961e-21, 1.28498e-20, 0, 
    -1.28498e-20, 7.709882e-21, 1.541976e-20, 7.709882e-21, 0, 5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, 0, -2.569961e-21, 
    -7.709882e-21, 1.28498e-20, 5.139921e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, -1.541976e-20, 
    -1.541976e-20, -5.139921e-21, 2.569961e-21, -7.709882e-21, 1.541976e-20, 
    0, 1.28498e-20, -1.003089e-36, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -1.28498e-20, 2.569961e-21, -1.28498e-20, -7.709882e-21, 
    1.003089e-36, -5.139921e-21, 0, -7.709882e-21, -1.027984e-20, 
    -1.003089e-36, -2.312965e-20, -1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 1.28498e-20, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    -2.055969e-20, -5.139921e-21, -1.541976e-20, 5.139921e-21, 1.798972e-20, 
    -1.28498e-20, 0, 2.569961e-21, 2.569961e-21, 1.027984e-20, 1.28498e-20, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    1.28498e-20, 1.003089e-36, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, -2.312965e-20, 7.709882e-21, 0, 
    -7.709882e-21, 1.027984e-20, -1.541976e-20, 1.541976e-20, 1.027984e-20, 
    0, 1.28498e-20, 7.709882e-21, 5.139921e-21, -1.28498e-20, -1.027984e-20, 
    -2.569961e-21, -1.027984e-20, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, 1.541976e-20, 1.28498e-20, 5.139921e-21, -2.055969e-20, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, 1.28498e-20, 1.28498e-20, 7.709882e-21, 7.709882e-21, 
    7.709882e-21, -2.569961e-21, -7.709882e-21, 2.569961e-21, -1.541976e-20, 
    2.569961e-21, -5.139921e-21, 2.055969e-20, 5.139921e-21, -5.139921e-21, 
    -2.055969e-20, 1.003089e-36, 1.28498e-20, 1.003089e-36, -2.569961e-21, 
    -1.027984e-20, -1.003089e-36, -5.139921e-21, -7.709882e-21, 
    -2.312965e-20, 5.139921e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, 
    -2.055969e-20, -7.709882e-21, 5.139921e-21, -1.798972e-20, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 2.055969e-20, 5.139921e-21, -7.709882e-21, 
    1.28498e-20, 2.569961e-21, -7.709882e-21, -5.139921e-21, -2.569961e-21, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, 1.027984e-20, -1.28498e-20, 
    -1.28498e-20, -1.798972e-20, -1.027984e-20, 7.709882e-21, 5.139921e-21, 
    1.027984e-20, -1.798972e-20, -1.541976e-20, -1.28498e-20, 5.139921e-21, 
    -1.28498e-20, 1.798972e-20, 7.709882e-21, -7.709882e-21, -1.027984e-20, 
    2.055969e-20, 1.798972e-20, -1.798972e-20, 5.139921e-21, 0, 5.139921e-21, 
    7.709882e-21, -7.709882e-21, 1.003089e-36, 5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 2.569961e-21, 2.569961e-20, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -1.003089e-36, -1.798972e-20, -7.709882e-21, 
    -2.055969e-20, -1.027984e-20, 1.798972e-20, 1.798972e-20, 1.28498e-20, 
    1.28498e-20, -1.541976e-20, -1.541976e-20, -1.027984e-20, -1.541976e-20, 
    -5.139921e-21, -1.027984e-20, -2.569961e-21, -2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, -7.709882e-21, 0, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, 2.569961e-21, 1.027984e-20, -7.709882e-21, -2.569961e-21, 
    -7.709882e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, -7.709882e-21, 
    2.569961e-21, -1.28498e-20, 2.055969e-20, -7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -1.798972e-20, -2.569961e-21, 1.28498e-20, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, 2.569961e-21, 7.709882e-21, 1.798972e-20, 5.139921e-21,
  -1.027984e-20, 7.709882e-21, -2.569961e-21, 1.027984e-20, -1.003089e-36, 
    -5.139921e-21, 2.569961e-21, -1.027984e-20, -1.28498e-20, -5.139921e-21, 
    7.709882e-21, -5.139921e-21, -5.139921e-21, -7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, 7.709882e-21, 5.139921e-21, 
    1.28498e-20, 2.569961e-21, 1.003089e-36, 0, 5.139921e-21, -1.027984e-20, 
    1.027984e-20, 2.569961e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, -7.709882e-21, 
    1.003089e-36, -2.569961e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, 1.027984e-20, 7.709882e-21, 
    1.027984e-20, -5.139921e-21, -7.709882e-21, -2.569961e-21, -1.541976e-20, 
    5.139921e-21, -1.28498e-20, 1.003089e-36, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 7.709882e-21, -2.569961e-21, 
    5.139921e-21, 0, -2.569961e-21, 1.003089e-36, -7.709882e-21, 
    -2.055969e-20, 0, 1.003089e-36, 2.569961e-21, 1.027984e-20, 
    -2.569961e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 0, 2.569961e-21, 1.027984e-20, -7.709882e-21, 
    -7.709882e-21, 5.139921e-21, 1.027984e-20, -7.709882e-21, -1.027984e-20, 
    7.709882e-21, 5.139921e-21, 1.027984e-20, -2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -2.569961e-21, 0, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 7.709882e-21, -1.003089e-36, 7.709882e-21, 0, 
    -1.28498e-20, 2.569961e-21, 1.28498e-20, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, 0, 5.139921e-21, 1.027984e-20, 0, 7.709882e-21, 
    -1.027984e-20, 0, -7.709882e-21, 1.798972e-20, -5.139921e-21, 0, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 5.139921e-21, 0, 
    0, -5.139921e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    5.139921e-21, 1.003089e-36, 5.139921e-21, -7.709882e-21, -2.569961e-21, 
    1.003089e-36, 0, 7.709882e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.28498e-20, -5.139921e-21, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    5.139921e-21, -7.709882e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    1.003089e-36, 1.798972e-20, 2.569961e-21, 1.28498e-20, -1.003089e-36, 
    2.569961e-21, 1.027984e-20, -1.28498e-20, -7.709882e-21, -1.003089e-36, 
    2.569961e-21, 0, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -2.569961e-21, 1.541976e-20, -5.139921e-21, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 0, 7.709882e-21, 7.709882e-21, -2.569961e-21, 0, 
    5.139921e-21, 7.709882e-21, 5.139921e-21, 5.139921e-21, 7.709882e-21, 
    -5.139921e-21, 0, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, 7.709882e-21, 
    -1.027984e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 0, 1.027984e-20, 7.709882e-21, 0, -5.139921e-21, 
    2.569961e-21, 0, -7.709882e-21, -1.027984e-20, -1.798972e-20, 
    7.709882e-21, 7.709882e-21, 0, -5.139921e-21, 0, 1.28498e-20, 
    7.709882e-21, 2.569961e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, 
    2.569961e-21, 1.28498e-20, 1.28498e-20, 2.569961e-21, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, -1.003089e-36, -1.027984e-20, 1.027984e-20, 
    5.139921e-21, 2.569961e-21, -1.003089e-36, 0, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    0, -7.709882e-21, 1.027984e-20, 1.003089e-36, 1.28498e-20, -5.139921e-21, 
    2.569961e-21, -1.027984e-20, -5.139921e-21, -7.709882e-21, 1.003089e-36, 
    -5.139921e-21, -1.28498e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, 0, 2.569961e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -1.798972e-20, -5.139921e-21, -5.139921e-21, -1.798972e-20, 
    -7.709882e-21, -1.027984e-20, 2.569961e-21, 0, 0, 5.139921e-21, 
    -1.28498e-20, -7.709882e-21, -5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, -1.003089e-36, 5.139921e-21, 5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, -2.569961e-21, 0, 0, 0, -2.569961e-21, -7.709882e-21, 
    1.28498e-20, 2.569961e-21, 1.798972e-20, 2.569961e-21, 0, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, -1.28498e-20, 2.569961e-21, -5.139921e-21, 
    -7.709882e-21, 0, 0, -1.027984e-20, 0, 1.027984e-20, 2.569961e-21, 
    5.139921e-21, 0, 1.003089e-36, -1.027984e-20, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 1.28498e-20, 
    -1.798972e-20, -5.139921e-21,
  1.027984e-20, 1.003089e-36, -7.709882e-21, 1.027984e-20, -7.709882e-21, 0, 
    -2.569961e-21, 7.709882e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    2.569961e-21, 1.28498e-20, 1.027984e-20, -7.709882e-21, -5.139921e-21, 
    5.139921e-21, -2.569961e-21, 5.139921e-21, 1.28498e-20, 1.28498e-20, 
    -1.28498e-20, 7.709882e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, 5.139921e-21, 1.28498e-20, 2.055969e-20, 1.28498e-20, 
    7.709882e-21, -2.569961e-21, 2.569961e-21, -1.027984e-20, -2.312965e-20, 
    -1.027984e-20, -5.139921e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, 1.003089e-36, -1.027984e-20, 
    2.569961e-21, -2.569961e-21, 0, -2.569961e-21, 7.709882e-21, 
    -7.709882e-21, 0, 5.139921e-21, 0, 7.709882e-21, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, 
    5.139921e-21, 0, 7.709882e-21, 5.139921e-21, 1.541976e-20, 1.003089e-36, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 1.027984e-20, 7.709882e-21, -1.798972e-20, 
    -2.569961e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, 0, 
    -1.28498e-20, -5.139921e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    1.027984e-20, -2.569961e-21, -5.139921e-21, 0, -7.709882e-21, 0, 
    -5.139921e-21, 2.569961e-21, 1.003089e-36, -2.569961e-21, 1.28498e-20, 
    1.798972e-20, -7.709882e-21, 5.139921e-21, 1.28498e-20, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, -5.139921e-21, 
    1.541976e-20, -7.709882e-21, -7.709882e-21, 2.055969e-20, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -1.027984e-20, -7.709882e-21, 0, 
    7.709882e-21, 5.139921e-21, 1.003089e-36, 0, -1.541976e-20, 1.003089e-36, 
    -1.027984e-20, 5.139921e-21, 7.709882e-21, 5.139921e-21, -7.709882e-21, 
    -2.569961e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -7.709882e-21, 1.798972e-20, 0, 5.139921e-21, 2.569961e-21, 
    -7.709882e-21, -1.541976e-20, -2.569961e-21, -2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, 
    2.569961e-21, -7.709882e-21, -2.569961e-21, 1.027984e-20, -1.003089e-36, 
    0, -7.709882e-21, -2.826957e-20, -1.541976e-20, -1.541976e-20, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 7.709882e-21, 1.003089e-36, 
    1.027984e-20, -1.027984e-20, 1.28498e-20, 7.709882e-21, 2.569961e-21, 0, 
    -2.569961e-21, 0, -1.28498e-20, -5.139921e-21, 7.709882e-21, 
    -5.139921e-21, 7.709882e-21, -7.709882e-21, -7.709882e-21, 7.709882e-21, 
    0, 7.709882e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    -1.798972e-20, -7.709882e-21, 1.28498e-20, 1.541976e-20, 2.569961e-21, 
    1.28498e-20, -5.139921e-21, -2.569961e-21, -1.003089e-36, 1.027984e-20, 
    -1.003089e-36, 0, 1.28498e-20, -7.709882e-21, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    7.709882e-21, 7.709882e-21, -2.569961e-21, -5.139921e-21, 0, 
    -5.139921e-21, 7.709882e-21, 5.139921e-21, -7.709882e-21, 7.709882e-21, 
    2.569961e-21, 2.055969e-20, 0, -5.139921e-21, -5.139921e-21, 
    7.709882e-21, 1.027984e-20, 7.709882e-21, -2.569961e-21, 0, 7.709882e-21, 
    0, 2.569961e-21, 7.709882e-21, 7.709882e-21, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, 1.541976e-20, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, -5.139921e-21, 1.798972e-20, 7.709882e-21, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, -1.541976e-20, 
    1.027984e-20, 1.28498e-20, 1.003089e-36, 7.709882e-21, -7.709882e-21, 
    2.055969e-20, -7.709882e-21, 1.027984e-20, -1.541976e-20, 1.003089e-36, 
    -7.709882e-21, -2.569961e-21, 1.28498e-20, -1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, 0, -5.139921e-21, 
    1.003089e-36, 0, -2.569961e-21, 1.027984e-20, -5.139921e-21, 
    5.139921e-21, 1.003089e-36, -2.055969e-20, 2.569961e-21, -5.139921e-21, 
    0, 1.027984e-20, -2.569961e-21, 1.541976e-20, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, 1.541976e-20, -5.139921e-21, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, -1.541976e-20, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, -1.28498e-20, 
    5.139921e-21, -1.798972e-20, -7.709882e-21, -2.569961e-21, 0, 
    -1.027984e-20, -7.709882e-21, 7.709882e-21, -1.027984e-20, 1.541976e-20, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -1.541976e-20, -1.541976e-20, 5.139921e-21, -7.709882e-21, 
    0, -5.139921e-21, -1.027984e-20, 1.28498e-20, 1.027984e-20, -1.28498e-20, 
    -5.139921e-21, -5.139921e-21, 1.003089e-36, -1.28498e-20, 0, 0, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20,
  -2.569961e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, -1.798972e-20, 
    -5.139921e-21, -1.28498e-20, -1.027984e-20, -1.027984e-20, -1.28498e-20, 
    -1.541976e-20, -7.709882e-21, 1.28498e-20, -5.139921e-21, 5.139921e-21, 
    7.709882e-21, -5.139921e-21, 1.003089e-36, 1.027984e-20, -2.312965e-20, 
    1.541976e-20, -1.541976e-20, 0, -1.28498e-20, -1.003089e-36, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, 1.798972e-20, 1.027984e-20, 
    -2.569961e-21, -1.027984e-20, 1.003089e-36, 1.28498e-20, 5.139921e-21, 
    1.027984e-20, 2.569961e-21, -1.28498e-20, 1.28498e-20, -1.027984e-20, 
    7.709882e-21, 1.027984e-20, -2.569961e-21, 1.027984e-20, -2.055969e-20, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, 0, -5.139921e-21, 
    1.541976e-20, -1.541976e-20, 1.28498e-20, 1.003089e-36, 5.139921e-21, 
    1.027984e-20, 0, 2.569961e-21, -1.003089e-36, 1.541976e-20, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, -7.709882e-21, 1.28498e-20, -2.569961e-21, 
    1.003089e-36, -1.28498e-20, -7.709882e-21, -2.569961e-21, 1.003089e-36, 
    -5.139921e-21, 7.709882e-21, 1.027984e-20, -7.709882e-21, -5.139921e-21, 
    -2.569961e-21, 1.28498e-20, 1.027984e-20, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, 1.027984e-20, 7.709882e-21, -2.569961e-21, -1.28498e-20, 
    -5.139921e-21, 2.055969e-20, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    -5.139921e-21, 7.709882e-21, 2.569961e-21, -7.709882e-21, 5.139921e-21, 
    7.709882e-21, -7.709882e-21, 2.569961e-21, 1.027984e-20, 1.798972e-20, 
    -1.798972e-20, 7.709882e-21, -1.541976e-20, 1.28498e-20, -2.569961e-20, 
    -1.003089e-36, 1.28498e-20, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 2.569961e-21, -1.798972e-20, 1.28498e-20, -2.569961e-21, 
    1.027984e-20, 1.541976e-20, -1.28498e-20, 7.709882e-21, 2.569961e-21, 
    5.139921e-21, 1.28498e-20, -1.027984e-20, -2.569961e-21, 1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 5.139921e-21, 0, 2.569961e-21, 1.027984e-20, 
    -5.139921e-21, -7.709882e-21, -1.027984e-20, 5.139921e-21, -2.312965e-20, 
    -2.569961e-21, 5.139921e-21, -1.28498e-20, 5.139921e-21, 1.28498e-20, 
    1.027984e-20, -2.569961e-21, 0, -5.139921e-21, -7.709882e-21, 
    -2.569961e-21, 1.027984e-20, 1.027984e-20, -1.798972e-20, 0, 
    -1.003089e-36, 0, -1.027984e-20, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -2.569961e-20, -5.139921e-21, -1.541976e-20, 
    -2.569961e-21, -1.541976e-20, 0, 7.709882e-21, 2.055969e-20, 
    2.569961e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    -1.003089e-36, -1.027984e-20, -7.709882e-21, 2.569961e-21, 1.541976e-20, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, 1.027984e-20, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, 1.798972e-20, 2.569961e-21, -1.28498e-20, 
    -2.569961e-21, -7.709882e-21, -1.28498e-20, 1.28498e-20, -2.569961e-21, 
    0, 2.569961e-21, -1.798972e-20, -1.003089e-36, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, -5.139921e-21, 0, 1.541976e-20, 
    -1.798972e-20, 2.569961e-21, 1.541976e-20, -5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 7.709882e-21, -7.709882e-21, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, 7.709882e-21, -2.569961e-21, 5.139921e-21, 1.003089e-36, 
    -7.709882e-21, 2.569961e-21, -2.312965e-20, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, 1.003089e-36, -1.28498e-20, -7.709882e-21, -1.28498e-20, 
    -7.709882e-21, 7.709882e-21, 1.28498e-20, 1.003089e-36, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, -1.28498e-20, -1.28498e-20, -1.541976e-20, 
    -2.569961e-21, 7.709882e-21, -1.28498e-20, 1.798972e-20, 2.569961e-21, 
    -1.003089e-36, 5.139921e-21, 1.003089e-36, 5.139921e-21, 1.28498e-20, 
    5.139921e-21, -1.798972e-20, -5.139921e-21, -1.003089e-36, 2.569961e-21, 
    -2.312965e-20, -2.569961e-21, -1.003089e-36, 7.709882e-21, 1.28498e-20, 
    -5.139921e-21, 5.139921e-21, -7.709882e-21, 7.709882e-21, 0, 
    5.139921e-21, -7.709882e-21, -7.709882e-21, -2.569961e-21, -1.027984e-20, 
    -7.709882e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, -7.709882e-21, 
    -7.709882e-21, 2.569961e-21, 2.569961e-21, 1.027984e-20, 2.569961e-21, 
    2.569961e-21, 7.709882e-21, 1.28498e-20, 0, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, -1.28498e-20, 
    -5.139921e-21, 5.139921e-21, -1.798972e-20, 7.709882e-21, -1.798972e-20, 
    0, 2.569961e-21, -1.28498e-20, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, -7.709882e-21, 7.709882e-21, 1.28498e-20, -1.027984e-20, 
    5.139921e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -1.28498e-20, 5.139921e-21, -7.709882e-21, 1.541976e-20, 2.569961e-21, 
    -1.027984e-20, 1.798972e-20, -2.569961e-20, 2.569961e-20, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -5.139921e-21, 5.139921e-21, -2.055969e-20, 
    1.003089e-36, 0, -1.003089e-36, 7.709882e-21, -7.709882e-21, 
    7.709882e-21, -1.027984e-20,
  5.139921e-21, -1.027984e-20, 0, -2.569961e-21, 2.569961e-21, 1.541976e-20, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, -2.055969e-20, 
    -7.709882e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, 2.312965e-20, 
    -5.139921e-21, -1.541976e-20, 1.28498e-20, 1.28498e-20, 2.055969e-20, 
    -2.569961e-21, -2.569961e-21, -3.009266e-36, -2.569961e-21, -1.28498e-20, 
    5.139921e-21, 2.312965e-20, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -1.28498e-20, -7.709882e-21, 1.541976e-20, 1.027984e-20, 1.798972e-20, 
    1.003089e-36, -2.569961e-21, 2.569961e-21, 1.003089e-36, 0, 
    -5.139921e-21, -2.312965e-20, -5.139921e-21, -7.709882e-21, 
    -1.798972e-20, -5.139921e-21, 5.139921e-21, -2.055969e-20, 2.569961e-21, 
    -1.28498e-20, 1.003089e-36, 5.139921e-21, 2.055969e-20, -1.541976e-20, 
    2.569961e-21, -2.312965e-20, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 1.027984e-20, -1.28498e-20, 5.139921e-21, 1.003089e-36, 
    1.541976e-20, -2.569961e-21, -1.027984e-20, 7.709882e-21, -1.027984e-20, 
    -7.709882e-21, 2.569961e-21, -2.569961e-20, -2.569961e-21, -2.312965e-20, 
    0, -5.139921e-21, 5.139921e-21, 7.709882e-21, -2.826957e-20, 
    1.027984e-20, -7.709882e-21, 1.027984e-20, 1.027984e-20, 2.569961e-20, 
    -3.083953e-20, 2.569961e-21, -1.027984e-20, -1.027984e-20, 5.139921e-21, 
    1.541976e-20, 1.28498e-20, -7.709882e-21, -1.027984e-20, -1.28498e-20, 
    -2.569961e-21, 1.541976e-20, 5.139921e-21, -1.541976e-20, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -1.003089e-36, 5.139921e-21, 0, 
    5.139921e-21, 1.027984e-20, 1.28498e-20, 7.709882e-21, -1.541976e-20, 
    -2.826957e-20, 1.541976e-20, -1.541976e-20, -5.139921e-21, -5.139921e-21, 
    -1.798972e-20, -1.003089e-36, 1.28498e-20, 7.709882e-21, -1.798972e-20, 
    7.709882e-21, -2.055969e-20, -1.003089e-36, 5.139921e-21, -1.027984e-20, 
    5.139921e-21, 0, -2.569961e-21, 2.569961e-21, -7.709882e-21, 
    -7.709882e-21, -3.083953e-20, -2.569961e-21, -5.139921e-21, -1.28498e-20, 
    2.055969e-20, 2.569961e-21, -7.709882e-21, 1.541976e-20, -2.569961e-21, 
    1.28498e-20, 1.28498e-20, 5.015443e-37, 7.709882e-21, -7.709882e-21, 
    -1.003089e-36, -2.826957e-20, 1.28498e-20, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, 3.083953e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -1.28498e-20, 1.28498e-20, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 1.027984e-20, 5.139921e-21, 0, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, 1.027984e-20, 2.826957e-20, -5.139921e-21, 
    -1.541976e-20, 1.541976e-20, 2.569961e-21, -7.709882e-21, 5.139921e-21, 
    2.312965e-20, -1.28498e-20, 2.569961e-21, 1.003089e-36, -1.28498e-20, 
    5.139921e-21, 7.709882e-21, 1.541976e-20, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, 1.027984e-20, 
    3.083953e-20, 0, 1.027984e-20, -7.709882e-21, -5.139921e-21, 
    2.569961e-20, 2.569961e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, -1.28498e-20, 7.709882e-21, -1.003089e-36, 7.709882e-21, 
    2.569961e-21, -5.139921e-21, 0, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -2.569961e-21, -3.340949e-20, 5.139921e-21, 7.709882e-21, 1.541976e-20, 
    7.709882e-21, 1.541976e-20, -3.009266e-36, 1.28498e-20, 5.139921e-21, 
    1.541976e-20, 2.569961e-21, -7.709882e-21, 7.709882e-21, 1.541976e-20, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, -1.28498e-20, 
    -2.569961e-21, 7.709882e-21, 1.28498e-20, 7.709882e-21, -1.28498e-20, 
    7.709882e-21, 1.027984e-20, 5.139921e-21, -2.569961e-21, -1.798972e-20, 
    -2.569961e-21, -5.139921e-21, -1.28498e-20, -7.709882e-21, -1.027984e-20, 
    -5.139921e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, 
    -7.709882e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, 2.055969e-20, 
    1.798972e-20, -7.709882e-21, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    7.709882e-21, 1.027984e-20, -1.003089e-36, 2.569961e-21, 1.541976e-20, 
    7.709882e-21, -1.798972e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -1.798972e-20, -2.312965e-20, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -1.003089e-36, 1.027984e-20, 1.027984e-20, 
    1.541976e-20, -1.003089e-36, -1.28498e-20, 2.569961e-21, 7.709882e-21, 
    -1.541976e-20, -1.28498e-20, -1.28498e-20, -1.027984e-20, -7.709882e-21, 
    7.709882e-21, -5.139921e-21, -2.055969e-20, 5.139921e-21, 1.003089e-36, 
    1.28498e-20, -2.569961e-21, 1.541976e-20, -2.826957e-20, -2.569961e-21, 
    7.709882e-21, 1.28498e-20, -7.709882e-21, 5.139921e-21, 1.003089e-36, 
    2.055969e-20, 2.569961e-21, -2.569961e-21, 5.139921e-21, 2.569961e-20, 
    7.709882e-21, 7.709882e-21, -1.28498e-20, 2.569961e-21, -1.003089e-36, 
    -1.027984e-20, -2.312965e-20, 1.027984e-20, -2.569961e-21, 1.027984e-20, 
    1.027984e-20, 1.28498e-20, -1.798972e-20, -1.28498e-20, -2.569961e-21, 
    5.139921e-21, 5.139921e-21, 7.709882e-21, 1.798972e-20, 7.709882e-21, 
    2.826957e-20, -2.569961e-21, -1.027984e-20, -1.027984e-20, -1.003089e-36, 
    -1.28498e-20, 7.709882e-21,
  6.259379e-29, 6.259386e-29, 6.259385e-29, 6.25939e-29, 6.259387e-29, 
    6.25939e-29, 6.259381e-29, 6.259386e-29, 6.259383e-29, 6.25938e-29, 
    6.259399e-29, 6.25939e-29, 6.25941e-29, 6.259404e-29, 6.259419e-29, 
    6.259408e-29, 6.25942e-29, 6.259418e-29, 6.259425e-29, 6.259423e-29, 
    6.259432e-29, 6.259426e-29, 6.259437e-29, 6.259431e-29, 6.259432e-29, 
    6.259426e-29, 6.259392e-29, 6.259398e-29, 6.259391e-29, 6.259392e-29, 
    6.259392e-29, 6.259387e-29, 6.259384e-29, 6.259379e-29, 6.25938e-29, 
    6.259384e-29, 6.259393e-29, 6.25939e-29, 6.259398e-29, 6.259397e-29, 
    6.259405e-29, 6.259402e-29, 6.259416e-29, 6.259412e-29, 6.259423e-29, 
    6.25942e-29, 6.259423e-29, 6.259422e-29, 6.259423e-29, 6.259419e-29, 
    6.259421e-29, 6.259417e-29, 6.259402e-29, 6.259407e-29, 6.259394e-29, 
    6.259386e-29, 6.259381e-29, 6.259378e-29, 6.259378e-29, 6.259379e-29, 
    6.259384e-29, 6.259388e-29, 6.259392e-29, 6.259394e-29, 6.259397e-29, 
    6.259404e-29, 6.259408e-29, 6.259417e-29, 6.259415e-29, 6.259417e-29, 
    6.25942e-29, 6.259425e-29, 6.259423e-29, 6.259425e-29, 6.259417e-29, 
    6.259423e-29, 6.259414e-29, 6.259417e-29, 6.259398e-29, 6.259391e-29, 
    6.259387e-29, 6.259385e-29, 6.259378e-29, 6.259383e-29, 6.259381e-29, 
    6.259385e-29, 6.259388e-29, 6.259387e-29, 6.259394e-29, 6.259391e-29, 
    6.259408e-29, 6.259401e-29, 6.25942e-29, 6.259416e-29, 6.259421e-29, 
    6.259418e-29, 6.259423e-29, 6.259419e-29, 6.259426e-29, 6.259428e-29, 
    6.259426e-29, 6.259431e-29, 6.259419e-29, 6.259423e-29, 6.259387e-29, 
    6.259387e-29, 6.259388e-29, 6.259384e-29, 6.259383e-29, 6.259379e-29, 
    6.259382e-29, 6.259384e-29, 6.259388e-29, 6.25939e-29, 6.259393e-29, 
    6.259398e-29, 6.259403e-29, 6.25941e-29, 6.259416e-29, 6.259419e-29, 
    6.259417e-29, 6.259419e-29, 6.259417e-29, 6.259416e-29, 6.259427e-29, 
    6.259421e-29, 6.259431e-29, 6.25943e-29, 6.259426e-29, 6.25943e-29, 
    6.259387e-29, 6.259385e-29, 6.259381e-29, 6.259385e-29, 6.259379e-29, 
    6.259382e-29, 6.259384e-29, 6.259391e-29, 6.259393e-29, 6.259395e-29, 
    6.259398e-29, 6.259402e-29, 6.259409e-29, 6.259415e-29, 6.25942e-29, 
    6.25942e-29, 6.25942e-29, 6.259421e-29, 6.259418e-29, 6.259422e-29, 
    6.259422e-29, 6.259421e-29, 6.25943e-29, 6.259427e-29, 6.25943e-29, 
    6.259428e-29, 6.259386e-29, 6.259388e-29, 6.259387e-29, 6.259389e-29, 
    6.259388e-29, 6.259394e-29, 6.259396e-29, 6.259406e-29, 6.259402e-29, 
    6.259408e-29, 6.259402e-29, 6.259404e-29, 6.259408e-29, 6.259403e-29, 
    6.259414e-29, 6.259407e-29, 6.259421e-29, 6.259413e-29, 6.259422e-29, 
    6.25942e-29, 6.259423e-29, 6.259425e-29, 6.259428e-29, 6.259433e-29, 
    6.259432e-29, 6.259437e-29, 6.259391e-29, 6.259394e-29, 6.259394e-29, 
    6.259397e-29, 6.259399e-29, 6.259404e-29, 6.259411e-29, 6.259408e-29, 
    6.259413e-29, 6.259414e-29, 6.259406e-29, 6.259411e-29, 6.259396e-29, 
    6.259398e-29, 6.259397e-29, 6.259391e-29, 6.259408e-29, 6.2594e-29, 
    6.259416e-29, 6.259411e-29, 6.259425e-29, 6.259418e-29, 6.259431e-29, 
    6.259437e-29, 6.259443e-29, 6.259449e-29, 6.259396e-29, 6.259394e-29, 
    6.259397e-29, 6.259402e-29, 6.259406e-29, 6.259411e-29, 6.259412e-29, 
    6.259413e-29, 6.259416e-29, 6.259418e-29, 6.259413e-29, 6.259419e-29, 
    6.259399e-29, 6.259409e-29, 6.259393e-29, 6.259398e-29, 6.259401e-29, 
    6.2594e-29, 6.259408e-29, 6.25941e-29, 6.259417e-29, 6.259413e-29, 
    6.259435e-29, 6.259426e-29, 6.259453e-29, 6.259446e-29, 6.259393e-29, 
    6.259396e-29, 6.259404e-29, 6.2594e-29, 6.259412e-29, 6.259414e-29, 
    6.259417e-29, 6.25942e-29, 6.25942e-29, 6.259422e-29, 6.259419e-29, 
    6.259422e-29, 6.259411e-29, 6.259416e-29, 6.259403e-29, 6.259407e-29, 
    6.259405e-29, 6.259403e-29, 6.259408e-29, 6.259413e-29, 6.259414e-29, 
    6.259415e-29, 6.25942e-29, 6.259412e-29, 6.259437e-29, 6.259422e-29, 
    6.259398e-29, 6.259403e-29, 6.259404e-29, 6.259402e-29, 6.259414e-29, 
    6.25941e-29, 6.259422e-29, 6.259419e-29, 6.259424e-29, 6.259422e-29, 
    6.259421e-29, 6.259417e-29, 6.259416e-29, 6.25941e-29, 6.259405e-29, 
    6.259402e-29, 6.259403e-29, 6.259407e-29, 6.259414e-29, 6.25942e-29, 
    6.259419e-29, 6.259423e-29, 6.259411e-29, 6.259416e-29, 6.259414e-29, 
    6.25942e-29, 6.259408e-29, 6.259418e-29, 6.259405e-29, 6.259406e-29, 
    6.25941e-29, 6.259417e-29, 6.259418e-29, 6.25942e-29, 6.259419e-29, 
    6.259414e-29, 6.259413e-29, 6.25941e-29, 6.259408e-29, 6.259406e-29, 
    6.259404e-29, 6.259406e-29, 6.259408e-29, 6.259414e-29, 6.259419e-29, 
    6.259425e-29, 6.259426e-29, 6.259434e-29, 6.259428e-29, 6.259437e-29, 
    6.259429e-29, 6.259443e-29, 6.259419e-29, 6.259429e-29, 6.25941e-29, 
    6.259412e-29, 6.259416e-29, 6.259424e-29, 6.25942e-29, 6.259425e-29, 
    6.259413e-29, 6.259407e-29, 6.259405e-29, 6.259402e-29, 6.259405e-29, 
    6.259405e-29, 6.259408e-29, 6.259407e-29, 6.259414e-29, 6.25941e-29, 
    6.259421e-29, 6.259425e-29, 6.259436e-29, 6.259443e-29, 6.25945e-29, 
    6.259453e-29, 6.259453e-29, 6.259454e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.145192e-10, 2.154657e-10, 2.152817e-10, 2.160452e-10, 2.156217e-10, 
    2.161216e-10, 2.147111e-10, 2.155033e-10, 2.149976e-10, 2.146044e-10, 
    2.175269e-10, 2.160793e-10, 2.190309e-10, 2.181075e-10, 2.204272e-10, 
    2.188872e-10, 2.207377e-10, 2.203828e-10, 2.214512e-10, 2.211451e-10, 
    2.225117e-10, 2.215925e-10, 2.232201e-10, 2.222922e-10, 2.224373e-10, 
    2.215621e-10, 2.163706e-10, 2.173466e-10, 2.163128e-10, 2.16452e-10, 
    2.163895e-10, 2.156304e-10, 2.152479e-10, 2.144469e-10, 2.145923e-10, 
    2.151806e-10, 2.165146e-10, 2.160618e-10, 2.17203e-10, 2.171772e-10, 
    2.184478e-10, 2.178749e-10, 2.200107e-10, 2.194037e-10, 2.211579e-10, 
    2.207167e-10, 2.211372e-10, 2.210097e-10, 2.211388e-10, 2.204918e-10, 
    2.20769e-10, 2.201997e-10, 2.179822e-10, 2.186339e-10, 2.166904e-10, 
    2.155218e-10, 2.147458e-10, 2.141952e-10, 2.14273e-10, 2.144214e-10, 
    2.151841e-10, 2.159012e-10, 2.164477e-10, 2.168133e-10, 2.171735e-10, 
    2.182638e-10, 2.18841e-10, 2.201334e-10, 2.199002e-10, 2.202953e-10, 
    2.206728e-10, 2.213066e-10, 2.212023e-10, 2.214815e-10, 2.202849e-10, 
    2.210801e-10, 2.197674e-10, 2.201264e-10, 2.172713e-10, 2.161839e-10, 
    2.157216e-10, 2.153171e-10, 2.143329e-10, 2.150125e-10, 2.147446e-10, 
    2.153821e-10, 2.157872e-10, 2.155868e-10, 2.168233e-10, 2.163426e-10, 
    2.188752e-10, 2.177843e-10, 2.206288e-10, 2.199481e-10, 2.207919e-10, 
    2.203613e-10, 2.210992e-10, 2.204351e-10, 2.215854e-10, 2.21836e-10, 
    2.216647e-10, 2.223223e-10, 2.203983e-10, 2.211372e-10, 2.155812e-10, 
    2.156139e-10, 2.157661e-10, 2.15097e-10, 2.15056e-10, 2.144429e-10, 
    2.149885e-10, 2.152208e-10, 2.158106e-10, 2.161595e-10, 2.164912e-10, 
    2.172204e-10, 2.180349e-10, 2.191738e-10, 2.199922e-10, 2.205408e-10, 
    2.202044e-10, 2.205014e-10, 2.201694e-10, 2.200138e-10, 2.217421e-10, 
    2.207716e-10, 2.222278e-10, 2.221472e-10, 2.214881e-10, 2.221563e-10, 
    2.156368e-10, 2.154488e-10, 2.14796e-10, 2.153069e-10, 2.143761e-10, 
    2.148971e-10, 2.151966e-10, 2.163526e-10, 2.166066e-10, 2.168421e-10, 
    2.173073e-10, 2.179043e-10, 2.189515e-10, 2.198628e-10, 2.206948e-10, 
    2.206338e-10, 2.206553e-10, 2.208411e-10, 2.203808e-10, 2.209167e-10, 
    2.210066e-10, 2.207715e-10, 2.221364e-10, 2.217465e-10, 2.221455e-10, 
    2.218916e-10, 2.155099e-10, 2.158263e-10, 2.156553e-10, 2.159768e-10, 
    2.157503e-10, 2.167574e-10, 2.170594e-10, 2.184724e-10, 2.178925e-10, 
    2.188154e-10, 2.179863e-10, 2.181332e-10, 2.188455e-10, 2.180311e-10, 
    2.198125e-10, 2.186047e-10, 2.208483e-10, 2.196421e-10, 2.209239e-10, 
    2.206912e-10, 2.210766e-10, 2.214217e-10, 2.218561e-10, 2.226573e-10, 
    2.224717e-10, 2.231419e-10, 2.16298e-10, 2.167083e-10, 2.166722e-10, 
    2.171017e-10, 2.174193e-10, 2.181078e-10, 2.19212e-10, 2.187968e-10, 
    2.195591e-10, 2.197122e-10, 2.18554e-10, 2.192651e-10, 2.16983e-10, 
    2.173516e-10, 2.171322e-10, 2.163303e-10, 2.188924e-10, 2.175775e-10, 
    2.200057e-10, 2.192933e-10, 2.213725e-10, 2.203384e-10, 2.223696e-10, 
    2.232379e-10, 2.240552e-10, 2.250102e-10, 2.169323e-10, 2.166535e-10, 
    2.171528e-10, 2.178435e-10, 2.184846e-10, 2.193368e-10, 2.19424e-10, 
    2.195836e-10, 2.199972e-10, 2.203449e-10, 2.196341e-10, 2.204321e-10, 
    2.174371e-10, 2.190066e-10, 2.16548e-10, 2.172883e-10, 2.178028e-10, 
    2.175771e-10, 2.187493e-10, 2.190256e-10, 2.201483e-10, 2.195679e-10, 
    2.230235e-10, 2.214946e-10, 2.257376e-10, 2.245517e-10, 2.165561e-10, 
    2.169314e-10, 2.182376e-10, 2.176161e-10, 2.193937e-10, 2.198312e-10, 
    2.20187e-10, 2.206417e-10, 2.206908e-10, 2.209602e-10, 2.205187e-10, 
    2.209428e-10, 2.193386e-10, 2.200555e-10, 2.180883e-10, 2.185671e-10, 
    2.183469e-10, 2.181053e-10, 2.188509e-10, 2.196453e-10, 2.196623e-10, 
    2.19917e-10, 2.206347e-10, 2.194009e-10, 2.232208e-10, 2.208615e-10, 
    2.173406e-10, 2.180635e-10, 2.181668e-10, 2.178868e-10, 2.197874e-10, 
    2.190987e-10, 2.209537e-10, 2.204523e-10, 2.212738e-10, 2.208656e-10, 
    2.208055e-10, 2.202813e-10, 2.199549e-10, 2.191303e-10, 2.184594e-10, 
    2.179274e-10, 2.180511e-10, 2.186355e-10, 2.196939e-10, 2.206952e-10, 
    2.204759e-10, 2.212113e-10, 2.192648e-10, 2.20081e-10, 2.197655e-10, 
    2.205881e-10, 2.187857e-10, 2.203204e-10, 2.183935e-10, 2.185624e-10, 
    2.19085e-10, 2.201363e-10, 2.20369e-10, 2.206173e-10, 2.204641e-10, 
    2.197208e-10, 2.19599e-10, 2.190723e-10, 2.189269e-10, 2.185256e-10, 
    2.181934e-10, 2.184969e-10, 2.188157e-10, 2.197211e-10, 2.20537e-10, 
    2.214266e-10, 2.216444e-10, 2.226838e-10, 2.218376e-10, 2.232339e-10, 
    2.220467e-10, 2.241019e-10, 2.204094e-10, 2.220119e-10, 2.191088e-10, 
    2.194216e-10, 2.199872e-10, 2.212846e-10, 2.205842e-10, 2.214034e-10, 
    2.195942e-10, 2.186556e-10, 2.184128e-10, 2.179598e-10, 2.184232e-10, 
    2.183855e-10, 2.188289e-10, 2.186864e-10, 2.197511e-10, 2.191792e-10, 
    2.20804e-10, 2.213969e-10, 2.230716e-10, 2.240982e-10, 2.251434e-10, 
    2.256048e-10, 2.257453e-10, 2.25804e-10 ;

 SOIL2N_TO_SOIL3N =
  1.53228e-11, 1.539041e-11, 1.537727e-11, 1.54318e-11, 1.540155e-11, 
    1.543726e-11, 1.533651e-11, 1.539309e-11, 1.535697e-11, 1.532889e-11, 
    1.553763e-11, 1.543423e-11, 1.564506e-11, 1.557911e-11, 1.57448e-11, 
    1.56348e-11, 1.576698e-11, 1.574163e-11, 1.581794e-11, 1.579608e-11, 
    1.589369e-11, 1.582803e-11, 1.59443e-11, 1.587801e-11, 1.588838e-11, 
    1.582587e-11, 1.545505e-11, 1.552476e-11, 1.545091e-11, 1.546085e-11, 
    1.545639e-11, 1.540217e-11, 1.537485e-11, 1.531763e-11, 1.532802e-11, 
    1.537005e-11, 1.546533e-11, 1.543298e-11, 1.55145e-11, 1.551266e-11, 
    1.560342e-11, 1.55625e-11, 1.571505e-11, 1.567169e-11, 1.579699e-11, 
    1.576548e-11, 1.579551e-11, 1.578641e-11, 1.579563e-11, 1.574941e-11, 
    1.576921e-11, 1.572855e-11, 1.557016e-11, 1.56167e-11, 1.547788e-11, 
    1.539442e-11, 1.533899e-11, 1.529965e-11, 1.530522e-11, 1.531581e-11, 
    1.537029e-11, 1.542152e-11, 1.546055e-11, 1.548667e-11, 1.55124e-11, 
    1.559027e-11, 1.56315e-11, 1.572381e-11, 1.570716e-11, 1.573538e-11, 
    1.576234e-11, 1.580761e-11, 1.580016e-11, 1.582011e-11, 1.573464e-11, 
    1.579144e-11, 1.569767e-11, 1.572332e-11, 1.551938e-11, 1.544171e-11, 
    1.540869e-11, 1.537979e-11, 1.530949e-11, 1.535804e-11, 1.53389e-11, 
    1.538444e-11, 1.541337e-11, 1.539906e-11, 1.548738e-11, 1.545304e-11, 
    1.563395e-11, 1.555602e-11, 1.57592e-11, 1.571058e-11, 1.577085e-11, 
    1.57401e-11, 1.57928e-11, 1.574537e-11, 1.582753e-11, 1.584543e-11, 
    1.583319e-11, 1.588017e-11, 1.574274e-11, 1.579551e-11, 1.539866e-11, 
    1.540099e-11, 1.541186e-11, 1.536407e-11, 1.536114e-11, 1.531735e-11, 
    1.535632e-11, 1.537291e-11, 1.541505e-11, 1.543997e-11, 1.546366e-11, 
    1.551574e-11, 1.557392e-11, 1.565528e-11, 1.571373e-11, 1.575291e-11, 
    1.572889e-11, 1.57501e-11, 1.572639e-11, 1.571527e-11, 1.583872e-11, 
    1.57694e-11, 1.587341e-11, 1.586766e-11, 1.582058e-11, 1.58683e-11, 
    1.540263e-11, 1.53892e-11, 1.534257e-11, 1.537906e-11, 1.531258e-11, 
    1.534979e-11, 1.537119e-11, 1.545376e-11, 1.54719e-11, 1.548872e-11, 
    1.552195e-11, 1.556459e-11, 1.56394e-11, 1.570449e-11, 1.576391e-11, 
    1.575956e-11, 1.576109e-11, 1.577437e-11, 1.574148e-11, 1.577976e-11, 
    1.578619e-11, 1.576939e-11, 1.586689e-11, 1.583903e-11, 1.586753e-11, 
    1.58494e-11, 1.539357e-11, 1.541616e-11, 1.540395e-11, 1.542691e-11, 
    1.541074e-11, 1.548267e-11, 1.550424e-11, 1.560517e-11, 1.556375e-11, 
    1.562967e-11, 1.557045e-11, 1.558094e-11, 1.563182e-11, 1.557365e-11, 
    1.57009e-11, 1.561462e-11, 1.577488e-11, 1.568872e-11, 1.578028e-11, 
    1.576366e-11, 1.579118e-11, 1.581584e-11, 1.584686e-11, 1.590409e-11, 
    1.589084e-11, 1.59387e-11, 1.544985e-11, 1.547916e-11, 1.547659e-11, 
    1.550726e-11, 1.552995e-11, 1.557913e-11, 1.5658e-11, 1.562834e-11, 
    1.56828e-11, 1.569373e-11, 1.5611e-11, 1.566179e-11, 1.549878e-11, 
    1.552512e-11, 1.550944e-11, 1.545217e-11, 1.563517e-11, 1.554125e-11, 
    1.571469e-11, 1.566381e-11, 1.581232e-11, 1.573846e-11, 1.588354e-11, 
    1.594556e-11, 1.600394e-11, 1.607216e-11, 1.549517e-11, 1.547525e-11, 
    1.551091e-11, 1.556025e-11, 1.560604e-11, 1.566691e-11, 1.567314e-11, 
    1.568455e-11, 1.571409e-11, 1.573892e-11, 1.568815e-11, 1.574515e-11, 
    1.553122e-11, 1.564333e-11, 1.546772e-11, 1.552059e-11, 1.555735e-11, 
    1.554122e-11, 1.562495e-11, 1.564469e-11, 1.572488e-11, 1.568343e-11, 
    1.593025e-11, 1.582104e-11, 1.612411e-11, 1.603941e-11, 1.546829e-11, 
    1.54951e-11, 1.55884e-11, 1.554401e-11, 1.567098e-11, 1.570223e-11, 
    1.572764e-11, 1.576012e-11, 1.576363e-11, 1.578287e-11, 1.575134e-11, 
    1.578163e-11, 1.566704e-11, 1.571825e-11, 1.557774e-11, 1.561194e-11, 
    1.55962e-11, 1.557895e-11, 1.563221e-11, 1.568895e-11, 1.569016e-11, 
    1.570836e-11, 1.575962e-11, 1.567149e-11, 1.594434e-11, 1.577582e-11, 
    1.552433e-11, 1.557597e-11, 1.558335e-11, 1.556334e-11, 1.56991e-11, 
    1.564991e-11, 1.57824e-11, 1.57466e-11, 1.580527e-11, 1.577611e-11, 
    1.577182e-11, 1.573438e-11, 1.571106e-11, 1.565216e-11, 1.560424e-11, 
    1.556624e-11, 1.557508e-11, 1.561682e-11, 1.569242e-11, 1.576394e-11, 
    1.574828e-11, 1.580081e-11, 1.566177e-11, 1.572007e-11, 1.569754e-11, 
    1.575629e-11, 1.562755e-11, 1.573717e-11, 1.559953e-11, 1.56116e-11, 
    1.564893e-11, 1.572402e-11, 1.574064e-11, 1.575838e-11, 1.574743e-11, 
    1.569434e-11, 1.568564e-11, 1.564802e-11, 1.563764e-11, 1.560897e-11, 
    1.558524e-11, 1.560692e-11, 1.562969e-11, 1.569436e-11, 1.575264e-11, 
    1.581619e-11, 1.583174e-11, 1.590598e-11, 1.584555e-11, 1.594528e-11, 
    1.586048e-11, 1.600728e-11, 1.574353e-11, 1.585799e-11, 1.565063e-11, 
    1.567297e-11, 1.571337e-11, 1.580605e-11, 1.575602e-11, 1.581453e-11, 
    1.56853e-11, 1.561826e-11, 1.560092e-11, 1.556856e-11, 1.560166e-11, 
    1.559896e-11, 1.563064e-11, 1.562046e-11, 1.569651e-11, 1.565566e-11, 
    1.577171e-11, 1.581407e-11, 1.593369e-11, 1.600702e-11, 1.608167e-11, 
    1.611463e-11, 1.612466e-11, 1.612886e-11 ;

 SOIL2N_vr =
  1.818724, 1.818725, 1.818725, 1.818726, 1.818726, 1.818726, 1.818724, 
    1.818725, 1.818725, 1.818724, 1.818729, 1.818726, 1.818731, 1.818729, 
    1.818733, 1.818731, 1.818733, 1.818733, 1.818735, 1.818734, 1.818736, 
    1.818735, 1.818737, 1.818736, 1.818736, 1.818735, 1.818727, 1.818728, 
    1.818727, 1.818727, 1.818727, 1.818726, 1.818725, 1.818724, 1.818724, 
    1.818725, 1.818727, 1.818726, 1.818728, 1.818728, 1.81873, 1.818729, 
    1.818732, 1.818731, 1.818734, 1.818733, 1.818734, 1.818734, 1.818734, 
    1.818733, 1.818734, 1.818733, 1.818729, 1.81873, 1.818727, 1.818725, 
    1.818724, 1.818723, 1.818723, 1.818724, 1.818725, 1.818726, 1.818727, 
    1.818727, 1.818728, 1.81873, 1.818731, 1.818733, 1.818732, 1.818733, 
    1.818733, 1.818734, 1.818734, 1.818735, 1.818733, 1.818734, 1.818732, 
    1.818733, 1.818728, 1.818726, 1.818726, 1.818725, 1.818724, 1.818725, 
    1.818724, 1.818725, 1.818726, 1.818725, 1.818727, 1.818727, 1.818731, 
    1.818729, 1.818733, 1.818732, 1.818734, 1.818733, 1.818734, 1.818733, 
    1.818735, 1.818735, 1.818735, 1.818736, 1.818733, 1.818734, 1.818725, 
    1.818725, 1.818726, 1.818725, 1.818725, 1.818724, 1.818725, 1.818725, 
    1.818726, 1.818726, 1.818727, 1.818728, 1.818729, 1.818731, 1.818732, 
    1.818733, 1.818733, 1.818733, 1.818733, 1.818732, 1.818735, 1.818734, 
    1.818736, 1.818736, 1.818735, 1.818736, 1.818726, 1.818725, 1.818724, 
    1.818725, 1.818724, 1.818724, 1.818725, 1.818727, 1.818727, 1.818727, 
    1.818728, 1.818729, 1.818731, 1.818732, 1.818733, 1.818733, 1.818733, 
    1.818734, 1.818733, 1.818734, 1.818734, 1.818734, 1.818736, 1.818735, 
    1.818736, 1.818735, 1.818725, 1.818726, 1.818726, 1.818726, 1.818726, 
    1.818727, 1.818728, 1.81873, 1.818729, 1.81873, 1.818729, 1.818729, 
    1.818731, 1.818729, 1.818732, 1.81873, 1.818734, 1.818732, 1.818734, 
    1.818733, 1.818734, 1.818735, 1.818735, 1.818736, 1.818736, 1.818737, 
    1.818727, 1.818727, 1.818727, 1.818728, 1.818728, 1.818729, 1.818731, 
    1.81873, 1.818732, 1.818732, 1.81873, 1.818731, 1.818728, 1.818728, 
    1.818728, 1.818727, 1.818731, 1.818729, 1.818732, 1.818731, 1.818735, 
    1.818733, 1.818736, 1.818737, 1.818739, 1.81874, 1.818728, 1.818727, 
    1.818728, 1.818729, 1.81873, 1.818731, 1.818731, 1.818732, 1.818732, 
    1.818733, 1.818732, 1.818733, 1.818728, 1.818731, 1.818727, 1.818728, 
    1.818729, 1.818729, 1.81873, 1.818731, 1.818733, 1.818732, 1.818737, 
    1.818735, 1.818741, 1.818739, 1.818727, 1.818728, 1.81873, 1.818729, 
    1.818731, 1.818732, 1.818733, 1.818733, 1.818733, 1.818734, 1.818733, 
    1.818734, 1.818731, 1.818733, 1.818729, 1.81873, 1.81873, 1.818729, 
    1.818731, 1.818732, 1.818732, 1.818732, 1.818733, 1.818731, 1.818737, 
    1.818734, 1.818728, 1.818729, 1.81873, 1.818729, 1.818732, 1.818731, 
    1.818734, 1.818733, 1.818734, 1.818734, 1.818734, 1.818733, 1.818732, 
    1.818731, 1.81873, 1.818729, 1.818729, 1.81873, 1.818732, 1.818733, 
    1.818733, 1.818734, 1.818731, 1.818733, 1.818732, 1.818733, 1.81873, 
    1.818733, 1.81873, 1.81873, 1.818731, 1.818733, 1.818733, 1.818733, 
    1.818733, 1.818732, 1.818732, 1.818731, 1.818731, 1.81873, 1.81873, 
    1.81873, 1.81873, 1.818732, 1.818733, 1.818735, 1.818735, 1.818737, 
    1.818735, 1.818737, 1.818736, 1.818739, 1.818733, 1.818735, 1.818731, 
    1.818731, 1.818732, 1.818734, 1.818733, 1.818735, 1.818732, 1.81873, 
    1.81873, 1.818729, 1.81873, 1.81873, 1.818731, 1.81873, 1.818732, 
    1.818731, 1.818734, 1.818735, 1.818737, 1.818739, 1.81874, 1.818741, 
    1.818741, 1.818741,
  1.818671, 1.818673, 1.818673, 1.818674, 1.818673, 1.818674, 1.818671, 
    1.818673, 1.818672, 1.818671, 1.818677, 1.818674, 1.81868, 1.818678, 
    1.818683, 1.81868, 1.818683, 1.818683, 1.818685, 1.818684, 1.818687, 
    1.818685, 1.818688, 1.818686, 1.818687, 1.818685, 1.818675, 1.818677, 
    1.818675, 1.818675, 1.818675, 1.818673, 1.818673, 1.818671, 1.818671, 
    1.818672, 1.818675, 1.818674, 1.818676, 1.818676, 1.818679, 1.818678, 
    1.818682, 1.818681, 1.818684, 1.818683, 1.818684, 1.818684, 1.818684, 
    1.818683, 1.818683, 1.818682, 1.818678, 1.818679, 1.818675, 1.818673, 
    1.818672, 1.818671, 1.818671, 1.818671, 1.818672, 1.818674, 1.818675, 
    1.818676, 1.818676, 1.818678, 1.81868, 1.818682, 1.818682, 1.818683, 
    1.818683, 1.818684, 1.818684, 1.818685, 1.818682, 1.818684, 1.818681, 
    1.818682, 1.818677, 1.818674, 1.818673, 1.818673, 1.818671, 1.818672, 
    1.818672, 1.818673, 1.818674, 1.818673, 1.818676, 1.818675, 1.81868, 
    1.818678, 1.818683, 1.818682, 1.818684, 1.818683, 1.818684, 1.818683, 
    1.818685, 1.818686, 1.818685, 1.818686, 1.818683, 1.818684, 1.818673, 
    1.818673, 1.818674, 1.818672, 1.818672, 1.818671, 1.818672, 1.818673, 
    1.818674, 1.818674, 1.818675, 1.818676, 1.818678, 1.81868, 1.818682, 
    1.818683, 1.818682, 1.818683, 1.818682, 1.818682, 1.818685, 1.818683, 
    1.818686, 1.818686, 1.818685, 1.818686, 1.818673, 1.818673, 1.818672, 
    1.818673, 1.818671, 1.818672, 1.818672, 1.818675, 1.818675, 1.818676, 
    1.818677, 1.818678, 1.81868, 1.818682, 1.818683, 1.818683, 1.818683, 
    1.818684, 1.818683, 1.818684, 1.818684, 1.818683, 1.818686, 1.818685, 
    1.818686, 1.818686, 1.818673, 1.818674, 1.818673, 1.818674, 1.818674, 
    1.818676, 1.818676, 1.818679, 1.818678, 1.81868, 1.818678, 1.818678, 
    1.81868, 1.818678, 1.818682, 1.818679, 1.818684, 1.818681, 1.818684, 
    1.818683, 1.818684, 1.818685, 1.818686, 1.818687, 1.818687, 1.818688, 
    1.818675, 1.818675, 1.818675, 1.818676, 1.818677, 1.818678, 1.81868, 
    1.81868, 1.818681, 1.818681, 1.818679, 1.818681, 1.818676, 1.818677, 
    1.818676, 1.818675, 1.81868, 1.818677, 1.818682, 1.818681, 1.818685, 
    1.818683, 1.818687, 1.818688, 1.81869, 1.818692, 1.818676, 1.818675, 
    1.818676, 1.818678, 1.818679, 1.818681, 1.818681, 1.818681, 1.818682, 
    1.818683, 1.818681, 1.818683, 1.818677, 1.81868, 1.818675, 1.818677, 
    1.818678, 1.818677, 1.818679, 1.81868, 1.818682, 1.818681, 1.818688, 
    1.818685, 1.818693, 1.818691, 1.818675, 1.818676, 1.818678, 1.818677, 
    1.818681, 1.818682, 1.818682, 1.818683, 1.818683, 1.818684, 1.818683, 
    1.818684, 1.818681, 1.818682, 1.818678, 1.818679, 1.818679, 1.818678, 
    1.81868, 1.818681, 1.818681, 1.818682, 1.818683, 1.818681, 1.818688, 
    1.818684, 1.818677, 1.818678, 1.818678, 1.818678, 1.818681, 1.81868, 
    1.818684, 1.818683, 1.818684, 1.818684, 1.818684, 1.818682, 1.818682, 
    1.81868, 1.818679, 1.818678, 1.818678, 1.818679, 1.818681, 1.818683, 
    1.818683, 1.818684, 1.818681, 1.818682, 1.818681, 1.818683, 1.81868, 
    1.818683, 1.818679, 1.818679, 1.81868, 1.818682, 1.818683, 1.818683, 
    1.818683, 1.818681, 1.818681, 1.81868, 1.81868, 1.818679, 1.818678, 
    1.818679, 1.81868, 1.818681, 1.818683, 1.818685, 1.818685, 1.818687, 
    1.818686, 1.818688, 1.818686, 1.81869, 1.818683, 1.818686, 1.81868, 
    1.818681, 1.818682, 1.818684, 1.818683, 1.818685, 1.818681, 1.818679, 
    1.818679, 1.818678, 1.818679, 1.818679, 1.81868, 1.818679, 1.818681, 
    1.81868, 1.818684, 1.818685, 1.818688, 1.81869, 1.818692, 1.818693, 
    1.818693, 1.818693,
  1.818642, 1.818644, 1.818643, 1.818645, 1.818644, 1.818645, 1.818642, 
    1.818644, 1.818643, 1.818642, 1.818648, 1.818645, 1.818651, 1.818649, 
    1.818654, 1.818651, 1.818655, 1.818654, 1.818657, 1.818656, 1.818659, 
    1.818657, 1.81866, 1.818658, 1.818659, 1.818657, 1.818646, 1.818648, 
    1.818645, 1.818646, 1.818646, 1.818644, 1.818643, 1.818642, 1.818642, 
    1.818643, 1.818646, 1.818645, 1.818647, 1.818647, 1.81865, 1.818649, 
    1.818653, 1.818652, 1.818656, 1.818655, 1.818656, 1.818656, 1.818656, 
    1.818655, 1.818655, 1.818654, 1.818649, 1.81865, 1.818646, 1.818644, 
    1.818642, 1.818641, 1.818641, 1.818641, 1.818643, 1.818645, 1.818646, 
    1.818647, 1.818647, 1.81865, 1.818651, 1.818654, 1.818653, 1.818654, 
    1.818655, 1.818656, 1.818656, 1.818657, 1.818654, 1.818656, 1.818653, 
    1.818654, 1.818648, 1.818645, 1.818644, 1.818643, 1.818641, 1.818643, 
    1.818642, 1.818644, 1.818644, 1.818644, 1.818647, 1.818646, 1.818651, 
    1.818649, 1.818655, 1.818653, 1.818655, 1.818654, 1.818656, 1.818654, 
    1.818657, 1.818657, 1.818657, 1.818658, 1.818654, 1.818656, 1.818644, 
    1.818644, 1.818644, 1.818643, 1.818643, 1.818642, 1.818643, 1.818643, 
    1.818644, 1.818645, 1.818646, 1.818648, 1.818649, 1.818652, 1.818653, 
    1.818655, 1.818654, 1.818655, 1.818654, 1.818653, 1.818657, 1.818655, 
    1.818658, 1.818658, 1.818657, 1.818658, 1.818644, 1.818644, 1.818642, 
    1.818643, 1.818641, 1.818642, 1.818643, 1.818646, 1.818646, 1.818647, 
    1.818648, 1.818649, 1.818651, 1.818653, 1.818655, 1.818655, 1.818655, 
    1.818655, 1.818654, 1.818655, 1.818656, 1.818655, 1.818658, 1.818657, 
    1.818658, 1.818658, 1.818644, 1.818645, 1.818644, 1.818645, 1.818644, 
    1.818646, 1.818647, 1.81865, 1.818649, 1.818651, 1.818649, 1.818649, 
    1.818651, 1.818649, 1.818653, 1.81865, 1.818655, 1.818653, 1.818655, 
    1.818655, 1.818656, 1.818656, 1.818657, 1.818659, 1.818659, 1.81866, 
    1.818645, 1.818646, 1.818646, 1.818647, 1.818648, 1.818649, 1.818652, 
    1.818651, 1.818653, 1.818653, 1.81865, 1.818652, 1.818647, 1.818648, 
    1.818647, 1.818646, 1.818651, 1.818648, 1.818653, 1.818652, 1.818656, 
    1.818654, 1.818658, 1.81866, 1.818662, 1.818664, 1.818647, 1.818646, 
    1.818647, 1.818649, 1.81865, 1.818652, 1.818652, 1.818653, 1.818653, 
    1.818654, 1.818653, 1.818654, 1.818648, 1.818651, 1.818646, 1.818648, 
    1.818649, 1.818648, 1.818651, 1.818651, 1.818654, 1.818653, 1.81866, 
    1.818657, 1.818666, 1.818663, 1.818646, 1.818647, 1.81865, 1.818648, 
    1.818652, 1.818653, 1.818654, 1.818655, 1.818655, 1.818655, 1.818655, 
    1.818655, 1.818652, 1.818654, 1.818649, 1.81865, 1.81865, 1.818649, 
    1.818651, 1.818653, 1.818653, 1.818653, 1.818655, 1.818652, 1.81866, 
    1.818655, 1.818648, 1.818649, 1.81865, 1.818649, 1.818653, 1.818652, 
    1.818655, 1.818654, 1.818656, 1.818655, 1.818655, 1.818654, 1.818653, 
    1.818652, 1.81865, 1.818649, 1.818649, 1.81865, 1.818653, 1.818655, 
    1.818654, 1.818656, 1.818652, 1.818654, 1.818653, 1.818655, 1.818651, 
    1.818654, 1.81865, 1.81865, 1.818651, 1.818654, 1.818654, 1.818655, 
    1.818654, 1.818653, 1.818653, 1.818651, 1.818651, 1.81865, 1.81865, 
    1.81865, 1.818651, 1.818653, 1.818655, 1.818656, 1.818657, 1.818659, 
    1.818657, 1.81866, 1.818658, 1.818662, 1.818654, 1.818658, 1.818652, 
    1.818652, 1.818653, 1.818656, 1.818655, 1.818656, 1.818653, 1.818651, 
    1.81865, 1.818649, 1.81865, 1.81865, 1.818651, 1.818651, 1.818653, 
    1.818652, 1.818655, 1.818656, 1.81866, 1.818662, 1.818664, 1.818665, 
    1.818666, 1.818666,
  1.818619, 1.818621, 1.818621, 1.818622, 1.818621, 1.818622, 1.818619, 
    1.818621, 1.81862, 1.818619, 1.818625, 1.818622, 1.818629, 1.818627, 
    1.818632, 1.818628, 1.818632, 1.818632, 1.818634, 1.818633, 1.818636, 
    1.818634, 1.818638, 1.818636, 1.818636, 1.818634, 1.818623, 1.818625, 
    1.818623, 1.818623, 1.818623, 1.818621, 1.81862, 1.818619, 1.818619, 
    1.81862, 1.818623, 1.818622, 1.818625, 1.818625, 1.818627, 1.818626, 
    1.818631, 1.81863, 1.818633, 1.818632, 1.818633, 1.818633, 1.818633, 
    1.818632, 1.818632, 1.818631, 1.818626, 1.818628, 1.818624, 1.818621, 
    1.818619, 1.818618, 1.818618, 1.818619, 1.81862, 1.818622, 1.818623, 
    1.818624, 1.818625, 1.818627, 1.818628, 1.818631, 1.818631, 1.818632, 
    1.818632, 1.818634, 1.818633, 1.818634, 1.818631, 1.818633, 1.81863, 
    1.818631, 1.818625, 1.818622, 1.818622, 1.818621, 1.818618, 1.81862, 
    1.818619, 1.818621, 1.818622, 1.818621, 1.818624, 1.818623, 1.818628, 
    1.818626, 1.818632, 1.818631, 1.818633, 1.818632, 1.818633, 1.818632, 
    1.818634, 1.818635, 1.818635, 1.818636, 1.818632, 1.818633, 1.818621, 
    1.818621, 1.818622, 1.81862, 1.81862, 1.818619, 1.81862, 1.81862, 
    1.818622, 1.818622, 1.818623, 1.818625, 1.818627, 1.818629, 1.818631, 
    1.818632, 1.818631, 1.818632, 1.818631, 1.818631, 1.818635, 1.818632, 
    1.818636, 1.818636, 1.818634, 1.818636, 1.818621, 1.818621, 1.818619, 
    1.818621, 1.818619, 1.81862, 1.81862, 1.818623, 1.818623, 1.818624, 
    1.818625, 1.818626, 1.818629, 1.818631, 1.818632, 1.818632, 1.818632, 
    1.818633, 1.818632, 1.818633, 1.818633, 1.818632, 1.818635, 1.818635, 
    1.818636, 1.818635, 1.818621, 1.818622, 1.818621, 1.818622, 1.818622, 
    1.818624, 1.818624, 1.818627, 1.818626, 1.818628, 1.818626, 1.818627, 
    1.818628, 1.818627, 1.81863, 1.818628, 1.818633, 1.81863, 1.818633, 
    1.818632, 1.818633, 1.818634, 1.818635, 1.818637, 1.818636, 1.818638, 
    1.818623, 1.818624, 1.818624, 1.818624, 1.818625, 1.818627, 1.818629, 
    1.818628, 1.81863, 1.81863, 1.818628, 1.818629, 1.818624, 1.818625, 
    1.818625, 1.818623, 1.818628, 1.818626, 1.818631, 1.818629, 1.818634, 
    1.818632, 1.818636, 1.818638, 1.81864, 1.818642, 1.818624, 1.818624, 
    1.818625, 1.818626, 1.818627, 1.818629, 1.81863, 1.81863, 1.818631, 
    1.818632, 1.81863, 1.818632, 1.818625, 1.818629, 1.818623, 1.818625, 
    1.818626, 1.818626, 1.818628, 1.818629, 1.818631, 1.81863, 1.818637, 
    1.818634, 1.818643, 1.818641, 1.818623, 1.818624, 1.818627, 1.818626, 
    1.81863, 1.81863, 1.818631, 1.818632, 1.818632, 1.818633, 1.818632, 
    1.818633, 1.818629, 1.818631, 1.818627, 1.818628, 1.818627, 1.818627, 
    1.818628, 1.81863, 1.81863, 1.818631, 1.818632, 1.81863, 1.818638, 
    1.818633, 1.818625, 1.818627, 1.818627, 1.818626, 1.81863, 1.818629, 
    1.818633, 1.818632, 1.818634, 1.818633, 1.818633, 1.818631, 1.818631, 
    1.818629, 1.818627, 1.818626, 1.818627, 1.818628, 1.81863, 1.818632, 
    1.818632, 1.818633, 1.818629, 1.818631, 1.81863, 1.818632, 1.818628, 
    1.818632, 1.818627, 1.818628, 1.818629, 1.818631, 1.818632, 1.818632, 
    1.818632, 1.81863, 1.81863, 1.818629, 1.818628, 1.818628, 1.818627, 
    1.818628, 1.818628, 1.81863, 1.818632, 1.818634, 1.818634, 1.818637, 
    1.818635, 1.818638, 1.818635, 1.81864, 1.818632, 1.818635, 1.818629, 
    1.81863, 1.818631, 1.818634, 1.818632, 1.818634, 1.81863, 1.818628, 
    1.818627, 1.818626, 1.818627, 1.818627, 1.818628, 1.818628, 1.81863, 
    1.818629, 1.818633, 1.818634, 1.818638, 1.81864, 1.818642, 1.818643, 
    1.818643, 1.818644,
  1.818569, 1.818571, 1.818571, 1.818572, 1.818571, 1.818572, 1.81857, 
    1.818571, 1.81857, 1.818569, 1.818575, 1.818572, 1.818578, 1.818576, 
    1.818581, 1.818578, 1.818581, 1.81858, 1.818582, 1.818582, 1.818584, 
    1.818583, 1.818586, 1.818584, 1.818584, 1.818583, 1.818573, 1.818575, 
    1.818573, 1.818573, 1.818573, 1.818571, 1.818571, 1.818569, 1.818569, 
    1.81857, 1.818573, 1.818572, 1.818574, 1.818574, 1.818577, 1.818576, 
    1.81858, 1.818578, 1.818582, 1.818581, 1.818582, 1.818582, 1.818582, 
    1.818581, 1.818581, 1.81858, 1.818576, 1.818577, 1.818573, 1.818571, 
    1.81857, 1.818569, 1.818569, 1.818569, 1.81857, 1.818572, 1.818573, 
    1.818574, 1.818574, 1.818576, 1.818577, 1.81858, 1.818579, 1.81858, 
    1.818581, 1.818582, 1.818582, 1.818583, 1.81858, 1.818582, 1.818579, 
    1.81858, 1.818574, 1.818572, 1.818571, 1.818571, 1.818569, 1.81857, 
    1.81857, 1.818571, 1.818572, 1.818571, 1.818574, 1.818573, 1.818578, 
    1.818575, 1.818581, 1.81858, 1.818581, 1.81858, 1.818582, 1.818581, 
    1.818583, 1.818583, 1.818583, 1.818584, 1.81858, 1.818582, 1.818571, 
    1.818571, 1.818572, 1.81857, 1.81857, 1.818569, 1.81857, 1.81857, 
    1.818572, 1.818572, 1.818573, 1.818574, 1.818576, 1.818578, 1.81858, 
    1.818581, 1.81858, 1.818581, 1.81858, 1.81858, 1.818583, 1.818581, 
    1.818584, 1.818584, 1.818583, 1.818584, 1.818571, 1.818571, 1.81857, 
    1.818571, 1.818569, 1.81857, 1.81857, 1.818573, 1.818573, 1.818574, 
    1.818575, 1.818576, 1.818578, 1.818579, 1.818581, 1.818581, 1.818581, 
    1.818581, 1.81858, 1.818581, 1.818582, 1.818581, 1.818584, 1.818583, 
    1.818584, 1.818583, 1.818571, 1.818572, 1.818571, 1.818572, 1.818572, 
    1.818573, 1.818574, 1.818577, 1.818576, 1.818577, 1.818576, 1.818576, 
    1.818577, 1.818576, 1.818579, 1.818577, 1.818581, 1.818579, 1.818581, 
    1.818581, 1.818582, 1.818582, 1.818583, 1.818585, 1.818584, 1.818586, 
    1.818573, 1.818573, 1.818573, 1.818574, 1.818575, 1.818576, 1.818578, 
    1.818577, 1.818579, 1.818579, 1.818577, 1.818578, 1.818574, 1.818575, 
    1.818574, 1.818573, 1.818578, 1.818575, 1.81858, 1.818578, 1.818582, 
    1.81858, 1.818584, 1.818586, 1.818587, 1.818589, 1.818574, 1.818573, 
    1.818574, 1.818576, 1.818577, 1.818578, 1.818579, 1.818579, 1.81858, 
    1.81858, 1.818579, 1.818581, 1.818575, 1.818578, 1.818573, 1.818574, 
    1.818576, 1.818575, 1.818577, 1.818578, 1.81858, 1.818579, 1.818586, 
    1.818583, 1.818591, 1.818588, 1.818573, 1.818574, 1.818576, 1.818575, 
    1.818578, 1.818579, 1.81858, 1.818581, 1.818581, 1.818581, 1.818581, 
    1.818581, 1.818578, 1.81858, 1.818576, 1.818577, 1.818576, 1.818576, 
    1.818577, 1.818579, 1.818579, 1.81858, 1.818581, 1.818578, 1.818586, 
    1.818581, 1.818575, 1.818576, 1.818576, 1.818576, 1.818579, 1.818578, 
    1.818581, 1.818581, 1.818582, 1.818581, 1.818581, 1.81858, 1.81858, 
    1.818578, 1.818577, 1.818576, 1.818576, 1.818577, 1.818579, 1.818581, 
    1.818581, 1.818582, 1.818578, 1.81858, 1.818579, 1.818581, 1.818577, 
    1.81858, 1.818577, 1.818577, 1.818578, 1.81858, 1.81858, 1.818581, 
    1.818581, 1.818579, 1.818579, 1.818578, 1.818578, 1.818577, 1.818576, 
    1.818577, 1.818577, 1.818579, 1.818581, 1.818582, 1.818583, 1.818585, 
    1.818583, 1.818586, 1.818584, 1.818588, 1.81858, 1.818583, 1.818578, 
    1.818579, 1.81858, 1.818582, 1.818581, 1.818582, 1.818579, 1.818577, 
    1.818577, 1.818576, 1.818577, 1.818577, 1.818577, 1.818577, 1.818579, 
    1.818578, 1.818581, 1.818582, 1.818586, 1.818588, 1.81859, 1.81859, 
    1.818591, 1.818591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.297841e-09, 1.303568e-09, 1.302455e-09, 1.307074e-09, 1.304511e-09, 
    1.307536e-09, 1.299002e-09, 1.303795e-09, 1.300735e-09, 1.298357e-09, 
    1.316038e-09, 1.30728e-09, 1.325137e-09, 1.319551e-09, 1.333584e-09, 
    1.324267e-09, 1.335463e-09, 1.333316e-09, 1.33978e-09, 1.337928e-09, 
    1.346196e-09, 1.340634e-09, 1.350482e-09, 1.344868e-09, 1.345746e-09, 
    1.340451e-09, 1.309042e-09, 1.314947e-09, 1.308692e-09, 1.309534e-09, 
    1.309157e-09, 1.304564e-09, 1.30225e-09, 1.297404e-09, 1.298283e-09, 
    1.301843e-09, 1.309913e-09, 1.307174e-09, 1.314078e-09, 1.313922e-09, 
    1.321609e-09, 1.318143e-09, 1.331065e-09, 1.327392e-09, 1.338005e-09, 
    1.335336e-09, 1.33788e-09, 1.337109e-09, 1.33789e-09, 1.333975e-09, 
    1.335652e-09, 1.332208e-09, 1.318792e-09, 1.322735e-09, 1.310977e-09, 
    1.303907e-09, 1.299212e-09, 1.295881e-09, 1.296352e-09, 1.29725e-09, 
    1.301864e-09, 1.306202e-09, 1.309509e-09, 1.311721e-09, 1.3139e-09, 
    1.320496e-09, 1.323988e-09, 1.331807e-09, 1.330396e-09, 1.332787e-09, 
    1.33507e-09, 1.338905e-09, 1.338274e-09, 1.339963e-09, 1.332724e-09, 
    1.337535e-09, 1.329593e-09, 1.331765e-09, 1.314491e-09, 1.307913e-09, 
    1.305116e-09, 1.302669e-09, 1.296714e-09, 1.300826e-09, 1.299205e-09, 
    1.303062e-09, 1.305512e-09, 1.3043e-09, 1.311781e-09, 1.308873e-09, 
    1.324195e-09, 1.317595e-09, 1.334804e-09, 1.330686e-09, 1.335791e-09, 
    1.333186e-09, 1.33765e-09, 1.333633e-09, 1.340592e-09, 1.342108e-09, 
    1.341072e-09, 1.34505e-09, 1.33341e-09, 1.33788e-09, 1.304266e-09, 
    1.304464e-09, 1.305385e-09, 1.301336e-09, 1.301089e-09, 1.297379e-09, 
    1.30068e-09, 1.302086e-09, 1.305654e-09, 1.307765e-09, 1.309772e-09, 
    1.314184e-09, 1.319111e-09, 1.326002e-09, 1.330953e-09, 1.334272e-09, 
    1.332237e-09, 1.334033e-09, 1.332025e-09, 1.331083e-09, 1.34154e-09, 
    1.335668e-09, 1.344478e-09, 1.343991e-09, 1.340003e-09, 1.344045e-09, 
    1.304603e-09, 1.303465e-09, 1.299516e-09, 1.302607e-09, 1.296975e-09, 
    1.300127e-09, 1.30194e-09, 1.308933e-09, 1.31047e-09, 1.311895e-09, 
    1.314709e-09, 1.318321e-09, 1.324657e-09, 1.33017e-09, 1.335203e-09, 
    1.334835e-09, 1.334964e-09, 1.336089e-09, 1.333304e-09, 1.336546e-09, 
    1.33709e-09, 1.335667e-09, 1.343925e-09, 1.341566e-09, 1.34398e-09, 
    1.342444e-09, 1.303835e-09, 1.305749e-09, 1.304715e-09, 1.30666e-09, 
    1.305289e-09, 1.311382e-09, 1.313209e-09, 1.321758e-09, 1.31825e-09, 
    1.323833e-09, 1.318817e-09, 1.319706e-09, 1.324015e-09, 1.319088e-09, 
    1.329866e-09, 1.322558e-09, 1.336133e-09, 1.328834e-09, 1.33659e-09, 
    1.335182e-09, 1.337513e-09, 1.339601e-09, 1.342229e-09, 1.347077e-09, 
    1.345954e-09, 1.350008e-09, 1.308603e-09, 1.311085e-09, 1.310867e-09, 
    1.313465e-09, 1.315387e-09, 1.319552e-09, 1.326233e-09, 1.323721e-09, 
    1.328333e-09, 1.329259e-09, 1.322252e-09, 1.326554e-09, 1.312747e-09, 
    1.314977e-09, 1.31365e-09, 1.308798e-09, 1.324299e-09, 1.316344e-09, 
    1.331035e-09, 1.326725e-09, 1.339304e-09, 1.333048e-09, 1.345336e-09, 
    1.350589e-09, 1.355534e-09, 1.361312e-09, 1.31244e-09, 1.310754e-09, 
    1.313774e-09, 1.317953e-09, 1.321832e-09, 1.326987e-09, 1.327515e-09, 
    1.328481e-09, 1.330983e-09, 1.333087e-09, 1.328786e-09, 1.333614e-09, 
    1.315494e-09, 1.32499e-09, 1.310116e-09, 1.314594e-09, 1.317707e-09, 
    1.316342e-09, 1.323433e-09, 1.325105e-09, 1.331897e-09, 1.328386e-09, 
    1.349292e-09, 1.340042e-09, 1.365712e-09, 1.358538e-09, 1.310164e-09, 
    1.312435e-09, 1.320338e-09, 1.316577e-09, 1.327332e-09, 1.329979e-09, 
    1.332131e-09, 1.334882e-09, 1.335179e-09, 1.336809e-09, 1.334138e-09, 
    1.336704e-09, 1.326998e-09, 1.331335e-09, 1.319434e-09, 1.322331e-09, 
    1.320999e-09, 1.319537e-09, 1.324048e-09, 1.328854e-09, 1.328957e-09, 
    1.330498e-09, 1.33484e-09, 1.327375e-09, 1.350486e-09, 1.336212e-09, 
    1.314911e-09, 1.319284e-09, 1.319909e-09, 1.318215e-09, 1.329714e-09, 
    1.325547e-09, 1.33677e-09, 1.333737e-09, 1.338706e-09, 1.336237e-09, 
    1.335873e-09, 1.332702e-09, 1.330727e-09, 1.325738e-09, 1.321679e-09, 
    1.318461e-09, 1.319209e-09, 1.322745e-09, 1.329148e-09, 1.335206e-09, 
    1.333879e-09, 1.338329e-09, 1.326552e-09, 1.33149e-09, 1.329581e-09, 
    1.334558e-09, 1.323654e-09, 1.332938e-09, 1.321281e-09, 1.322303e-09, 
    1.325464e-09, 1.331825e-09, 1.333232e-09, 1.334735e-09, 1.333808e-09, 
    1.329311e-09, 1.328574e-09, 1.325388e-09, 1.324508e-09, 1.32208e-09, 
    1.32007e-09, 1.321906e-09, 1.323835e-09, 1.329313e-09, 1.334249e-09, 
    1.339631e-09, 1.340948e-09, 1.347237e-09, 1.342118e-09, 1.350565e-09, 
    1.343383e-09, 1.355817e-09, 1.333477e-09, 1.343172e-09, 1.325608e-09, 
    1.3275e-09, 1.330922e-09, 1.338772e-09, 1.334535e-09, 1.33949e-09, 
    1.328545e-09, 1.322866e-09, 1.321398e-09, 1.318657e-09, 1.32146e-09, 
    1.321232e-09, 1.323915e-09, 1.323053e-09, 1.329494e-09, 1.326034e-09, 
    1.335864e-09, 1.339451e-09, 1.349583e-09, 1.355794e-09, 1.362118e-09, 
    1.364909e-09, 1.365759e-09, 1.366114e-09 ;

 SOIL2_HR_S3 =
  9.270293e-11, 9.311198e-11, 9.303247e-11, 9.336239e-11, 9.317938e-11, 
    9.339542e-11, 9.278587e-11, 9.312821e-11, 9.290967e-11, 9.273977e-11, 
    9.400268e-11, 9.337712e-11, 9.465263e-11, 9.425361e-11, 9.525603e-11, 
    9.459052e-11, 9.539023e-11, 9.523686e-11, 9.569855e-11, 9.556628e-11, 
    9.615683e-11, 9.57596e-11, 9.646299e-11, 9.606198e-11, 9.612471e-11, 
    9.574649e-11, 9.350302e-11, 9.392478e-11, 9.347803e-11, 9.353818e-11, 
    9.351119e-11, 9.318316e-11, 9.301784e-11, 9.267168e-11, 9.273453e-11, 
    9.298878e-11, 9.356522e-11, 9.336956e-11, 9.386273e-11, 9.385159e-11, 
    9.440067e-11, 9.41531e-11, 9.507604e-11, 9.481373e-11, 9.557181e-11, 
    9.538115e-11, 9.556285e-11, 9.550775e-11, 9.556356e-11, 9.528395e-11, 
    9.540374e-11, 9.515771e-11, 9.419946e-11, 9.448106e-11, 9.364121e-11, 
    9.313622e-11, 9.280088e-11, 9.256291e-11, 9.259655e-11, 9.266068e-11, 
    9.299026e-11, 9.330017e-11, 9.353635e-11, 9.369432e-11, 9.385e-11, 
    9.432115e-11, 9.457059e-11, 9.512908e-11, 9.50283e-11, 9.519904e-11, 
    9.536218e-11, 9.563605e-11, 9.559098e-11, 9.571164e-11, 9.519455e-11, 
    9.55382e-11, 9.49709e-11, 9.512605e-11, 9.389224e-11, 9.342235e-11, 
    9.322256e-11, 9.304775e-11, 9.262242e-11, 9.291613e-11, 9.280034e-11, 
    9.307583e-11, 9.325088e-11, 9.316431e-11, 9.369865e-11, 9.34909e-11, 
    9.458537e-11, 9.411392e-11, 9.534315e-11, 9.504899e-11, 9.541366e-11, 
    9.522758e-11, 9.554642e-11, 9.525947e-11, 9.575656e-11, 9.586482e-11, 
    9.579083e-11, 9.607501e-11, 9.524356e-11, 9.556284e-11, 9.316188e-11, 
    9.317599e-11, 9.324178e-11, 9.295261e-11, 9.293492e-11, 9.266996e-11, 
    9.290573e-11, 9.300613e-11, 9.326103e-11, 9.34118e-11, 9.355512e-11, 
    9.387026e-11, 9.422221e-11, 9.471442e-11, 9.506806e-11, 9.530512e-11, 
    9.515976e-11, 9.528809e-11, 9.514463e-11, 9.50774e-11, 9.582427e-11, 
    9.540486e-11, 9.603414e-11, 9.599933e-11, 9.571451e-11, 9.600325e-11, 
    9.318591e-11, 9.310466e-11, 9.282256e-11, 9.304333e-11, 9.26411e-11, 
    9.286624e-11, 9.299569e-11, 9.349523e-11, 9.360501e-11, 9.370677e-11, 
    9.390779e-11, 9.416577e-11, 9.461834e-11, 9.501214e-11, 9.537168e-11, 
    9.534533e-11, 9.535461e-11, 9.543492e-11, 9.523598e-11, 9.546758e-11, 
    9.550644e-11, 9.540482e-11, 9.599466e-11, 9.582615e-11, 9.599858e-11, 
    9.588887e-11, 9.313107e-11, 9.326779e-11, 9.319391e-11, 9.333283e-11, 
    9.323496e-11, 9.367016e-11, 9.380065e-11, 9.441128e-11, 9.416069e-11, 
    9.455953e-11, 9.420121e-11, 9.426469e-11, 9.457251e-11, 9.422058e-11, 
    9.499042e-11, 9.446845e-11, 9.543803e-11, 9.491674e-11, 9.54707e-11, 
    9.537012e-11, 9.553666e-11, 9.568581e-11, 9.587351e-11, 9.621975e-11, 
    9.613958e-11, 9.642916e-11, 9.347162e-11, 9.364895e-11, 9.363335e-11, 
    9.381895e-11, 9.39562e-11, 9.425372e-11, 9.473091e-11, 9.455147e-11, 
    9.488092e-11, 9.494705e-11, 9.444655e-11, 9.475383e-11, 9.376765e-11, 
    9.392696e-11, 9.383211e-11, 9.34856e-11, 9.45928e-11, 9.402455e-11, 
    9.50739e-11, 9.476604e-11, 9.566455e-11, 9.521768e-11, 9.609544e-11, 
    9.647065e-11, 9.682385e-11, 9.723657e-11, 9.374575e-11, 9.362525e-11, 
    9.384102e-11, 9.413953e-11, 9.441654e-11, 9.478482e-11, 9.482251e-11, 
    9.48915e-11, 9.507022e-11, 9.522049e-11, 9.49133e-11, 9.525816e-11, 
    9.396388e-11, 9.464213e-11, 9.357969e-11, 9.389958e-11, 9.412194e-11, 
    9.402441e-11, 9.453096e-11, 9.465035e-11, 9.513552e-11, 9.488472e-11, 
    9.637803e-11, 9.57173e-11, 9.755088e-11, 9.703843e-11, 9.358315e-11, 
    9.374534e-11, 9.430983e-11, 9.404125e-11, 9.480941e-11, 9.49985e-11, 
    9.515223e-11, 9.534873e-11, 9.536995e-11, 9.548638e-11, 9.529559e-11, 
    9.547885e-11, 9.47856e-11, 9.50954e-11, 9.424532e-11, 9.44522e-11, 
    9.435704e-11, 9.425263e-11, 9.457485e-11, 9.491813e-11, 9.492549e-11, 
    9.503556e-11, 9.53457e-11, 9.481253e-11, 9.646326e-11, 9.544373e-11, 
    9.39222e-11, 9.42346e-11, 9.427924e-11, 9.415822e-11, 9.497955e-11, 
    9.468194e-11, 9.548354e-11, 9.52669e-11, 9.562188e-11, 9.544548e-11, 
    9.541953e-11, 9.519297e-11, 9.505192e-11, 9.469558e-11, 9.440566e-11, 
    9.417579e-11, 9.422924e-11, 9.448176e-11, 9.493914e-11, 9.537186e-11, 
    9.527707e-11, 9.55949e-11, 9.475371e-11, 9.510642e-11, 9.497009e-11, 
    9.532557e-11, 9.45467e-11, 9.520987e-11, 9.437718e-11, 9.445019e-11, 
    9.467603e-11, 9.513032e-11, 9.523087e-11, 9.533818e-11, 9.527197e-11, 
    9.495076e-11, 9.489814e-11, 9.467055e-11, 9.46077e-11, 9.443429e-11, 
    9.429073e-11, 9.442189e-11, 9.455964e-11, 9.495089e-11, 9.530349e-11, 
    9.568794e-11, 9.578203e-11, 9.623121e-11, 9.586556e-11, 9.646894e-11, 
    9.59559e-11, 9.684404e-11, 9.524835e-11, 9.594085e-11, 9.468631e-11, 
    9.482146e-11, 9.506589e-11, 9.562658e-11, 9.53239e-11, 9.567789e-11, 
    9.489608e-11, 9.449046e-11, 9.438554e-11, 9.418975e-11, 9.439002e-11, 
    9.437373e-11, 9.456536e-11, 9.450378e-11, 9.496388e-11, 9.471673e-11, 
    9.541887e-11, 9.56751e-11, 9.639881e-11, 9.684245e-11, 9.729411e-11, 
    9.749351e-11, 9.75542e-11, 9.757958e-11 ;

 SOIL3C =
  5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611 ;

 SOIL3C_TO_SOIL1C =
  2.559307e-11, 2.570598e-11, 2.568403e-11, 2.57751e-11, 2.572458e-11, 
    2.578421e-11, 2.561596e-11, 2.571046e-11, 2.565014e-11, 2.560324e-11, 
    2.595182e-11, 2.577916e-11, 2.613122e-11, 2.602108e-11, 2.629777e-11, 
    2.611408e-11, 2.633481e-11, 2.629248e-11, 2.641991e-11, 2.63834e-11, 
    2.65464e-11, 2.643676e-11, 2.66309e-11, 2.652022e-11, 2.653753e-11, 
    2.643314e-11, 2.581391e-11, 2.593033e-11, 2.580701e-11, 2.582361e-11, 
    2.581617e-11, 2.572562e-11, 2.567999e-11, 2.558445e-11, 2.560179e-11, 
    2.567197e-11, 2.583108e-11, 2.577707e-11, 2.59132e-11, 2.591012e-11, 
    2.606168e-11, 2.599334e-11, 2.624809e-11, 2.617568e-11, 2.638493e-11, 
    2.63323e-11, 2.638245e-11, 2.636725e-11, 2.638265e-11, 2.630547e-11, 
    2.633854e-11, 2.627063e-11, 2.600614e-11, 2.608386e-11, 2.585205e-11, 
    2.571267e-11, 2.562011e-11, 2.555442e-11, 2.556371e-11, 2.558141e-11, 
    2.567238e-11, 2.575792e-11, 2.582311e-11, 2.586671e-11, 2.590968e-11, 
    2.603973e-11, 2.610858e-11, 2.626273e-11, 2.623491e-11, 2.628204e-11, 
    2.632707e-11, 2.640266e-11, 2.639022e-11, 2.642352e-11, 2.62808e-11, 
    2.637565e-11, 2.621907e-11, 2.626189e-11, 2.592134e-11, 2.579164e-11, 
    2.57365e-11, 2.568825e-11, 2.557085e-11, 2.565192e-11, 2.561996e-11, 
    2.5696e-11, 2.574431e-11, 2.572042e-11, 2.586791e-11, 2.581057e-11, 
    2.611266e-11, 2.598253e-11, 2.632181e-11, 2.624062e-11, 2.634128e-11, 
    2.628991e-11, 2.637792e-11, 2.629872e-11, 2.643592e-11, 2.64658e-11, 
    2.644538e-11, 2.652382e-11, 2.629433e-11, 2.638245e-11, 2.571975e-11, 
    2.572365e-11, 2.57418e-11, 2.566199e-11, 2.56571e-11, 2.558397e-11, 
    2.564905e-11, 2.567676e-11, 2.574712e-11, 2.578873e-11, 2.582829e-11, 
    2.591527e-11, 2.601242e-11, 2.614827e-11, 2.624589e-11, 2.631132e-11, 
    2.62712e-11, 2.630662e-11, 2.626702e-11, 2.624846e-11, 2.645461e-11, 
    2.633885e-11, 2.651254e-11, 2.650293e-11, 2.642431e-11, 2.650401e-11, 
    2.572638e-11, 2.570396e-11, 2.562609e-11, 2.568703e-11, 2.557601e-11, 
    2.563815e-11, 2.567388e-11, 2.581176e-11, 2.584206e-11, 2.587015e-11, 
    2.592563e-11, 2.599684e-11, 2.612176e-11, 2.623045e-11, 2.632969e-11, 
    2.632242e-11, 2.632498e-11, 2.634714e-11, 2.629223e-11, 2.635616e-11, 
    2.636688e-11, 2.633884e-11, 2.650164e-11, 2.645513e-11, 2.650272e-11, 
    2.647244e-11, 2.571125e-11, 2.574898e-11, 2.572859e-11, 2.576694e-11, 
    2.573992e-11, 2.586004e-11, 2.589606e-11, 2.60646e-11, 2.599544e-11, 
    2.610552e-11, 2.600662e-11, 2.602414e-11, 2.610911e-11, 2.601197e-11, 
    2.622445e-11, 2.608039e-11, 2.6348e-11, 2.620412e-11, 2.635702e-11, 
    2.632926e-11, 2.637523e-11, 2.64164e-11, 2.64682e-11, 2.656377e-11, 
    2.654164e-11, 2.662157e-11, 2.580524e-11, 2.585419e-11, 2.584988e-11, 
    2.590111e-11, 2.5939e-11, 2.602112e-11, 2.615283e-11, 2.61033e-11, 
    2.619423e-11, 2.621248e-11, 2.607434e-11, 2.615915e-11, 2.588695e-11, 
    2.593092e-11, 2.590475e-11, 2.58091e-11, 2.611471e-11, 2.595786e-11, 
    2.62475e-11, 2.616253e-11, 2.641052e-11, 2.628718e-11, 2.652946e-11, 
    2.663302e-11, 2.673051e-11, 2.684442e-11, 2.588091e-11, 2.584765e-11, 
    2.59072e-11, 2.59896e-11, 2.606606e-11, 2.616771e-11, 2.617811e-11, 
    2.619715e-11, 2.624648e-11, 2.628796e-11, 2.620317e-11, 2.629836e-11, 
    2.594111e-11, 2.612832e-11, 2.583507e-11, 2.592337e-11, 2.598474e-11, 
    2.595782e-11, 2.609764e-11, 2.613059e-11, 2.62645e-11, 2.619528e-11, 
    2.660745e-11, 2.642509e-11, 2.693117e-11, 2.678973e-11, 2.583603e-11, 
    2.588079e-11, 2.60366e-11, 2.596247e-11, 2.617449e-11, 2.622669e-11, 
    2.626912e-11, 2.632335e-11, 2.632921e-11, 2.636135e-11, 2.630869e-11, 
    2.635927e-11, 2.616792e-11, 2.625343e-11, 2.60188e-11, 2.60759e-11, 
    2.604963e-11, 2.602082e-11, 2.610975e-11, 2.62045e-11, 2.620653e-11, 
    2.623692e-11, 2.632252e-11, 2.617536e-11, 2.663098e-11, 2.634958e-11, 
    2.592961e-11, 2.601584e-11, 2.602816e-11, 2.599476e-11, 2.622145e-11, 
    2.613931e-11, 2.636056e-11, 2.630077e-11, 2.639875e-11, 2.635006e-11, 
    2.634289e-11, 2.628036e-11, 2.624143e-11, 2.614308e-11, 2.606305e-11, 
    2.59996e-11, 2.601436e-11, 2.608406e-11, 2.62103e-11, 2.632974e-11, 
    2.630358e-11, 2.63913e-11, 2.615912e-11, 2.625647e-11, 2.621884e-11, 
    2.631696e-11, 2.610198e-11, 2.628503e-11, 2.605519e-11, 2.607534e-11, 
    2.613768e-11, 2.626307e-11, 2.629082e-11, 2.632044e-11, 2.630217e-11, 
    2.621351e-11, 2.619898e-11, 2.613617e-11, 2.611882e-11, 2.607096e-11, 
    2.603133e-11, 2.606753e-11, 2.610556e-11, 2.621355e-11, 2.631087e-11, 
    2.641698e-11, 2.644295e-11, 2.656693e-11, 2.6466e-11, 2.663255e-11, 
    2.649094e-11, 2.673608e-11, 2.629565e-11, 2.648679e-11, 2.614052e-11, 
    2.617782e-11, 2.624529e-11, 2.640004e-11, 2.63165e-11, 2.641421e-11, 
    2.619841e-11, 2.608646e-11, 2.60575e-11, 2.600346e-11, 2.605874e-11, 
    2.605424e-11, 2.610713e-11, 2.609014e-11, 2.621713e-11, 2.614891e-11, 
    2.634271e-11, 2.641344e-11, 2.661319e-11, 2.673564e-11, 2.68603e-11, 
    2.691534e-11, 2.693209e-11, 2.69391e-11 ;

 SOIL3C_vr =
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  7.709882e-21, -5.139921e-21, -2.569961e-21, 0, 1.28498e-20, -1.541976e-20, 
    1.027984e-20, 1.541976e-20, -2.569961e-21, 1.28498e-20, -2.569961e-21, 
    -1.541976e-20, 2.569961e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 
    -1.027984e-20, -7.709882e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    7.709882e-21, -7.709882e-21, -5.139921e-21, -1.541976e-20, -5.139921e-21, 
    2.569961e-21, 5.139921e-21, -1.28498e-20, -7.709882e-21, -7.709882e-21, 
    -2.569961e-21, -7.709882e-21, 1.541976e-20, 5.139921e-21, 7.709882e-21, 
    -5.139921e-21, 0, -5.139921e-21, -1.003089e-36, -1.541976e-20, 
    -1.798972e-20, -1.798972e-20, 0, -1.798972e-20, 2.055969e-20, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, -1.28498e-20, 7.709882e-21, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, 0, -1.798972e-20, 5.139921e-21, 
    1.541976e-20, -1.027984e-20, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    1.541976e-20, 7.709882e-21, 1.027984e-20, -1.541976e-20, 2.569961e-21, 0, 
    0, 2.569961e-21, -7.709882e-21, 1.003089e-36, 2.569961e-21, -1.28498e-20, 
    1.28498e-20, -2.055969e-20, 1.541976e-20, 7.709882e-21, -7.709882e-21, 
    5.139921e-21, -7.709882e-21, 7.709882e-21, 1.541976e-20, 7.709882e-21, 
    1.027984e-20, 1.027984e-20, 0, -2.569961e-21, -2.569961e-21, 
    1.541976e-20, -5.139921e-21, 5.139921e-21, 1.003089e-36, -1.28498e-20, 0, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 1.003089e-36, -1.003089e-36, 
    -1.027984e-20, 5.139921e-21, -1.003089e-36, 1.003089e-36, -1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 1.003089e-36, 1.027984e-20, 
    -5.139921e-21, 0, -1.027984e-20, -1.28498e-20, -5.139921e-21, 
    7.709882e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, 
    1.027984e-20, -1.28498e-20, -1.28498e-20, 2.569961e-21, 1.798972e-20, 
    2.569961e-21, 1.541976e-20, -1.003089e-36, 5.139921e-21, 1.027984e-20, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, -2.055969e-20, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    -2.569961e-21, 1.027984e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, 5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -1.003089e-36, 2.569961e-21, -2.569961e-21, 1.798972e-20, 
    1.541976e-20, 2.312965e-20, 2.569961e-21, -1.003089e-36, -1.003089e-36, 
    5.139921e-21, 7.709882e-21, 2.055969e-20, 2.569961e-21, -2.569961e-21, 
    1.28498e-20, 1.798972e-20, 5.139921e-21, -3.083953e-20, 7.709882e-21, 
    -1.541976e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, -1.798972e-20, 
    5.139921e-21, -5.139921e-21, -2.055969e-20, 7.709882e-21, 7.709882e-21, 
    -1.28498e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -1.28498e-20, -1.003089e-36, 0, 2.055969e-20, -5.139921e-21, 
    5.139921e-21, 1.003089e-36, -1.027984e-20, 0, -1.003089e-36, 
    2.569961e-21, 0, -1.003089e-36, -1.003089e-36, 5.139921e-21, 
    5.139921e-21, 1.003089e-36, 1.541976e-20, -1.28498e-20, -1.027984e-20, 
    7.709882e-21, 1.798972e-20, -1.027984e-20, -2.569961e-21, -1.28498e-20, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, -7.709882e-21, -1.027984e-20, 
    7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, -1.541976e-20, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, 1.28498e-20, 1.28498e-20, 
    1.541976e-20, -7.709882e-21, -1.28498e-20, 5.139921e-21, 7.709882e-21, 
    -1.027984e-20, 2.569961e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -1.28498e-20, -7.709882e-21, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, -1.28498e-20, -1.28498e-20, -1.28498e-20, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, -7.709882e-21, 2.055969e-20, 
    1.003089e-36, 5.139921e-21, -7.709882e-21, -1.28498e-20, 1.28498e-20, 
    7.709882e-21, -5.139921e-21, -7.709882e-21, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 
    1.027984e-20, 1.28498e-20, 7.709882e-21, 7.709882e-21, -2.569961e-21, 
    1.027984e-20, -5.139921e-21, 1.003089e-36, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, -1.541976e-20, 2.569961e-21, 
    -7.709882e-21, 1.003089e-36, 7.709882e-21, 1.28498e-20, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, -2.569961e-20, -7.709882e-21, 1.003089e-36, 
    1.027984e-20, 1.027984e-20, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -1.28498e-20, -7.709882e-21, -7.709882e-21, 
    -1.003089e-36, 5.139921e-21, -2.569961e-21, -1.027984e-20, 1.027984e-20, 
    -1.027984e-20, -1.28498e-20, 2.569961e-21, -1.798972e-20, -2.569961e-21, 
    2.312965e-20, -5.139921e-21, -7.709882e-21, 1.541976e-20, -1.541976e-20, 
    1.027984e-20, -1.798972e-20, -2.569961e-21, -1.798972e-20, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 0, 
    -1.027984e-20, 2.569961e-21, -1.027984e-20, 5.139921e-21,
  1.28498e-20, -5.139921e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, -5.139921e-21, -1.003089e-36, 2.569961e-21, 5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, 2.569961e-21, 1.027984e-20, 
    7.709882e-21, 7.709882e-21, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    2.569961e-21, 2.569961e-21, 0, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -1.027984e-20, -1.28498e-20, -5.139921e-21, 5.139921e-21, 
    -1.003089e-36, 2.569961e-21, -1.28498e-20, 2.569961e-21, -1.541976e-20, 
    -1.541976e-20, -2.569961e-21, -1.28498e-20, 0, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -1.541976e-20, 7.709882e-21, 5.139921e-21, 
    0, 7.709882e-21, 1.027984e-20, -1.027984e-20, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, 1.541976e-20, -5.139921e-21, 7.709882e-21, 0, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, -7.709882e-21, 
    -1.28498e-20, -5.139921e-21, 5.139921e-21, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, 0, -5.139921e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    7.709882e-21, 1.28498e-20, 7.709882e-21, -1.027984e-20, -1.027984e-20, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, 5.139921e-21, 0, 
    2.569961e-21, 1.541976e-20, -1.027984e-20, 0, -7.709882e-21, 
    5.139921e-21, -1.003089e-36, 1.027984e-20, -1.027984e-20, 1.28498e-20, 
    7.709882e-21, 0, 5.139921e-21, 5.139921e-21, 0, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, 1.28498e-20, 1.027984e-20, 1.003089e-36, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, -2.569961e-21, 7.709882e-21, 
    0, -2.569961e-21, 7.709882e-21, -1.28498e-20, -2.569961e-21, 
    1.027984e-20, -1.003089e-36, -7.709882e-21, -7.709882e-21, -5.139921e-21, 
    -5.139921e-21, 7.709882e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 1.003089e-36, -2.569961e-21, 0, 1.28498e-20, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 0, 5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 0, -7.709882e-21, 1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, -1.28498e-20, 
    1.28498e-20, -5.139921e-21, 1.027984e-20, -2.569961e-21, 0, 1.28498e-20, 
    -1.027984e-20, 0, -1.28498e-20, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, -1.027984e-20, -7.709882e-21, -2.569961e-21, -7.709882e-21, 
    0, -1.003089e-36, -2.569961e-21, 5.139921e-21, 1.28498e-20, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, 
    5.139921e-21, 2.569961e-21, 1.28498e-20, 0, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, -1.027984e-20, 7.709882e-21, 0, 
    -2.569961e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 1.541976e-20, 
    2.569961e-21, -1.28498e-20, -5.139921e-21, -7.709882e-21, -2.569961e-21, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, -1.28498e-20, -7.709882e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 1.003089e-36, 2.569961e-21, 
    1.28498e-20, 1.003089e-36, -1.28498e-20, 2.569961e-21, 5.139921e-21, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, -7.709882e-21, -1.027984e-20, 
    1.28498e-20, 2.569961e-21, -7.709882e-21, -7.709882e-21, 1.798972e-20, 
    2.055969e-20, -1.027984e-20, 1.28498e-20, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 1.003089e-36, -7.709882e-21, 1.027984e-20, -5.139921e-21, 
    0, 5.139921e-21, -2.569961e-21, -1.798972e-20, -5.139921e-21, 
    7.709882e-21, 0, -1.027984e-20, 7.709882e-21, 1.28498e-20, 1.027984e-20, 
    1.027984e-20, 1.28498e-20, -2.569961e-21, 1.003089e-36, -7.709882e-21, 
    5.139921e-21, 1.027984e-20, -2.569961e-21, -7.709882e-21, 5.139921e-21, 
    1.541976e-20, 1.798972e-20, -2.569961e-21, -7.709882e-21, 5.139921e-21, 
    0, 0, -1.28498e-20, 1.28498e-20, 5.139921e-21, 2.569961e-21, 
    -1.003089e-36, -2.569961e-21, -1.027984e-20, -1.28498e-20, -2.569961e-21, 
    -5.139921e-21, 1.541976e-20, 2.569961e-21, 0, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 2.569961e-21, -1.28498e-20, 0, 
    5.139921e-21, 5.139921e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -1.541976e-20, -5.139921e-21, 0, -1.003089e-36, -7.709882e-21, 
    5.139921e-21, 2.569961e-21, 0, 0, 7.709882e-21, -5.139921e-21, 
    1.541976e-20, 2.569961e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, 0, -1.28498e-20, -7.709882e-21, -1.027984e-20, 
    2.569961e-21, 5.139921e-21, -1.28498e-20, 0, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -7.709882e-21, -1.027984e-20, 0, -1.798972e-20, 
    5.139921e-21, 2.569961e-21,
  -2.569961e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, -1.027984e-20, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    2.569961e-21, 7.709882e-21, -7.709882e-21, 1.027984e-20, -2.569961e-21, 
    2.569961e-21, 5.139921e-21, 1.541976e-20, 0, 5.139921e-21, 5.139921e-21, 
    -1.28498e-20, 0, -2.569961e-21, 2.569961e-21, 2.569961e-21, 1.027984e-20, 
    1.003089e-36, -7.709882e-21, 1.027984e-20, -1.28498e-20, 1.28498e-20, 0, 
    2.569961e-21, -5.139921e-21, 1.541976e-20, -7.709882e-21, -2.312965e-20, 
    1.798972e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, 0, 
    -2.569961e-21, -7.709882e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, 1.003089e-36, -2.569961e-21, 
    0, 2.569961e-21, 7.709882e-21, -2.569961e-21, 5.139921e-21, 1.798972e-20, 
    -2.312965e-20, 1.027984e-20, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 0, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, 0, 5.139921e-21, -1.541976e-20, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, -1.003089e-36, 2.569961e-20, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    7.709882e-21, -1.28498e-20, -1.541976e-20, 2.569961e-21, 0, 
    -1.027984e-20, -1.003089e-36, -1.003089e-36, 2.569961e-21, 1.28498e-20, 
    0, -2.569961e-21, -1.027984e-20, 5.139921e-21, -1.28498e-20, 1.28498e-20, 
    1.027984e-20, -5.139921e-21, 0, 1.798972e-20, 7.709882e-21, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, -1.28498e-20, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, 5.139921e-21, 1.003089e-36, -2.569961e-21, 
    2.569961e-21, -5.139921e-21, 1.027984e-20, -5.139921e-21, 0, 
    5.139921e-21, -7.709882e-21, 7.709882e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, -1.541976e-20, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 
    5.139921e-21, 0, 5.139921e-21, -1.027984e-20, 0, -1.28498e-20, 
    7.709882e-21, 2.569961e-21, 0, -2.569961e-21, -1.28498e-20, 1.027984e-20, 
    2.569961e-21, 5.139921e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, -1.541976e-20, -1.798972e-20, -2.569961e-21, -5.139921e-21, 
    1.027984e-20, 2.569961e-21, 1.28498e-20, 0, 1.28498e-20, 1.541976e-20, 
    -2.569961e-21, 0, -7.709882e-21, -7.709882e-21, 7.709882e-21, 
    -1.28498e-20, -5.139921e-21, -1.027984e-20, 1.541976e-20, -1.28498e-20, 
    -5.139921e-21, 1.28498e-20, -1.541976e-20, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -1.28498e-20, -1.28498e-20, 7.709882e-21, 7.709882e-21, 
    -7.709882e-21, -1.027984e-20, 1.541976e-20, 1.027984e-20, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, 0, -1.28498e-20, 1.28498e-20, 
    -7.709882e-21, 2.569961e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    1.027984e-20, -1.027984e-20, 5.139921e-21, 1.798972e-20, 7.709882e-21, 
    -5.139921e-21, 1.28498e-20, -1.027984e-20, 1.28498e-20, 0, -7.709882e-21, 
    -1.003089e-36, -1.027984e-20, -1.003089e-36, 0, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 1.541976e-20, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, -1.027984e-20, 2.569961e-21, 
    -7.709882e-21, -7.709882e-21, 5.139921e-21, -1.541976e-20, 1.541976e-20, 
    1.027984e-20, -2.569961e-21, 2.569961e-21, -1.003089e-36, -7.709882e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, 1.027984e-20, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, 0, 0, 0, 5.139921e-21, 
    -1.798972e-20, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.003089e-36, 1.28498e-20, 0, 5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 1.28498e-20, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, 1.027984e-20, -1.003089e-36, 
    -1.027984e-20, 2.569961e-21, 0, -2.569961e-21, 1.027984e-20, 
    -1.003089e-36, 7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 1.027984e-20, 
    -2.569961e-21, -1.027984e-20, -7.709882e-21, -2.569961e-20, 2.569961e-21, 
    5.139921e-21, -1.003089e-36, -1.003089e-36, -1.003089e-36, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -1.28498e-20, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, 1.003089e-36, 1.003089e-36, 
    5.139921e-21, -5.139921e-21, 1.28498e-20, -7.709882e-21, 0, 2.569961e-21, 
    -2.569961e-21, -1.003089e-36, -1.027984e-20, 0, -2.569961e-21, 
    -1.003089e-36, -5.139921e-21, 7.709882e-21, 1.027984e-20, 1.027984e-20, 
    -2.826957e-20, -2.055969e-20, 1.003089e-36, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, -1.798972e-20, 7.709882e-21, 
    1.027984e-20, 7.709882e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 
    7.709882e-21,
  2.569961e-21, -2.569961e-20, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, 5.139921e-21, 1.027984e-20, 1.798972e-20, 0, -1.003089e-36, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, -1.28498e-20, -2.569961e-21, 
    2.569961e-21, -5.139921e-21, -2.569961e-21, 1.027984e-20, -1.28498e-20, 
    1.28498e-20, 2.569961e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    7.709882e-21, 2.569961e-21, 1.003089e-36, -7.709882e-21, 2.569961e-21, 
    -1.027984e-20, 2.312965e-20, 1.28498e-20, 1.28498e-20, 0, 2.569961e-21, 
    1.28498e-20, -2.569961e-21, -1.003089e-36, -5.139921e-21, -1.027984e-20, 
    1.798972e-20, -2.569961e-20, 7.709882e-21, 2.569961e-21, 7.709882e-21, 
    -5.139921e-21, 1.003089e-36, -5.139921e-21, 7.709882e-21, 5.139921e-21, 
    1.003089e-36, 0, -1.027984e-20, 1.541976e-20, 7.709882e-21, 5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, -7.709882e-21, 
    2.312965e-20, -1.28498e-20, -2.569961e-21, 7.709882e-21, 7.709882e-21, 
    1.027984e-20, -5.139921e-21, -1.28498e-20, -2.569961e-21, -1.541976e-20, 
    1.027984e-20, 0, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -1.541976e-20, -7.709882e-21, -1.28498e-20, -1.541976e-20, 1.541976e-20, 
    -2.312965e-20, 0, 1.28498e-20, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, -1.798972e-20, -7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    7.709882e-21, 1.28498e-20, 5.139921e-21, -1.28498e-20, 1.28498e-20, 
    7.709882e-21, 2.055969e-20, 5.139921e-21, 2.569961e-21, -7.709882e-21, 
    1.28498e-20, -1.28498e-20, 5.139921e-21, 1.28498e-20, 1.541976e-20, 
    1.027984e-20, -7.709882e-21, 7.709882e-21, -1.541976e-20, -5.139921e-21, 
    2.569961e-21, 0, -7.709882e-21, 1.027984e-20, 7.709882e-21, 1.541976e-20, 
    -5.139921e-21, 7.709882e-21, 0, -7.709882e-21, -1.541976e-20, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, -2.569961e-21, 5.139921e-21, -1.027984e-20, 7.709882e-21, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    1.027984e-20, 2.055969e-20, 1.027984e-20, 5.139921e-21, 1.003089e-36, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 1.541976e-20, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, -1.798972e-20, 2.569961e-21, 1.027984e-20, 2.312965e-20, 
    1.28498e-20, -2.569961e-21, -2.569961e-21, -1.798972e-20, -2.569961e-21, 
    1.28498e-20, -2.569961e-20, 2.569961e-21, 2.055969e-20, -2.569961e-21, 
    1.798972e-20, -5.139921e-21, -2.569961e-21, 7.709882e-21, 1.28498e-20, 0, 
    -2.055969e-20, 7.709882e-21, -5.139921e-21, -1.798972e-20, -7.709882e-21, 
    2.569961e-21, 2.569961e-21, -2.569961e-21, 1.28498e-20, -7.709882e-21, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, 1.541976e-20, -5.139921e-21, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, 7.709882e-21, 1.003089e-36, 
    -7.709882e-21, 5.139921e-21, -2.312965e-20, 1.003089e-36, -7.709882e-21, 
    1.003089e-36, 7.709882e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, -7.709882e-21, 0, 
    -5.139921e-21, -1.541976e-20, 2.569961e-21, 7.709882e-21, 0, 
    -5.139921e-21, -2.569961e-21, 1.027984e-20, -2.055969e-20, 1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 1.28498e-20, -5.139921e-21, 1.28498e-20, 
    2.569961e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    -1.003089e-36, 1.027984e-20, -5.139921e-21, -1.541976e-20, -1.541976e-20, 
    -2.569961e-21, -1.798972e-20, 7.709882e-21, -5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, -1.003089e-36, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    1.027984e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    1.027984e-20, 1.28498e-20, -1.28498e-20, -5.139921e-21, -5.139921e-21, 
    -1.28498e-20, -1.28498e-20, -1.027984e-20, 2.569961e-21, -1.28498e-20, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, -1.798972e-20, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 1.28498e-20, 
    -7.709882e-21, -1.003089e-36, 1.541976e-20, 7.709882e-21, -7.709882e-21, 
    -5.139921e-21, -1.027984e-20, -1.541976e-20, -1.798972e-20, 0, 
    -1.003089e-36, 2.569961e-21, 2.569961e-21, -7.709882e-21, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, -7.709882e-21, -7.709882e-21, 
    2.312965e-20, -1.28498e-20, -2.312965e-20, -5.139921e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    1.003089e-36, -7.709882e-21, 2.055969e-20, -2.569961e-21, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 
    0, 5.139921e-21, -1.28498e-20,
  -1.003089e-36, -1.798972e-20, 1.28498e-20, -7.709882e-21, 5.139921e-21, 
    -1.28498e-20, 2.569961e-21, 1.003089e-36, -2.569961e-21, 1.003089e-36, 
    1.027984e-20, 7.709882e-21, -7.709882e-21, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, 1.541976e-20, -5.139921e-21, 1.28498e-20, -2.569961e-21, 
    5.139921e-21, 1.541976e-20, 2.055969e-20, -1.027984e-20, -1.027984e-20, 
    -1.541976e-20, -1.003089e-36, -1.027984e-20, 5.139921e-21, -7.709882e-21, 
    -1.027984e-20, -2.055969e-20, 7.709882e-21, -7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, 7.709882e-21, -1.027984e-20, -2.569961e-21, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, -1.541976e-20, -5.139921e-21, 
    1.003089e-36, 5.139921e-21, 5.139921e-21, -2.055969e-20, -1.28498e-20, 
    -5.139921e-21, -1.027984e-20, 1.027984e-20, 1.541976e-20, -5.139921e-21, 
    7.709882e-21, -1.541976e-20, -2.312965e-20, 0, -2.569961e-21, 
    -5.139921e-21, -1.28498e-20, -1.003089e-36, 7.709882e-21, -2.569961e-21, 
    1.027984e-20, 7.709882e-21, 2.312965e-20, -1.28498e-20, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, -1.798972e-20, -1.541976e-20, 
    5.139921e-21, 2.055969e-20, 2.569961e-21, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, 5.139921e-21, -1.798972e-20, -1.027984e-20, 5.139921e-21, 
    7.709882e-21, -7.709882e-21, -1.027984e-20, -5.139921e-21, -7.709882e-21, 
    -1.28498e-20, 1.28498e-20, 5.139921e-21, -1.541976e-20, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 1.541976e-20, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, 5.139921e-21, 1.28498e-20, 0, -2.569961e-21, 7.709882e-21, 
    -1.798972e-20, 1.541976e-20, 7.709882e-21, 1.28498e-20, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, -7.709882e-21, -1.027984e-20, 
    2.569961e-21, 1.28498e-20, 1.798972e-20, 2.569961e-21, -1.027984e-20, 0, 
    7.709882e-21, 1.027984e-20, 1.798972e-20, 2.569961e-21, -7.709882e-21, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 
    7.709882e-21, -1.28498e-20, 7.709882e-21, 1.541976e-20, 5.139921e-21, 
    -2.312965e-20, -1.541976e-20, 1.003089e-36, 1.28498e-20, 1.28498e-20, 
    -2.826957e-20, -1.798972e-20, -1.027984e-20, 7.709882e-21, -2.569961e-21, 
    5.139921e-21, 1.027984e-20, -1.798972e-20, 2.569961e-21, -2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 1.28498e-20, 7.709882e-21, -1.027984e-20, 
    -2.569961e-21, 1.027984e-20, -1.027984e-20, 1.027984e-20, -2.569961e-21, 
    -1.798972e-20, 5.139921e-21, 1.027984e-20, 1.28498e-20, 1.28498e-20, 
    7.709882e-21, 5.139921e-21, -1.28498e-20, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, -1.28498e-20, 2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, -1.027984e-20, -1.541976e-20, 
    -7.709882e-21, 2.569961e-21, -1.28498e-20, 1.28498e-20, -1.798972e-20, 
    7.709882e-21, -1.003089e-36, 1.003089e-36, -1.798972e-20, 1.798972e-20, 
    2.569961e-21, 1.003089e-36, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -2.569961e-21, -2.569961e-20, 2.055969e-20, 1.28498e-20, 7.709882e-21, 
    -2.055969e-20, -5.139921e-21, 1.28498e-20, -7.709882e-21, 1.798972e-20, 
    1.504633e-36, -1.798972e-20, -1.027984e-20, -5.139921e-21, 0, 
    -1.798972e-20, 1.027984e-20, -5.139921e-21, -2.569961e-21, -1.027984e-20, 
    0, -2.569961e-21, 1.28498e-20, 1.003089e-36, -5.139921e-21, 5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -1.28498e-20, -2.055969e-20, -5.139921e-21, 
    5.139921e-21, 1.541976e-20, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -1.541976e-20, -1.027984e-20, -1.798972e-20, 2.569961e-21, -2.569961e-21, 
    1.28498e-20, -1.027984e-20, -2.569961e-21, 5.139921e-21, 2.569961e-20, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 2.312965e-20, 
    -7.709882e-21, -2.312965e-20, -1.027984e-20, 7.709882e-21, 2.569961e-21, 
    -1.003089e-36, 1.027984e-20, -1.28498e-20, -1.28498e-20, -5.139921e-21, 
    7.709882e-21, -5.139921e-21, -2.569961e-21, -1.027984e-20, -5.139921e-21, 
    -2.569961e-21, 1.798972e-20, -1.541976e-20, -7.709882e-21, 1.027984e-20, 
    -7.709882e-21, -2.569961e-21, 7.709882e-21, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, 7.709882e-21, -7.709882e-21, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -1.003089e-36, 1.003089e-36, 1.003089e-36, 7.709882e-21, 
    2.569961e-21, -7.709882e-21, -1.541976e-20, -1.027984e-20, 5.139921e-21, 
    2.569961e-21, 1.003089e-36, 5.139921e-21, -2.569961e-21, 1.28498e-20, 
    1.28498e-20, -2.569961e-21, -5.139921e-21, 1.28498e-20, -2.569961e-21, 
    1.798972e-20, 1.541976e-20, 1.027984e-20, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, -1.28498e-20, -1.003089e-36, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -1.798972e-20, 2.569961e-21, -7.709882e-21, 
    1.027984e-20, -1.003089e-36, -7.709882e-21, 2.569961e-21, -1.003089e-36, 
    -7.709882e-21, 1.027984e-20, 2.312965e-20, -1.28498e-20, 2.569961e-21, 
    5.139921e-21, -1.027984e-20, 2.569961e-21, -1.28498e-20, 1.027984e-20, 
    -7.709882e-21, 2.569961e-21, 7.709882e-21, 1.027984e-20, 7.709882e-21, 
    1.28498e-20, -2.826957e-20, 1.541976e-20, -2.569961e-21, -1.28498e-20,
  6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.170318e-12, 5.193127e-12, 5.188693e-12, 5.20709e-12, 5.196885e-12, 
    5.208931e-12, 5.174943e-12, 5.194032e-12, 5.181846e-12, 5.172372e-12, 
    5.242793e-12, 5.207911e-12, 5.279034e-12, 5.256785e-12, 5.31268e-12, 
    5.275571e-12, 5.320164e-12, 5.311611e-12, 5.337356e-12, 5.32998e-12, 
    5.362909e-12, 5.34076e-12, 5.379981e-12, 5.357621e-12, 5.361118e-12, 
    5.340029e-12, 5.214932e-12, 5.238449e-12, 5.213538e-12, 5.216892e-12, 
    5.215387e-12, 5.197095e-12, 5.187877e-12, 5.168575e-12, 5.172079e-12, 
    5.186257e-12, 5.218399e-12, 5.207489e-12, 5.234989e-12, 5.234368e-12, 
    5.264985e-12, 5.25118e-12, 5.302644e-12, 5.288017e-12, 5.330288e-12, 
    5.319657e-12, 5.329789e-12, 5.326716e-12, 5.329829e-12, 5.314237e-12, 
    5.320917e-12, 5.307198e-12, 5.253765e-12, 5.269468e-12, 5.222637e-12, 
    5.194479e-12, 5.17578e-12, 5.16251e-12, 5.164386e-12, 5.167962e-12, 
    5.18634e-12, 5.20362e-12, 5.21679e-12, 5.225599e-12, 5.234279e-12, 
    5.260551e-12, 5.27446e-12, 5.305601e-12, 5.299982e-12, 5.309502e-12, 
    5.318599e-12, 5.333871e-12, 5.331357e-12, 5.338085e-12, 5.309252e-12, 
    5.328414e-12, 5.296781e-12, 5.305433e-12, 5.236634e-12, 5.210433e-12, 
    5.199293e-12, 5.189545e-12, 5.165828e-12, 5.182206e-12, 5.17575e-12, 
    5.191111e-12, 5.200872e-12, 5.196045e-12, 5.22584e-12, 5.214256e-12, 
    5.275284e-12, 5.248996e-12, 5.317538e-12, 5.301136e-12, 5.32147e-12, 
    5.311094e-12, 5.328872e-12, 5.312872e-12, 5.34059e-12, 5.346627e-12, 
    5.342501e-12, 5.358347e-12, 5.311985e-12, 5.329788e-12, 5.195909e-12, 
    5.196696e-12, 5.200364e-12, 5.18424e-12, 5.183254e-12, 5.168479e-12, 
    5.181626e-12, 5.187224e-12, 5.201438e-12, 5.209845e-12, 5.217837e-12, 
    5.235409e-12, 5.255034e-12, 5.28248e-12, 5.302199e-12, 5.315417e-12, 
    5.307312e-12, 5.314468e-12, 5.306469e-12, 5.30272e-12, 5.344365e-12, 
    5.320979e-12, 5.356068e-12, 5.354127e-12, 5.338245e-12, 5.354345e-12, 
    5.197249e-12, 5.192719e-12, 5.176988e-12, 5.189299e-12, 5.16687e-12, 
    5.179424e-12, 5.186642e-12, 5.214497e-12, 5.220618e-12, 5.226293e-12, 
    5.237502e-12, 5.251887e-12, 5.277122e-12, 5.299081e-12, 5.319129e-12, 
    5.31766e-12, 5.318177e-12, 5.322655e-12, 5.311562e-12, 5.324476e-12, 
    5.326643e-12, 5.320977e-12, 5.353867e-12, 5.344471e-12, 5.354085e-12, 
    5.347968e-12, 5.194191e-12, 5.201815e-12, 5.197695e-12, 5.205442e-12, 
    5.199984e-12, 5.224251e-12, 5.231527e-12, 5.265577e-12, 5.251603e-12, 
    5.273843e-12, 5.253863e-12, 5.257403e-12, 5.274567e-12, 5.254943e-12, 
    5.29787e-12, 5.268765e-12, 5.322829e-12, 5.293762e-12, 5.32465e-12, 
    5.319042e-12, 5.328328e-12, 5.336645e-12, 5.347111e-12, 5.366418e-12, 
    5.361947e-12, 5.378094e-12, 5.213181e-12, 5.223069e-12, 5.222199e-12, 
    5.232547e-12, 5.240201e-12, 5.256791e-12, 5.283399e-12, 5.273394e-12, 
    5.291764e-12, 5.295451e-12, 5.267543e-12, 5.284677e-12, 5.229687e-12, 
    5.23857e-12, 5.233282e-12, 5.21396e-12, 5.275698e-12, 5.244013e-12, 
    5.302525e-12, 5.285359e-12, 5.33546e-12, 5.310542e-12, 5.359486e-12, 
    5.380408e-12, 5.400103e-12, 5.423116e-12, 5.228466e-12, 5.221747e-12, 
    5.233779e-12, 5.250423e-12, 5.26587e-12, 5.286405e-12, 5.288507e-12, 
    5.292354e-12, 5.30232e-12, 5.310698e-12, 5.293569e-12, 5.312799e-12, 
    5.240629e-12, 5.278449e-12, 5.219207e-12, 5.237044e-12, 5.249443e-12, 
    5.244004e-12, 5.27225e-12, 5.278908e-12, 5.305961e-12, 5.291976e-12, 
    5.375243e-12, 5.338401e-12, 5.440641e-12, 5.412067e-12, 5.2194e-12, 
    5.228444e-12, 5.25992e-12, 5.244943e-12, 5.287777e-12, 5.29832e-12, 
    5.306893e-12, 5.317849e-12, 5.319033e-12, 5.325525e-12, 5.314887e-12, 
    5.325105e-12, 5.286449e-12, 5.303723e-12, 5.256323e-12, 5.267859e-12, 
    5.262552e-12, 5.25673e-12, 5.274698e-12, 5.293839e-12, 5.294249e-12, 
    5.300387e-12, 5.317681e-12, 5.28795e-12, 5.379996e-12, 5.323146e-12, 
    5.238305e-12, 5.255725e-12, 5.258214e-12, 5.251466e-12, 5.297263e-12, 
    5.280669e-12, 5.325366e-12, 5.313286e-12, 5.33308e-12, 5.323244e-12, 
    5.321797e-12, 5.309164e-12, 5.301299e-12, 5.281429e-12, 5.265263e-12, 
    5.252445e-12, 5.255426e-12, 5.269506e-12, 5.29501e-12, 5.319139e-12, 
    5.313854e-12, 5.331576e-12, 5.284671e-12, 5.304338e-12, 5.296736e-12, 
    5.316558e-12, 5.273127e-12, 5.310107e-12, 5.263675e-12, 5.267746e-12, 
    5.28034e-12, 5.305671e-12, 5.311277e-12, 5.317261e-12, 5.313569e-12, 
    5.295658e-12, 5.292724e-12, 5.280033e-12, 5.276529e-12, 5.26686e-12, 
    5.258855e-12, 5.266169e-12, 5.273849e-12, 5.295666e-12, 5.315327e-12, 
    5.336764e-12, 5.34201e-12, 5.367057e-12, 5.346668e-12, 5.380313e-12, 
    5.351706e-12, 5.401228e-12, 5.312252e-12, 5.350866e-12, 5.280913e-12, 
    5.288448e-12, 5.302078e-12, 5.333342e-12, 5.316465e-12, 5.336203e-12, 
    5.292609e-12, 5.269991e-12, 5.264141e-12, 5.253224e-12, 5.264391e-12, 
    5.263483e-12, 5.274168e-12, 5.270734e-12, 5.29639e-12, 5.282609e-12, 
    5.32176e-12, 5.336048e-12, 5.376402e-12, 5.401139e-12, 5.426324e-12, 
    5.437443e-12, 5.440827e-12, 5.442242e-12 ;

 SOIL3N_vr =
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818189, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818189, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818188, 1.818189, 1.818188, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818189, 1.818188, 1.818189, 1.818188, 1.818188, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 1.818189, 
    1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 
    1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.128042e-11, 3.141842e-11, 3.139159e-11, 3.150289e-11, 3.144116e-11, 
    3.151403e-11, 3.13084e-11, 3.142389e-11, 3.135017e-11, 3.129285e-11, 
    3.171889e-11, 3.150786e-11, 3.193816e-11, 3.180355e-11, 3.214172e-11, 
    3.191721e-11, 3.218699e-11, 3.213525e-11, 3.2291e-11, 3.224638e-11, 
    3.24456e-11, 3.23116e-11, 3.254888e-11, 3.241361e-11, 3.243476e-11, 
    3.230717e-11, 3.155034e-11, 3.169262e-11, 3.15419e-11, 3.156219e-11, 
    3.155309e-11, 3.144243e-11, 3.138666e-11, 3.126988e-11, 3.129108e-11, 
    3.137685e-11, 3.157132e-11, 3.150531e-11, 3.167169e-11, 3.166793e-11, 
    3.185316e-11, 3.176964e-11, 3.2081e-11, 3.19925e-11, 3.224824e-11, 
    3.218393e-11, 3.224522e-11, 3.222663e-11, 3.224546e-11, 3.215113e-11, 
    3.219155e-11, 3.210854e-11, 3.178528e-11, 3.188028e-11, 3.159695e-11, 
    3.142659e-11, 3.131347e-11, 3.123318e-11, 3.124453e-11, 3.126617e-11, 
    3.137736e-11, 3.14819e-11, 3.156158e-11, 3.161487e-11, 3.166739e-11, 
    3.182633e-11, 3.191048e-11, 3.209889e-11, 3.206489e-11, 3.212249e-11, 
    3.217752e-11, 3.226992e-11, 3.225471e-11, 3.229542e-11, 3.212098e-11, 
    3.223691e-11, 3.204553e-11, 3.209787e-11, 3.168164e-11, 3.152312e-11, 
    3.145572e-11, 3.139675e-11, 3.125326e-11, 3.135235e-11, 3.131329e-11, 
    3.140622e-11, 3.146527e-11, 3.143607e-11, 3.161633e-11, 3.154625e-11, 
    3.191547e-11, 3.175643e-11, 3.217111e-11, 3.207187e-11, 3.219489e-11, 
    3.213212e-11, 3.223968e-11, 3.214288e-11, 3.231057e-11, 3.234709e-11, 
    3.232213e-11, 3.2418e-11, 3.213751e-11, 3.224522e-11, 3.143525e-11, 
    3.144001e-11, 3.14622e-11, 3.136465e-11, 3.135868e-11, 3.12693e-11, 
    3.134884e-11, 3.138271e-11, 3.14687e-11, 3.151956e-11, 3.156791e-11, 
    3.167422e-11, 3.179296e-11, 3.1959e-11, 3.207831e-11, 3.215828e-11, 
    3.210924e-11, 3.215253e-11, 3.210414e-11, 3.208145e-11, 3.233341e-11, 
    3.219192e-11, 3.240421e-11, 3.239247e-11, 3.229638e-11, 3.239379e-11, 
    3.144336e-11, 3.141595e-11, 3.132078e-11, 3.139525e-11, 3.125956e-11, 
    3.133551e-11, 3.137918e-11, 3.154771e-11, 3.158474e-11, 3.161907e-11, 
    3.168689e-11, 3.177391e-11, 3.192659e-11, 3.205944e-11, 3.218073e-11, 
    3.217184e-11, 3.217497e-11, 3.220206e-11, 3.213495e-11, 3.221308e-11, 
    3.222619e-11, 3.219191e-11, 3.239089e-11, 3.233405e-11, 3.239222e-11, 
    3.235521e-11, 3.142486e-11, 3.147098e-11, 3.144606e-11, 3.149292e-11, 
    3.14599e-11, 3.160672e-11, 3.165074e-11, 3.185674e-11, 3.17722e-11, 
    3.190675e-11, 3.178587e-11, 3.180729e-11, 3.191113e-11, 3.179241e-11, 
    3.205211e-11, 3.187603e-11, 3.220312e-11, 3.202726e-11, 3.221414e-11, 
    3.21802e-11, 3.223639e-11, 3.22867e-11, 3.235002e-11, 3.246683e-11, 
    3.243978e-11, 3.253747e-11, 3.153974e-11, 3.159957e-11, 3.15943e-11, 
    3.165691e-11, 3.170322e-11, 3.180358e-11, 3.196457e-11, 3.190403e-11, 
    3.201517e-11, 3.203748e-11, 3.186864e-11, 3.19723e-11, 3.163961e-11, 
    3.169335e-11, 3.166135e-11, 3.154446e-11, 3.191798e-11, 3.172628e-11, 
    3.208028e-11, 3.197642e-11, 3.227953e-11, 3.212878e-11, 3.242489e-11, 
    3.255147e-11, 3.267062e-11, 3.280985e-11, 3.163222e-11, 3.159157e-11, 
    3.166436e-11, 3.176506e-11, 3.185852e-11, 3.198275e-11, 3.199547e-11, 
    3.201874e-11, 3.207903e-11, 3.212973e-11, 3.20261e-11, 3.214243e-11, 
    3.17058e-11, 3.193461e-11, 3.15762e-11, 3.168411e-11, 3.175913e-11, 
    3.172623e-11, 3.189711e-11, 3.193739e-11, 3.210106e-11, 3.201646e-11, 
    3.252022e-11, 3.229733e-11, 3.291588e-11, 3.274301e-11, 3.157737e-11, 
    3.163208e-11, 3.182251e-11, 3.173191e-11, 3.199105e-11, 3.205484e-11, 
    3.21067e-11, 3.217299e-11, 3.218015e-11, 3.221943e-11, 3.215506e-11, 
    3.221689e-11, 3.198302e-11, 3.208753e-11, 3.180075e-11, 3.187054e-11, 
    3.183844e-11, 3.180322e-11, 3.191192e-11, 3.202772e-11, 3.203021e-11, 
    3.206734e-11, 3.217197e-11, 3.19921e-11, 3.254898e-11, 3.220504e-11, 
    3.169175e-11, 3.179713e-11, 3.18122e-11, 3.177137e-11, 3.204844e-11, 
    3.194804e-11, 3.221847e-11, 3.214538e-11, 3.226514e-11, 3.220563e-11, 
    3.219687e-11, 3.212045e-11, 3.207286e-11, 3.195265e-11, 3.185484e-11, 
    3.177729e-11, 3.179533e-11, 3.188051e-11, 3.203481e-11, 3.218079e-11, 
    3.214881e-11, 3.225603e-11, 3.197226e-11, 3.209124e-11, 3.204525e-11, 
    3.216518e-11, 3.190242e-11, 3.212615e-11, 3.184523e-11, 3.186986e-11, 
    3.194605e-11, 3.209931e-11, 3.213323e-11, 3.216943e-11, 3.214709e-11, 
    3.203873e-11, 3.202098e-11, 3.19442e-11, 3.1923e-11, 3.18645e-11, 
    3.181607e-11, 3.186032e-11, 3.190679e-11, 3.203878e-11, 3.215773e-11, 
    3.228742e-11, 3.231916e-11, 3.247069e-11, 3.234734e-11, 3.255089e-11, 
    3.237782e-11, 3.267743e-11, 3.213912e-11, 3.237274e-11, 3.194952e-11, 
    3.199511e-11, 3.207757e-11, 3.226672e-11, 3.216461e-11, 3.228403e-11, 
    3.202029e-11, 3.188345e-11, 3.184806e-11, 3.178201e-11, 3.184956e-11, 
    3.184407e-11, 3.190872e-11, 3.188794e-11, 3.204316e-11, 3.195979e-11, 
    3.219665e-11, 3.228309e-11, 3.252723e-11, 3.267689e-11, 3.282926e-11, 
    3.289653e-11, 3.2917e-11, 3.292556e-11 ;

 SOILC =
  17.3448, 17.34478, 17.34479, 17.34477, 17.34478, 17.34477, 17.34479, 
    17.34478, 17.34479, 17.3448, 17.34476, 17.34477, 17.34473, 17.34475, 
    17.34471, 17.34474, 17.34471, 17.34472, 17.3447, 17.3447, 17.34468, 
    17.3447, 17.34468, 17.34469, 17.34469, 17.3447, 17.34477, 17.34476, 
    17.34477, 17.34477, 17.34477, 17.34478, 17.34479, 17.3448, 17.3448, 
    17.34479, 17.34477, 17.34477, 17.34476, 17.34476, 17.34474, 17.34475, 
    17.34472, 17.34473, 17.3447, 17.34471, 17.3447, 17.34471, 17.3447, 
    17.34471, 17.34471, 17.34472, 17.34475, 17.34474, 17.34477, 17.34478, 
    17.34479, 17.3448, 17.3448, 17.3448, 17.34479, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34472, 17.34472, 17.34472, 
    17.34471, 17.3447, 17.3447, 17.3447, 17.34472, 17.34471, 17.34472, 
    17.34472, 17.34476, 17.34477, 17.34478, 17.34479, 17.3448, 17.34479, 
    17.34479, 17.34478, 17.34478, 17.34478, 17.34476, 17.34477, 17.34474, 
    17.34475, 17.34471, 17.34472, 17.34471, 17.34472, 17.34471, 17.34471, 
    17.3447, 17.34469, 17.3447, 17.34469, 17.34472, 17.3447, 17.34478, 
    17.34478, 17.34478, 17.34479, 17.34479, 17.3448, 17.34479, 17.34479, 
    17.34478, 17.34477, 17.34477, 17.34476, 17.34475, 17.34473, 17.34472, 
    17.34471, 17.34472, 17.34471, 17.34472, 17.34472, 17.3447, 17.34471, 
    17.34469, 17.34469, 17.3447, 17.34469, 17.34478, 17.34478, 17.34479, 
    17.34479, 17.3448, 17.34479, 17.34479, 17.34477, 17.34477, 17.34476, 
    17.34476, 17.34475, 17.34473, 17.34472, 17.34471, 17.34471, 17.34471, 
    17.34471, 17.34472, 17.34471, 17.34471, 17.34471, 17.34469, 17.3447, 
    17.34469, 17.34469, 17.34478, 17.34478, 17.34478, 17.34478, 17.34478, 
    17.34476, 17.34476, 17.34474, 17.34475, 17.34474, 17.34475, 17.34475, 
    17.34474, 17.34475, 17.34472, 17.34474, 17.34471, 17.34472, 17.34471, 
    17.34471, 17.34471, 17.3447, 17.34469, 17.34468, 17.34469, 17.34468, 
    17.34477, 17.34476, 17.34477, 17.34476, 17.34476, 17.34475, 17.34473, 
    17.34474, 17.34473, 17.34472, 17.34474, 17.34473, 17.34476, 17.34476, 
    17.34476, 17.34477, 17.34474, 17.34475, 17.34472, 17.34473, 17.3447, 
    17.34472, 17.34469, 17.34468, 17.34466, 17.34465, 17.34476, 17.34477, 
    17.34476, 17.34475, 17.34474, 17.34473, 17.34473, 17.34473, 17.34472, 
    17.34472, 17.34472, 17.34471, 17.34476, 17.34473, 17.34477, 17.34476, 
    17.34475, 17.34475, 17.34474, 17.34473, 17.34472, 17.34473, 17.34468, 
    17.3447, 17.34464, 17.34466, 17.34477, 17.34476, 17.34474, 17.34475, 
    17.34473, 17.34472, 17.34472, 17.34471, 17.34471, 17.34471, 17.34471, 
    17.34471, 17.34473, 17.34472, 17.34475, 17.34474, 17.34474, 17.34475, 
    17.34474, 17.34472, 17.34472, 17.34472, 17.34471, 17.34473, 17.34468, 
    17.34471, 17.34476, 17.34475, 17.34475, 17.34475, 17.34472, 17.34473, 
    17.34471, 17.34471, 17.3447, 17.34471, 17.34471, 17.34472, 17.34472, 
    17.34473, 17.34474, 17.34475, 17.34475, 17.34474, 17.34472, 17.34471, 
    17.34471, 17.3447, 17.34473, 17.34472, 17.34472, 17.34471, 17.34474, 
    17.34472, 17.34474, 17.34474, 17.34473, 17.34472, 17.34472, 17.34471, 
    17.34471, 17.34472, 17.34472, 17.34473, 17.34473, 17.34474, 17.34475, 
    17.34474, 17.34474, 17.34472, 17.34471, 17.3447, 17.3447, 17.34468, 
    17.34469, 17.34468, 17.34469, 17.34466, 17.34472, 17.34469, 17.34473, 
    17.34473, 17.34472, 17.3447, 17.34471, 17.3447, 17.34472, 17.34474, 
    17.34474, 17.34475, 17.34474, 17.34474, 17.34474, 17.34474, 17.34472, 
    17.34473, 17.34471, 17.3447, 17.34468, 17.34466, 17.34465, 17.34464, 
    17.34464, 17.34464 ;

 SOILC_HR =
  6.215665e-08, 6.243071e-08, 6.237744e-08, 6.25985e-08, 6.247588e-08, 
    6.262062e-08, 6.221222e-08, 6.244159e-08, 6.229516e-08, 6.218133e-08, 
    6.302749e-08, 6.260836e-08, 6.346296e-08, 6.319562e-08, 6.386725e-08, 
    6.342135e-08, 6.395716e-08, 6.38544e-08, 6.416374e-08, 6.407512e-08, 
    6.447078e-08, 6.420464e-08, 6.467591e-08, 6.440724e-08, 6.444926e-08, 
    6.419586e-08, 6.269272e-08, 6.29753e-08, 6.267597e-08, 6.271627e-08, 
    6.269819e-08, 6.247841e-08, 6.236764e-08, 6.213571e-08, 6.217782e-08, 
    6.234817e-08, 6.273439e-08, 6.260329e-08, 6.293373e-08, 6.292627e-08, 
    6.329415e-08, 6.312828e-08, 6.374665e-08, 6.357089e-08, 6.407881e-08, 
    6.395107e-08, 6.407281e-08, 6.40359e-08, 6.407329e-08, 6.388595e-08, 
    6.396621e-08, 6.380137e-08, 6.315934e-08, 6.334801e-08, 6.27853e-08, 
    6.244696e-08, 6.222228e-08, 6.206283e-08, 6.208537e-08, 6.212834e-08, 
    6.234917e-08, 6.255681e-08, 6.271505e-08, 6.28209e-08, 6.29252e-08, 
    6.324087e-08, 6.3408e-08, 6.378219e-08, 6.371467e-08, 6.382906e-08, 
    6.393837e-08, 6.412186e-08, 6.409167e-08, 6.41725e-08, 6.382605e-08, 
    6.40563e-08, 6.36762e-08, 6.378016e-08, 6.29535e-08, 6.263866e-08, 
    6.25048e-08, 6.238768e-08, 6.21027e-08, 6.22995e-08, 6.222191e-08, 
    6.24065e-08, 6.252378e-08, 6.246577e-08, 6.282379e-08, 6.26846e-08, 
    6.34179e-08, 6.310203e-08, 6.392562e-08, 6.372853e-08, 6.397286e-08, 
    6.384818e-08, 6.40618e-08, 6.386955e-08, 6.42026e-08, 6.427513e-08, 
    6.422556e-08, 6.441596e-08, 6.385889e-08, 6.407281e-08, 6.246415e-08, 
    6.247361e-08, 6.251769e-08, 6.232393e-08, 6.231208e-08, 6.213455e-08, 
    6.229253e-08, 6.23598e-08, 6.253058e-08, 6.263159e-08, 6.272763e-08, 
    6.293877e-08, 6.317458e-08, 6.350436e-08, 6.37413e-08, 6.390013e-08, 
    6.380274e-08, 6.388873e-08, 6.37926e-08, 6.374756e-08, 6.424796e-08, 
    6.396696e-08, 6.438858e-08, 6.436525e-08, 6.417443e-08, 6.436788e-08, 
    6.248025e-08, 6.242581e-08, 6.223679e-08, 6.238472e-08, 6.211522e-08, 
    6.226607e-08, 6.23528e-08, 6.26875e-08, 6.276105e-08, 6.282924e-08, 
    6.296392e-08, 6.313677e-08, 6.343999e-08, 6.370384e-08, 6.394473e-08, 
    6.392708e-08, 6.393329e-08, 6.398709e-08, 6.385381e-08, 6.400898e-08, 
    6.403502e-08, 6.396693e-08, 6.436213e-08, 6.424923e-08, 6.436476e-08, 
    6.429125e-08, 6.244351e-08, 6.253511e-08, 6.248561e-08, 6.257869e-08, 
    6.251312e-08, 6.28047e-08, 6.289213e-08, 6.330126e-08, 6.313336e-08, 
    6.340058e-08, 6.316051e-08, 6.320305e-08, 6.340928e-08, 6.317349e-08, 
    6.368928e-08, 6.333956e-08, 6.398919e-08, 6.363992e-08, 6.401108e-08, 
    6.394369e-08, 6.405527e-08, 6.41552e-08, 6.428095e-08, 6.451294e-08, 
    6.445922e-08, 6.465324e-08, 6.267168e-08, 6.279049e-08, 6.278004e-08, 
    6.290439e-08, 6.299635e-08, 6.319569e-08, 6.351541e-08, 6.339518e-08, 
    6.361591e-08, 6.366022e-08, 6.332489e-08, 6.353077e-08, 6.287001e-08, 
    6.297676e-08, 6.291321e-08, 6.268105e-08, 6.342287e-08, 6.304215e-08, 
    6.374522e-08, 6.353896e-08, 6.414095e-08, 6.384155e-08, 6.442965e-08, 
    6.468104e-08, 6.491769e-08, 6.519421e-08, 6.285535e-08, 6.277462e-08, 
    6.291918e-08, 6.311918e-08, 6.330479e-08, 6.355153e-08, 6.357678e-08, 
    6.362301e-08, 6.374275e-08, 6.384343e-08, 6.363761e-08, 6.386867e-08, 
    6.300149e-08, 6.345593e-08, 6.274409e-08, 6.295841e-08, 6.31074e-08, 
    6.304205e-08, 6.338144e-08, 6.346144e-08, 6.37865e-08, 6.361847e-08, 
    6.461898e-08, 6.41763e-08, 6.540478e-08, 6.506145e-08, 6.27464e-08, 
    6.285507e-08, 6.323329e-08, 6.305333e-08, 6.356801e-08, 6.36947e-08, 
    6.37977e-08, 6.392935e-08, 6.394357e-08, 6.402158e-08, 6.389375e-08, 
    6.401653e-08, 6.355206e-08, 6.375961e-08, 6.319006e-08, 6.332868e-08, 
    6.326491e-08, 6.319497e-08, 6.341085e-08, 6.364085e-08, 6.364578e-08, 
    6.371953e-08, 6.392733e-08, 6.35701e-08, 6.467609e-08, 6.399301e-08, 
    6.297358e-08, 6.318288e-08, 6.321279e-08, 6.313171e-08, 6.368199e-08, 
    6.34826e-08, 6.401968e-08, 6.387452e-08, 6.411236e-08, 6.399417e-08, 
    6.397678e-08, 6.3825e-08, 6.373049e-08, 6.349174e-08, 6.329749e-08, 
    6.314347e-08, 6.317929e-08, 6.334847e-08, 6.365492e-08, 6.394485e-08, 
    6.388134e-08, 6.409429e-08, 6.353069e-08, 6.3767e-08, 6.367566e-08, 
    6.391384e-08, 6.339199e-08, 6.383632e-08, 6.327841e-08, 6.332733e-08, 
    6.347864e-08, 6.378302e-08, 6.385039e-08, 6.392229e-08, 6.387792e-08, 
    6.366271e-08, 6.362745e-08, 6.347497e-08, 6.343286e-08, 6.331668e-08, 
    6.322048e-08, 6.330837e-08, 6.340066e-08, 6.36628e-08, 6.389904e-08, 
    6.415662e-08, 6.421966e-08, 6.452062e-08, 6.427562e-08, 6.46799e-08, 
    6.433616e-08, 6.493121e-08, 6.38621e-08, 6.432608e-08, 6.348553e-08, 
    6.357608e-08, 6.373985e-08, 6.411551e-08, 6.391272e-08, 6.414989e-08, 
    6.362608e-08, 6.335431e-08, 6.328401e-08, 6.315283e-08, 6.328701e-08, 
    6.32761e-08, 6.340449e-08, 6.336324e-08, 6.367151e-08, 6.350592e-08, 
    6.397634e-08, 6.414802e-08, 6.46329e-08, 6.493014e-08, 6.523275e-08, 
    6.536635e-08, 6.540701e-08, 6.542402e-08 ;

 SOILC_LOSS =
  6.215665e-08, 6.243071e-08, 6.237744e-08, 6.25985e-08, 6.247588e-08, 
    6.262062e-08, 6.221222e-08, 6.244159e-08, 6.229516e-08, 6.218133e-08, 
    6.302749e-08, 6.260836e-08, 6.346296e-08, 6.319562e-08, 6.386725e-08, 
    6.342135e-08, 6.395716e-08, 6.38544e-08, 6.416374e-08, 6.407512e-08, 
    6.447078e-08, 6.420464e-08, 6.467591e-08, 6.440724e-08, 6.444926e-08, 
    6.419586e-08, 6.269272e-08, 6.29753e-08, 6.267597e-08, 6.271627e-08, 
    6.269819e-08, 6.247841e-08, 6.236764e-08, 6.213571e-08, 6.217782e-08, 
    6.234817e-08, 6.273439e-08, 6.260329e-08, 6.293373e-08, 6.292627e-08, 
    6.329415e-08, 6.312828e-08, 6.374665e-08, 6.357089e-08, 6.407881e-08, 
    6.395107e-08, 6.407281e-08, 6.40359e-08, 6.407329e-08, 6.388595e-08, 
    6.396621e-08, 6.380137e-08, 6.315934e-08, 6.334801e-08, 6.27853e-08, 
    6.244696e-08, 6.222228e-08, 6.206283e-08, 6.208537e-08, 6.212834e-08, 
    6.234917e-08, 6.255681e-08, 6.271505e-08, 6.28209e-08, 6.29252e-08, 
    6.324087e-08, 6.3408e-08, 6.378219e-08, 6.371467e-08, 6.382906e-08, 
    6.393837e-08, 6.412186e-08, 6.409167e-08, 6.41725e-08, 6.382605e-08, 
    6.40563e-08, 6.36762e-08, 6.378016e-08, 6.29535e-08, 6.263866e-08, 
    6.25048e-08, 6.238768e-08, 6.21027e-08, 6.22995e-08, 6.222191e-08, 
    6.24065e-08, 6.252378e-08, 6.246577e-08, 6.282379e-08, 6.26846e-08, 
    6.34179e-08, 6.310203e-08, 6.392562e-08, 6.372853e-08, 6.397286e-08, 
    6.384818e-08, 6.40618e-08, 6.386955e-08, 6.42026e-08, 6.427513e-08, 
    6.422556e-08, 6.441596e-08, 6.385889e-08, 6.407281e-08, 6.246415e-08, 
    6.247361e-08, 6.251769e-08, 6.232393e-08, 6.231208e-08, 6.213455e-08, 
    6.229253e-08, 6.23598e-08, 6.253058e-08, 6.263159e-08, 6.272763e-08, 
    6.293877e-08, 6.317458e-08, 6.350436e-08, 6.37413e-08, 6.390013e-08, 
    6.380274e-08, 6.388873e-08, 6.37926e-08, 6.374756e-08, 6.424796e-08, 
    6.396696e-08, 6.438858e-08, 6.436525e-08, 6.417443e-08, 6.436788e-08, 
    6.248025e-08, 6.242581e-08, 6.223679e-08, 6.238472e-08, 6.211522e-08, 
    6.226607e-08, 6.23528e-08, 6.26875e-08, 6.276105e-08, 6.282924e-08, 
    6.296392e-08, 6.313677e-08, 6.343999e-08, 6.370384e-08, 6.394473e-08, 
    6.392708e-08, 6.393329e-08, 6.398709e-08, 6.385381e-08, 6.400898e-08, 
    6.403502e-08, 6.396693e-08, 6.436213e-08, 6.424923e-08, 6.436476e-08, 
    6.429125e-08, 6.244351e-08, 6.253511e-08, 6.248561e-08, 6.257869e-08, 
    6.251312e-08, 6.28047e-08, 6.289213e-08, 6.330126e-08, 6.313336e-08, 
    6.340058e-08, 6.316051e-08, 6.320305e-08, 6.340928e-08, 6.317349e-08, 
    6.368928e-08, 6.333956e-08, 6.398919e-08, 6.363992e-08, 6.401108e-08, 
    6.394369e-08, 6.405527e-08, 6.41552e-08, 6.428095e-08, 6.451294e-08, 
    6.445922e-08, 6.465324e-08, 6.267168e-08, 6.279049e-08, 6.278004e-08, 
    6.290439e-08, 6.299635e-08, 6.319569e-08, 6.351541e-08, 6.339518e-08, 
    6.361591e-08, 6.366022e-08, 6.332489e-08, 6.353077e-08, 6.287001e-08, 
    6.297676e-08, 6.291321e-08, 6.268105e-08, 6.342287e-08, 6.304215e-08, 
    6.374522e-08, 6.353896e-08, 6.414095e-08, 6.384155e-08, 6.442965e-08, 
    6.468104e-08, 6.491769e-08, 6.519421e-08, 6.285535e-08, 6.277462e-08, 
    6.291918e-08, 6.311918e-08, 6.330479e-08, 6.355153e-08, 6.357678e-08, 
    6.362301e-08, 6.374275e-08, 6.384343e-08, 6.363761e-08, 6.386867e-08, 
    6.300149e-08, 6.345593e-08, 6.274409e-08, 6.295841e-08, 6.31074e-08, 
    6.304205e-08, 6.338144e-08, 6.346144e-08, 6.37865e-08, 6.361847e-08, 
    6.461898e-08, 6.41763e-08, 6.540478e-08, 6.506145e-08, 6.27464e-08, 
    6.285507e-08, 6.323329e-08, 6.305333e-08, 6.356801e-08, 6.36947e-08, 
    6.37977e-08, 6.392935e-08, 6.394357e-08, 6.402158e-08, 6.389375e-08, 
    6.401653e-08, 6.355206e-08, 6.375961e-08, 6.319006e-08, 6.332868e-08, 
    6.326491e-08, 6.319497e-08, 6.341085e-08, 6.364085e-08, 6.364578e-08, 
    6.371953e-08, 6.392733e-08, 6.35701e-08, 6.467609e-08, 6.399301e-08, 
    6.297358e-08, 6.318288e-08, 6.321279e-08, 6.313171e-08, 6.368199e-08, 
    6.34826e-08, 6.401968e-08, 6.387452e-08, 6.411236e-08, 6.399417e-08, 
    6.397678e-08, 6.3825e-08, 6.373049e-08, 6.349174e-08, 6.329749e-08, 
    6.314347e-08, 6.317929e-08, 6.334847e-08, 6.365492e-08, 6.394485e-08, 
    6.388134e-08, 6.409429e-08, 6.353069e-08, 6.3767e-08, 6.367566e-08, 
    6.391384e-08, 6.339199e-08, 6.383632e-08, 6.327841e-08, 6.332733e-08, 
    6.347864e-08, 6.378302e-08, 6.385039e-08, 6.392229e-08, 6.387792e-08, 
    6.366271e-08, 6.362745e-08, 6.347497e-08, 6.343286e-08, 6.331668e-08, 
    6.322048e-08, 6.330837e-08, 6.340066e-08, 6.36628e-08, 6.389904e-08, 
    6.415662e-08, 6.421966e-08, 6.452062e-08, 6.427562e-08, 6.46799e-08, 
    6.433616e-08, 6.493121e-08, 6.38621e-08, 6.432608e-08, 6.348553e-08, 
    6.357608e-08, 6.373985e-08, 6.411551e-08, 6.391272e-08, 6.414989e-08, 
    6.362608e-08, 6.335431e-08, 6.328401e-08, 6.315283e-08, 6.328701e-08, 
    6.32761e-08, 6.340449e-08, 6.336324e-08, 6.367151e-08, 6.350592e-08, 
    6.397634e-08, 6.414802e-08, 6.46329e-08, 6.493014e-08, 6.523275e-08, 
    6.536635e-08, 6.540701e-08, 6.542402e-08 ;

 SOILICE =
  95.04456, 95.48095, 95.396, 95.74871, 95.55294, 95.78405, 95.13291, 
    95.49832, 95.26494, 95.08376, 96.43555, 95.76446, 97.13544, 96.70526, 
    97.78803, 97.06846, 97.9335, 97.76717, 98.26815, 98.12447, 98.84444, 
    98.3345, 99.17878, 98.7409, 98.80936, 98.32026, 95.89923, 96.35187, 
    95.87247, 95.93692, 95.90798, 95.557, 95.38046, 95.01122, 95.07818, 
    95.34939, 95.9659, 95.75632, 96.28497, 96.27301, 96.86364, 96.59707, 
    97.59303, 97.30932, 98.13046, 97.92358, 98.12074, 98.06093, 98.12153, 
    97.81821, 97.9481, 97.68143, 96.64697, 96.95032, 96.04733, 95.50695, 
    95.14893, 94.89542, 94.93123, 94.99954, 95.35098, 95.68208, 95.9349, 
    96.10426, 96.27129, 96.77813, 97.04691, 97.65048, 97.54134, 97.72624, 
    97.903, 98.20026, 98.15129, 98.2824, 97.72132, 98.09402, 97.47922, 
    97.64716, 96.31693, 95.81282, 95.59921, 95.41233, 94.95878, 95.27187, 
    95.14837, 95.44229, 95.62936, 95.5368, 96.10889, 95.88623, 97.06286, 
    96.55497, 97.88238, 97.56374, 97.95883, 97.7571, 98.10293, 97.79165, 
    98.33121, 98.52591, 98.36848, 98.75506, 97.77441, 98.12077, 95.53422, 
    95.54932, 95.61963, 95.31078, 95.2919, 95.00939, 95.26073, 95.3679, 
    95.64021, 95.80154, 95.95504, 96.29308, 96.67149, 97.20211, 97.58437, 
    97.84113, 97.68362, 97.82267, 97.66725, 97.59445, 98.48169, 97.94932, 
    98.71049, 98.67251, 98.28553, 98.67679, 95.55991, 95.47308, 95.17203, 
    95.40757, 94.97866, 95.21862, 95.35678, 95.89092, 96.00848, 96.11763, 
    96.33337, 96.6107, 97.09839, 97.5239, 97.91328, 97.88472, 97.89478, 
    97.9819, 97.7662, 98.01733, 98.05954, 97.94924, 98.66743, 98.48371, 
    98.67171, 98.55209, 95.50129, 95.64745, 95.56846, 95.71704, 95.61237, 
    96.07842, 96.21843, 96.87514, 96.60525, 97.03495, 96.64883, 96.71719, 
    97.04907, 96.66965, 97.50045, 96.93681, 97.98528, 97.42082, 98.02073, 
    97.9116, 98.0923, 98.25433, 98.53535, 98.91306, 98.82553, 99.14176, 
    95.86558, 96.05565, 96.03886, 96.23797, 96.38539, 96.70535, 97.21989, 
    97.02619, 97.38193, 97.45345, 96.91305, 97.24467, 96.18295, 96.35404, 
    96.25212, 95.88058, 97.07085, 96.45891, 97.59071, 97.25783, 98.23122, 
    97.74645, 98.77737, 99.18722, 99.57362, 100.0264, 96.15943, 96.03018, 
    96.26166, 96.58253, 96.88074, 97.27811, 97.31881, 97.39339, 97.58669, 
    97.74942, 97.41702, 97.79023, 96.39382, 97.12407, 95.98138, 96.32465, 
    96.56359, 96.45869, 97.00406, 97.13288, 97.65744, 97.38604, 99.08601, 
    98.28863, 100.3719, 99.80894, 95.98505, 96.15897, 96.76581, 96.47678, 
    97.30466, 97.50911, 97.67548, 97.88844, 97.91142, 98.03775, 97.8308, 
    98.02956, 97.27896, 97.61396, 96.69628, 96.91918, 96.81659, 96.70416, 
    97.05141, 97.42226, 97.43012, 97.54923, 97.88544, 97.30802, 99.17932, 
    97.99172, 96.34884, 96.68485, 96.73283, 96.60256, 97.4886, 97.167, 
    98.03467, 97.7997, 98.18484, 97.99335, 97.9652, 97.7196, 97.56691, 
    97.18175, 96.86902, 96.62144, 96.67897, 96.95105, 97.44495, 97.91354, 
    97.81078, 98.15554, 97.24449, 97.62592, 97.47841, 97.86331, 97.02106, 
    97.73819, 96.83829, 96.91698, 97.16062, 97.65187, 97.76066, 97.87701, 
    97.8052, 97.4575, 97.40057, 97.15469, 97.08689, 96.89983, 96.74517, 
    96.88649, 97.03505, 97.45762, 97.83941, 98.25665, 98.35889, 98.9257, 
    98.52679, 99.18554, 98.62547, 99.59597, 97.77975, 98.60892, 97.1717, 
    97.31767, 97.58209, 98.19006, 97.8615, 98.24579, 97.39835, 96.96047, 
    96.84731, 96.6365, 96.85213, 96.83457, 97.04117, 96.97475, 97.47166, 
    97.20455, 97.96451, 98.24274, 99.10861, 99.59409, 100.0895, 100.3087, 
    100.3755, 100.4034,
  94.71748, 95.18745, 95.09595, 95.47588, 95.26497, 95.51395, 94.8126, 
    95.20617, 94.95478, 94.75967, 96.21598, 95.49284, 96.95303, 96.50356, 
    97.63499, 96.88307, 97.78702, 97.61314, 98.13679, 97.98659, 98.66016, 
    98.20615, 99.00941, 98.55196, 98.62347, 98.19128, 95.63801, 96.12579, 
    95.60918, 95.67862, 95.64744, 95.26936, 95.07925, 94.68155, 94.75365, 
    95.04575, 95.70986, 95.48404, 96.05359, 96.0407, 96.66901, 96.38992, 
    97.43114, 97.13464, 97.99285, 97.7766, 97.9827, 97.92017, 97.98352, 
    97.66647, 97.80224, 97.52351, 96.44267, 96.75958, 95.79758, 95.21551, 
    94.82986, 94.55685, 94.59541, 94.66898, 95.04746, 95.40408, 95.67642, 
    95.85888, 96.03885, 96.57977, 96.86053, 97.49121, 97.37711, 97.57037, 
    97.7551, 98.06584, 98.01463, 98.15171, 97.56521, 97.95479, 97.31218, 
    97.48769, 96.08815, 95.54491, 95.31487, 95.11354, 94.62508, 94.96226, 
    94.82925, 95.14578, 95.3473, 95.24758, 95.86387, 95.624, 96.87719, 
    96.34457, 97.73354, 97.40051, 97.81345, 97.60258, 97.9641, 97.6387, 
    98.20273, 98.3275, 98.24171, 98.56671, 97.6207, 97.98274, 95.2448, 
    95.26107, 95.3368, 95.00418, 94.98383, 94.67959, 94.95025, 95.06567, 
    95.35896, 95.53276, 95.69813, 96.06234, 96.46832, 97.02266, 97.42209, 
    97.69041, 97.5258, 97.67113, 97.50869, 97.4326, 98.28137, 97.80353, 
    98.52016, 98.4805, 98.15498, 98.48497, 95.27248, 95.17894, 94.85472, 
    95.10839, 94.64648, 94.90491, 95.05373, 95.62908, 95.7557, 95.8733, 
    96.10575, 96.40462, 96.91428, 97.3589, 97.76583, 97.73598, 97.74649, 
    97.83757, 97.61211, 97.8746, 97.91874, 97.80343, 98.47519, 98.28344, 
    98.47966, 98.35477, 95.20933, 95.36678, 95.28168, 95.44175, 95.32899, 
    95.83109, 95.98195, 96.68108, 96.39874, 96.84801, 96.4446, 96.51603, 
    96.86283, 96.46635, 97.33443, 96.74551, 97.84111, 97.25126, 97.87815, 
    97.76408, 97.95296, 98.12236, 98.33731, 98.73177, 98.64033, 98.9707, 
    95.60175, 95.80653, 95.78843, 96.00296, 96.16182, 96.50363, 97.04122, 
    96.83882, 97.21052, 97.28526, 96.72061, 97.06712, 95.94369, 96.12807, 
    96.01822, 95.61793, 96.88554, 96.24107, 97.42871, 97.08085, 98.09821, 
    97.59151, 98.59003, 99.01829, 99.42205, 99.89554, 95.91834, 95.77908, 
    96.02847, 96.37429, 96.68688, 97.10206, 97.14456, 97.2225, 97.4245, 
    97.59457, 97.24722, 97.63721, 96.17099, 96.94112, 95.72651, 96.09641, 
    96.35386, 96.24081, 96.81569, 96.95029, 97.49847, 97.21481, 98.91254, 
    98.15826, 100.2567, 99.6681, 95.73046, 95.91783, 96.56683, 96.26029, 
    97.12978, 97.34344, 97.51728, 97.7399, 97.7639, 97.89596, 97.67962, 
    97.88737, 97.10294, 97.453, 96.49416, 96.72704, 96.61983, 96.50239, 
    96.86517, 97.25271, 97.26089, 97.38538, 97.73693, 97.13329, 99.01015, 
    97.84798, 96.12241, 96.48229, 96.53236, 96.39583, 97.32201, 96.98595, 
    97.89272, 97.64712, 98.04971, 97.84953, 97.82011, 97.56341, 97.40383, 
    97.00137, 96.67464, 96.41598, 96.47607, 96.76034, 97.27641, 97.76612, 
    97.65874, 98.01907, 97.06691, 97.46553, 97.31138, 97.71362, 96.83347, 
    97.58299, 96.64251, 96.72472, 96.97929, 97.49268, 97.60632, 97.72795, 
    97.65286, 97.28952, 97.23002, 96.97307, 96.90225, 96.7068, 96.54523, 
    96.69288, 96.84811, 97.28963, 97.68864, 98.12479, 98.23166, 98.74508, 
    98.3285, 99.01666, 98.43165, 99.44556, 97.62637, 98.41425, 96.99084, 
    97.14337, 97.41975, 98.05522, 97.71172, 98.11346, 97.22768, 96.77021, 
    96.65192, 96.43172, 96.65697, 96.63863, 96.85446, 96.78506, 97.30431, 
    97.02517, 97.8194, 98.11026, 98.93609, 99.4435, 99.96143, 100.1907, 
    100.2605, 100.2897,
  128.8469, 129.5346, 129.4007, 129.9567, 129.648, 130.0124, 128.9861, 
    129.562, 129.1941, 128.9087, 131.0403, 129.9816, 132.1454, 131.466, 
    133.1768, 132.0396, 133.4069, 133.1438, 133.9362, 133.7089, 134.7264, 
    134.0412, 135.2553, 134.5626, 134.6708, 134.0187, 130.194, 130.9083, 
    130.1518, 130.2535, 130.2079, 129.6544, 129.3762, 128.7944, 128.8999, 
    129.3272, 130.2992, 129.9687, 130.8026, 130.7837, 131.716, 131.2952, 
    132.8685, 132.4201, 133.7184, 133.3911, 133.703, 133.6084, 133.7043, 
    133.2245, 133.4299, 133.0082, 131.3739, 131.853, 130.4277, 129.5756, 
    129.0114, 128.612, 128.6684, 128.776, 129.3297, 129.8516, 130.2503, 
    130.5174, 130.781, 131.5811, 132.0056, 132.9594, 132.7868, 133.0791, 
    133.3586, 133.8288, 133.7514, 133.9588, 133.0713, 133.6608, 132.6886, 
    132.9541, 130.8531, 130.0578, 129.7211, 129.4264, 128.7118, 129.2051, 
    129.0105, 129.4736, 129.7685, 129.6226, 130.5247, 130.1736, 132.0307, 
    131.2287, 133.326, 132.8222, 133.4469, 133.1279, 133.6749, 133.1825, 
    134.036, 134.2228, 134.095, 134.5849, 133.1553, 133.7031, 129.6185, 
    129.6423, 129.7532, 129.2664, 129.2366, 128.7915, 129.1875, 129.3564, 
    129.7856, 130.04, 130.2821, 130.8154, 131.4127, 132.2507, 132.8548, 
    133.2607, 133.0117, 133.2316, 132.9858, 132.8707, 134.1529, 133.4319, 
    134.5144, 134.4544, 133.9638, 134.4612, 129.659, 129.5221, 129.0477, 
    129.4189, 128.7431, 129.1212, 129.3389, 130.181, 130.3664, 130.5385, 
    130.8789, 131.3167, 132.0869, 132.7592, 133.3749, 133.3297, 133.3456, 
    133.4834, 133.1423, 133.5394, 133.6062, 133.4317, 134.4464, 134.1561, 
    134.4531, 134.2641, 129.5666, 129.797, 129.6725, 129.9068, 129.7417, 
    130.4767, 130.6976, 131.7343, 131.3081, 131.9866, 131.3769, 131.4848, 
    132.009, 131.4097, 132.7222, 131.8316, 133.4888, 132.5964, 133.5448, 
    133.3722, 133.658, 133.9144, 134.2376, 134.8348, 134.6964, 135.1967, 
    130.141, 130.4408, 130.4143, 130.7284, 130.961, 131.4661, 132.2788, 
    131.9728, 132.5348, 132.6479, 131.7941, 132.3179, 130.6416, 130.9116, 
    130.7507, 130.1647, 132.0434, 131.0771, 132.8648, 132.3387, 133.8778, 
    133.1111, 134.6202, 135.2687, 135.8805, 136.5981, 130.6045, 130.4006, 
    130.7658, 131.2722, 131.7431, 132.3708, 132.4351, 132.5529, 132.8585, 
    133.1157, 132.5903, 133.1803, 130.9745, 132.1274, 130.3236, 130.8652, 
    131.2423, 131.0767, 131.9378, 132.1413, 132.9703, 132.5413, 135.1086, 
    133.9687, 137.1457, 136.2533, 130.3294, 130.6038, 131.5616, 131.1053, 
    132.4127, 132.7358, 132.9988, 133.3356, 133.3719, 133.5717, 133.2444, 
    133.5588, 132.3721, 132.9016, 131.4518, 131.8038, 131.6417, 131.4642, 
    132.0126, 132.5986, 132.611, 132.7993, 133.331, 132.418, 135.2564, 
    133.4991, 130.9033, 131.4338, 131.5095, 131.3038, 132.7034, 132.1952, 
    133.5668, 133.1952, 133.8044, 133.5015, 133.457, 133.0686, 132.8272, 
    132.2185, 131.7245, 131.3336, 131.4244, 131.8541, 132.6345, 133.3753, 
    133.2128, 133.7581, 132.3176, 132.9205, 132.6873, 133.2958, 131.9647, 
    133.0981, 131.676, 131.8003, 132.1852, 132.9616, 133.1335, 133.3175, 
    133.2039, 132.6543, 132.5643, 132.1758, 132.0687, 131.7732, 131.529, 
    131.7521, 131.9868, 132.6544, 133.258, 133.9181, 134.0798, 134.8549, 
    134.2242, 135.2662, 134.3803, 135.916, 133.1638, 134.354, 132.2026, 
    132.4333, 132.8512, 133.8127, 133.293, 133.9009, 132.5608, 131.869, 
    131.6902, 131.3574, 131.6978, 131.6701, 131.9964, 131.8915, 132.6767, 
    132.2545, 133.4559, 133.8961, 135.1443, 135.9129, 136.698, 137.0455, 
    137.1514, 137.1957,
  193.9548, 195.0306, 194.8211, 195.6913, 195.2081, 195.7785, 194.1725, 
    195.0734, 194.4979, 194.0514, 197.3885, 195.7302, 199.1213, 198.0557, 
    200.7402, 198.9553, 201.1015, 200.6883, 201.9332, 201.576, 203.1748, 
    202.0982, 204.0069, 202.9172, 203.0874, 202.0628, 196.0629, 197.1815, 
    195.9968, 196.156, 196.0845, 195.2182, 194.7828, 193.8727, 194.0377, 
    194.7061, 196.2276, 195.71, 197.016, 196.9865, 198.4479, 197.788, 
    200.256, 199.5522, 201.5909, 201.0768, 201.5667, 201.418, 201.5687, 
    200.8151, 201.1377, 200.4754, 197.9115, 198.6625, 196.4287, 195.0948, 
    194.212, 193.5875, 193.6757, 193.8439, 194.7101, 195.5268, 196.151, 
    196.5694, 196.9822, 198.2362, 198.9019, 200.3987, 200.1278, 200.5867, 
    201.0257, 201.7644, 201.6427, 201.9687, 200.5745, 201.5003, 199.9736, 
    200.3904, 197.0951, 195.8495, 195.3224, 194.8613, 193.7435, 194.515, 
    194.2106, 194.9352, 195.3967, 195.1683, 196.5808, 196.0308, 198.9414, 
    197.6838, 200.9744, 200.1833, 201.1644, 200.6633, 201.5224, 200.7491, 
    202.09, 202.3829, 202.1828, 202.9524, 200.7063, 201.5668, 195.162, 
    195.1992, 195.3727, 194.611, 194.5644, 193.8682, 194.4875, 194.7518, 
    195.4235, 195.8217, 196.2007, 197.0361, 197.9722, 199.2865, 200.2346, 
    200.872, 200.4809, 200.8261, 200.4403, 200.2596, 202.2732, 201.1407, 
    202.8415, 202.7471, 201.9764, 202.7578, 195.2254, 195.0111, 194.2689, 
    194.8496, 193.7925, 194.3838, 194.7244, 196.0424, 196.3327, 196.6024, 
    197.1357, 197.8217, 199.0294, 200.0845, 201.0512, 200.9802, 201.0052, 
    201.2217, 200.6859, 201.3097, 201.4146, 201.1405, 202.7345, 202.2781, 
    202.7451, 202.4479, 195.0807, 195.4413, 195.2464, 195.6131, 195.3548, 
    196.5056, 196.8516, 198.4764, 197.8082, 198.8722, 197.916, 198.0853, 
    198.9072, 197.9676, 200.0264, 198.6291, 201.2301, 199.8288, 201.3181, 
    201.047, 201.496, 201.8988, 202.4063, 203.3454, 203.1276, 203.9147, 
    195.9798, 196.4493, 196.4078, 196.8998, 197.2643, 198.0559, 199.3305, 
    198.8505, 199.7323, 199.9097, 198.5702, 199.392, 196.7639, 197.1868, 
    196.9348, 196.0169, 198.9612, 197.4462, 200.2503, 199.4246, 201.8414, 
    200.6369, 203.0078, 204.028, 204.991, 206.1212, 196.7057, 196.3864, 
    196.9584, 197.752, 198.4902, 199.4749, 199.5758, 199.7607, 200.2403, 
    200.6442, 199.8194, 200.7456, 197.2852, 199.093, 196.2658, 197.1142, 
    197.7051, 197.4456, 198.7956, 199.1149, 200.4159, 199.7425, 203.776, 
    201.9842, 206.9845, 205.5781, 196.2749, 196.7046, 198.2056, 197.4904, 
    199.5407, 200.0478, 200.4607, 200.9895, 201.0466, 201.3605, 200.8463, 
    201.3401, 199.477, 200.308, 198.0335, 198.5854, 198.3313, 198.053, 
    198.913, 199.8324, 199.8519, 200.1474, 200.9822, 199.549, 204.0084, 
    201.2462, 197.1739, 198.0052, 198.124, 197.8015, 199.9969, 199.1994, 
    201.3528, 200.7691, 201.7261, 201.2501, 201.1802, 200.5702, 200.1912, 
    199.236, 198.4612, 197.8483, 197.9906, 198.6643, 199.8887, 201.0518, 
    200.7966, 201.6532, 199.3915, 200.3377, 199.9717, 200.9271, 198.8378, 
    200.6165, 198.3851, 198.5799, 199.1836, 200.4021, 200.6722, 200.9611, 
    200.7827, 199.9198, 199.7786, 199.1689, 199.0009, 198.5375, 198.1545, 
    198.5044, 198.8725, 199.9201, 200.8677, 201.9046, 202.1589, 203.3769, 
    202.3852, 204.0239, 202.6305, 205.0468, 200.7196, 202.5892, 199.2111, 
    199.573, 200.2289, 201.7391, 200.9226, 201.8776, 199.773, 198.6877, 
    198.4074, 197.8855, 198.4193, 198.3759, 198.8876, 198.723, 199.9549, 
    199.2925, 201.1785, 201.87, 203.8322, 205.0421, 206.2788, 206.8266, 
    206.9935, 207.0634,
  318.312, 320.1113, 319.7607, 321.2175, 320.4086, 321.3636, 318.676, 
    320.183, 319.2202, 318.4735, 324.0625, 321.2826, 326.9049, 325.1748, 
    329.5376, 326.6352, 330.1258, 329.4533, 331.4809, 330.8988, 333.506, 
    331.7499, 334.8651, 333.0857, 333.3635, 331.6922, 321.8401, 323.7153, 
    321.7293, 321.996, 321.8763, 320.4253, 319.6966, 318.1748, 318.4505, 
    319.5684, 322.116, 321.2489, 323.4379, 323.3883, 325.8113, 324.7332, 
    328.7498, 327.6053, 330.9231, 330.0857, 330.8837, 330.6415, 330.8869, 
    329.6595, 330.1849, 329.1068, 324.9405, 326.1598, 322.4531, 320.2187, 
    318.742, 317.6981, 317.8455, 318.1267, 319.575, 320.9421, 321.9877, 
    322.6889, 323.3812, 325.4676, 326.5485, 328.9819, 328.5412, 329.2879, 
    330.0024, 331.2058, 331.0074, 331.5387, 329.268, 330.7755, 328.2905, 
    328.9684, 323.5703, 321.4826, 320.5997, 319.8281, 317.9589, 319.2487, 
    318.7397, 319.9518, 320.7243, 320.3419, 322.7081, 321.7863, 326.6127, 
    324.5583, 329.919, 328.6316, 330.2283, 329.4126, 330.8116, 329.5522, 
    331.7366, 332.2141, 331.8878, 333.1431, 329.4826, 330.8838, 320.3313, 
    320.3936, 320.6841, 319.4092, 319.3313, 318.1673, 319.2028, 319.6448, 
    320.769, 321.4359, 322.071, 323.4715, 325.0392, 327.1734, 328.7149, 
    329.7522, 329.1157, 329.6776, 329.0496, 328.7556, 332.0352, 330.1898, 
    332.9623, 332.8082, 331.5514, 332.8256, 320.4374, 320.0788, 318.8372, 
    319.8085, 318.0407, 319.0292, 319.5989, 321.8057, 322.2922, 322.7443, 
    323.6386, 324.7899, 326.7557, 328.4708, 330.044, 329.9285, 329.9692, 
    330.3216, 329.4494, 330.4651, 330.6359, 330.1895, 332.7876, 332.0433, 
    332.805, 332.3201, 320.1953, 320.799, 320.4727, 321.0866, 320.654, 
    322.5819, 323.162, 325.8575, 324.7672, 326.5003, 324.9482, 325.2227, 
    326.5572, 325.0318, 328.3762, 326.1055, 330.3354, 328.0549, 330.4788, 
    330.0372, 330.7685, 331.4249, 332.2523, 333.7846, 333.4292, 334.7144, 
    321.7008, 322.4875, 322.4181, 323.243, 323.8544, 325.1751, 327.245, 
    326.4651, 327.8981, 328.1866, 326.0099, 327.3448, 323.0149, 323.7243, 
    323.3017, 321.7629, 326.6449, 324.1595, 328.7405, 327.3978, 331.3313, 
    329.3695, 333.2337, 334.8995, 336.474, 338.3241, 322.9175, 322.3821, 
    323.3412, 324.6728, 325.88, 327.4796, 327.6436, 327.9443, 328.7243, 
    329.3815, 328.0396, 329.5465, 323.8893, 326.8591, 322.18, 323.6024, 
    324.5941, 324.1586, 326.376, 326.8946, 329.0099, 327.9147, 334.4877, 
    331.5639, 339.739, 337.4348, 322.1953, 322.9156, 325.4181, 324.2337, 
    327.5866, 328.4111, 329.0828, 329.9436, 330.0365, 330.5477, 329.7105, 
    330.5145, 327.483, 328.8344, 325.1388, 326.0346, 325.6221, 325.1704, 
    326.5666, 328.0607, 328.0925, 328.5731, 329.9314, 327.6001, 334.8674, 
    330.3614, 323.7028, 325.0929, 325.2856, 324.756, 328.3284, 327.032, 
    330.5352, 329.5847, 331.1434, 330.368, 330.2541, 329.2611, 328.6444, 
    327.0913, 325.8329, 324.8345, 325.0692, 326.1628, 328.1523, 330.045, 
    329.6295, 331.0247, 327.3441, 328.8827, 328.2873, 329.8419, 326.4445, 
    329.3362, 325.7094, 326.0258, 327.0063, 328.9874, 329.427, 329.8973, 
    329.607, 328.2029, 327.9733, 326.9824, 326.7094, 325.9568, 325.3351, 
    325.9032, 326.5008, 328.2034, 329.7453, 331.4343, 331.8488, 333.836, 
    332.2178, 334.8927, 332.6177, 336.5652, 329.5041, 332.5505, 327.0509, 
    327.639, 328.7057, 331.1645, 329.8346, 331.3903, 327.9643, 326.2007, 
    325.7456, 324.897, 325.765, 325.6944, 326.5254, 326.2581, 328.26, 
    327.1832, 330.2513, 331.3779, 334.5796, 336.5575, 338.5823, 339.4802, 
    339.7539, 339.8684,
  524.2802, 527.5528, 526.9146, 529.5684, 528.0942, 529.8349, 524.9416, 
    527.6833, 525.931, 524.5736, 534.7657, 529.6872, 540.1031, 536.8177, 
    545.1176, 539.5904, 546.2406, 544.9568, 548.8311, 547.7177, 552.7115, 
    549.3459, 555.3222, 551.9052, 552.4382, 549.2354, 530.7042, 534.1304, 
    530.5021, 530.9888, 530.7702, 528.1247, 526.7978, 524.0309, 524.5319, 
    526.5646, 531.2078, 529.6258, 533.6231, 533.5324, 538.0255, 535.9939, 
    543.6154, 541.4355, 547.7641, 546.1639, 547.6888, 547.2258, 547.6949, 
    545.3505, 546.3534, 544.296, 536.3737, 538.6873, 531.8234, 527.7482, 
    525.0615, 523.1646, 523.4329, 523.9435, 526.5765, 529.0663, 530.9736, 
    532.254, 533.5194, 537.3729, 539.4256, 544.0576, 543.2178, 544.6412, 
    546.0051, 548.3048, 547.9254, 548.9417, 544.6034, 547.4819, 542.7401, 
    544.032, 533.8652, 530.0519, 528.4423, 527.0372, 523.6387, 525.9829, 
    525.0573, 527.2623, 528.6694, 527.9728, 532.2891, 530.606, 539.5476, 
    535.6736, 545.8458, 543.39, 546.4364, 544.8792, 547.5509, 545.1456, 
    549.3204, 550.2349, 549.6097, 552.0154, 545.0127, 547.689, 527.9534, 
    528.0669, 528.5961, 526.2748, 526.1332, 524.0172, 525.8994, 526.7035, 
    528.751, 529.9668, 531.1257, 533.6846, 536.5605, 540.6136, 543.5488, 
    545.5273, 544.313, 545.3849, 544.1868, 543.6263, 549.8921, 546.3629, 
    551.6686, 551.3733, 548.9659, 551.4066, 528.1466, 527.4937, 525.2346, 
    527.0015, 523.7874, 525.5837, 526.6201, 530.6414, 531.5296, 532.3553, 
    533.9902, 536.0977, 539.8195, 543.0836, 546.0845, 545.8639, 545.9415, 
    546.6147, 544.9494, 546.8887, 547.2151, 546.3623, 551.3338, 549.9077, 
    551.367, 550.4379, 527.7057, 528.8055, 528.2109, 529.3298, 528.5413, 
    532.0585, 533.1186, 538.1132, 536.0562, 539.3342, 536.3879, 536.9086, 
    539.442, 536.5466, 542.9032, 538.584, 546.6409, 542.2913, 546.9149, 
    546.0715, 547.4687, 548.7239, 550.308, 553.2464, 552.5641, 555.0326, 
    530.4501, 531.8862, 531.7594, 533.2668, 534.385, 536.8184, 540.7499, 
    539.2672, 541.9928, 542.5421, 538.4026, 540.9398, 532.8499, 534.147, 
    533.3741, 530.5634, 539.6088, 534.9434, 543.5975, 541.0406, 548.5448, 
    544.797, 552.1891, 555.3882, 558.3942, 561.8449, 532.6718, 531.6937, 
    533.4464, 535.8833, 538.156, 541.1962, 541.5084, 542.0807, 543.5667, 
    544.8199, 542.2621, 545.1347, 534.4489, 540.016, 531.3247, 533.924, 
    535.7391, 534.9417, 539.098, 540.0835, 544.1112, 542.0244, 554.5967, 
    548.9899, 564.4904, 560.185, 531.3525, 532.6683, 537.2792, 535.0792, 
    541.3998, 542.9698, 544.2502, 545.8926, 546.0701, 547.0466, 545.4477, 
    546.9832, 541.2028, 543.7764, 536.7494, 538.4495, 537.6664, 536.8093, 
    539.4601, 542.3024, 542.3629, 543.2784, 545.8692, 541.4256, 555.3264, 
    546.6904, 534.1076, 536.6622, 537.0278, 536.0358, 542.8122, 540.3447, 
    547.0227, 545.2077, 548.1854, 546.7032, 546.4856, 544.5902, 543.4144, 
    540.4576, 538.0665, 536.1794, 536.6175, 538.6929, 542.4767, 546.0864, 
    545.2932, 547.9583, 540.9385, 543.8685, 542.7338, 545.6986, 539.228, 
    544.7332, 537.832, 538.4327, 540.2959, 544.0682, 544.9067, 545.8044, 
    545.2501, 542.5731, 542.1359, 540.2504, 539.7314, 538.3018, 537.1219, 
    538.1999, 539.335, 542.5741, 545.514, 548.7419, 549.5353, 553.3449, 
    550.2418, 555.375, 551.0078, 558.564, 545.0538, 550.8792, 540.3807, 
    541.4996, 543.5312, 548.2256, 545.6846, 548.6576, 542.1188, 538.7648, 
    537.9008, 536.294, 537.9376, 537.8036, 539.3818, 538.874, 542.6821, 
    540.6324, 546.4802, 548.634, 554.7734, 558.5497, 562.3273, 564.006, 
    564.5182, 564.7325,
  947.2507, 954.1235, 952.7804, 958.3742, 955.2639, 958.9371, 948.6368, 
    954.3984, 950.7131, 947.8654, 969.252, 958.625, 980.2917, 973.4848, 
    990.7531, 979.2271, 993.1078, 990.4163, 998.5573, 996.2121, 1006.765, 
    999.6431, 1012.319, 1005.055, 1006.185, 999.4099, 960.7752, 967.944, 
    960.3477, 961.3776, 960.915, 955.3281, 952.5348, 946.7285, 947.7778, 
    952.0444, 961.8413, 958.4954, 966.9009, 966.7145, 975.9829, 971.7838, 
    987.6099, 983.0631, 996.3098, 992.947, 996.1514, 995.1776, 996.1641, 
    991.241, 993.3447, 989.033, 972.5678, 977.3539, 963.1456, 954.5349, 
    948.8883, 944.9172, 945.4769, 946.5455, 952.0695, 957.3141, 961.3454, 
    964.0589, 966.6877, 974.6326, 978.8851, 988.5344, 986.7792, 989.7555, 
    992.6136, 997.4482, 996.6493, 998.7903, 989.6763, 995.7162, 985.7823, 
    988.4808, 967.3987, 959.3959, 955.9976, 953.0384, 945.9076, 950.8221, 
    948.8795, 953.512, 956.4765, 955.0082, 964.1333, 960.5676, 979.1383, 
    971.123, 992.2795, 987.139, 993.519, 990.2537, 995.8612, 990.8118, 
    999.5892, 1001.52, 1000.2, 1005.289, 990.5333, 996.1517, 954.9672, 
    955.2064, 956.3219, 951.4355, 951.1379, 946.6998, 950.6468, 952.3365, 
    956.6487, 959.2159, 961.6675, 967.0273, 972.9534, 981.353, 987.4707, 
    991.6118, 989.0685, 991.3132, 988.8046, 987.6328, 1000.796, 993.3645, 
    1004.554, 1003.929, 998.8414, 1003.999, 955.3744, 953.999, 949.2512, 
    952.9633, 946.2187, 949.9839, 952.161, 960.6424, 962.5231, 964.2736, 
    967.6558, 971.9979, 979.7028, 986.499, 992.7803, 992.3174, 992.4803, 
    993.8933, 990.4006, 994.4689, 995.155, 993.3633, 1003.845, 1000.829, 
    1003.915, 1001.949, 954.4456, 956.7637, 955.5099, 957.8702, 956.2065, 
    963.6442, 965.8643, 976.1646, 971.9122, 978.6954, 972.5971, 973.6727, 
    978.9192, 972.9247, 986.1225, 977.1398, 993.9483, 984.8461, 994.524, 
    992.753, 995.6882, 998.3313, 1001.675, 1007.901, 1006.453, 1011.702, 
    960.2377, 963.2789, 963.01, 966.1687, 968.4681, 973.4862, 981.6363, 
    978.5566, 984.2238, 985.3691, 976.7642, 982.0312, 965.3124, 967.9783, 
    966.389, 960.4773, 979.2653, 969.6177, 987.5725, 982.2411, 997.9537, 
    990.0816, 1005.657, 1012.46, 1018.94, 1026.619, 964.9453, 962.8708, 
    966.5376, 971.5555, 976.2532, 982.5649, 983.2147, 984.4072, 987.5081, 
    990.1296, 984.7853, 990.7888, 968.5995, 980.1109, 962.089, 967.5195, 
    971.2582, 969.6144, 978.2056, 980.2512, 988.6464, 984.2896, 1010.773, 
    998.892, 1032.424, 1022.919, 962.1479, 964.9379, 974.4387, 969.8976, 
    982.9887, 986.2617, 988.9371, 992.3777, 992.7501, 994.8007, 991.4447, 
    994.6675, 982.5784, 987.9465, 973.3437, 976.8611, 975.2399, 973.4677, 
    978.9567, 984.8691, 984.9954, 986.9059, 992.3286, 983.0424, 1012.328, 
    994.0522, 967.8973, 973.1636, 973.9192, 971.8702, 985.9327, 980.794, 
    994.7505, 990.9418, 997.1965, 994.0793, 993.6223, 989.6486, 987.1899, 
    981.0286, 976.0679, 972.1667, 973.0712, 977.3655, 985.2327, 992.7842, 
    991.1209, 996.7186, 982.0285, 988.139, 985.7692, 991.9708, 978.4752, 
    989.9479, 975.5825, 976.8263, 980.6924, 988.5566, 990.3112, 992.1926, 
    991.0307, 985.4338, 984.5222, 980.598, 979.52, 976.5552, 974.1135, 
    976.3441, 978.697, 985.4359, 991.5839, 998.3691, 1000.043, 1008.11, 
    1001.535, 1012.431, 1003.155, 1019.317, 990.6193, 1002.883, 980.8688, 
    983.1965, 987.434, 997.2814, 991.9415, 998.1915, 984.4865, 977.5147, 
    975.7249, 972.4033, 975.8011, 975.5239, 978.7942, 977.741, 985.6611, 
    981.392, 993.611, 998.1417, 1011.149, 1019.285, 1027.696, 1031.374, 
    1032.485, 1032.95,
  1829.891, 1849.353, 1845.525, 1861.55, 1852.613, 1863.174, 1833.791, 
    1850.138, 1839.656, 1831.619, 1893.772, 1862.273, 1928.094, 1906.814, 
    1960.69, 1924.74, 1968.121, 1959.631, 1985.506, 1977.992, 2012.212, 
    1989.003, 2030.647, 2006.595, 2010.303, 1988.251, 1868.494, 1889.771, 
    1867.255, 1870.243, 1868.9, 1852.797, 1844.826, 1828.425, 1831.373, 
    1843.432, 1871.59, 1861.899, 1886.589, 1886.021, 1914.579, 1901.555, 
    1950.847, 1936.758, 1978.304, 1967.612, 1977.798, 1974.693, 1977.839, 
    1962.226, 1968.871, 1955.293, 1903.976, 1918.863, 1875.39, 1850.528, 
    1834.5, 1823.354, 1824.918, 1827.912, 1843.504, 1858.496, 1870.149, 
    1878.057, 1885.94, 1910.375, 1923.665, 1953.734, 1948.26, 1957.557, 
    1966.557, 1981.946, 1979.389, 1986.256, 1957.309, 1976.409, 1945.163, 
    1953.566, 1888.106, 1864.5, 1854.715, 1846.259, 1826.124, 1839.965, 
    1834.475, 1847.609, 1856.089, 1851.881, 1878.275, 1867.892, 1924.461, 
    1899.519, 1965.501, 1949.38, 1969.423, 1959.12, 1976.872, 1960.875, 
    1988.829, 1995.073, 1990.8, 2007.361, 1959.999, 1977.799, 1851.764, 
    1852.448, 1855.646, 1841.704, 1840.86, 1828.345, 1839.469, 1844.262, 
    1856.583, 1863.979, 1871.085, 1886.974, 1905.169, 1931.447, 1950.413, 
    1963.394, 1955.404, 1962.453, 1954.578, 1950.919, 1992.728, 1968.934, 
    2004.954, 2002.91, 1986.421, 2003.14, 1852.929, 1848.998, 1835.524, 
    1846.045, 1826.996, 1837.593, 1843.764, 1868.109, 1873.575, 1878.685, 
    1888.891, 1902.216, 1926.238, 1947.389, 1967.084, 1965.621, 1966.136, 
    1970.61, 1959.582, 1972.438, 1974.621, 1968.93, 2002.636, 1992.834, 
    2002.866, 1996.466, 1850.273, 1856.914, 1853.318, 1860.097, 1855.314, 
    1876.845, 1883.436, 1915.146, 1901.952, 1923.069, 1904.067, 1907.396, 
    1923.772, 1905.08, 1946.219, 1918.193, 1970.785, 1942.262, 1972.613, 
    1966.998, 1976.32, 1984.78, 1995.575, 2015.957, 2011.182, 2028.583, 
    1866.936, 1875.779, 1874.994, 1884.361, 1891.372, 1906.818, 1932.344, 
    1922.633, 1940.339, 1943.882, 1917.018, 1933.585, 1881.76, 1889.875, 
    1885.031, 1867.63, 1924.861, 1894.893, 1950.731, 1934.23, 1983.568, 
    1958.58, 2008.569, 2031.119, 2053.034, 2079.239, 1880.652, 1874.588, 
    1885.483, 1900.852, 1915.422, 1935.225, 1937.225, 1940.905, 1950.53, 
    1958.731, 1942.074, 1960.803, 1891.774, 1927.524, 1872.311, 1888.475, 
    1899.935, 1894.883, 1921.531, 1927.966, 1954.084, 1940.542, 2025.485, 
    1986.583, 2099.508, 2066.705, 1872.483, 1880.63, 1909.773, 1895.752, 
    1936.529, 1946.652, 1954.993, 1965.812, 1966.989, 1973.493, 1962.868, 
    1973.07, 1935.267, 1951.897, 1906.377, 1917.321, 1912.264, 1906.761, 
    1923.89, 1942.334, 1942.724, 1948.654, 1965.656, 1936.695, 2030.677, 
    1971.115, 1889.628, 1905.819, 1908.16, 1901.822, 1945.63, 1929.68, 
    1973.333, 1961.284, 1981.14, 1971.2, 1969.75, 1957.222, 1949.539, 
    1930.421, 1914.844, 1902.737, 1905.533, 1918.899, 1943.46, 1967.097, 
    1961.848, 1979.61, 1933.577, 1952.498, 1945.122, 1964.527, 1922.377, 
    1958.161, 1913.331, 1917.212, 1929.359, 1953.803, 1959.301, 1965.227, 
    1961.564, 1944.083, 1941.261, 1929.061, 1925.662, 1916.365, 1908.763, 
    1915.706, 1923.074, 1944.089, 1963.306, 1984.902, 1990.293, 2016.649, 
    1995.121, 2031.024, 2000.386, 2054.32, 1960.269, 1999.5, 1929.916, 
    1937.17, 1950.299, 1981.412, 1964.434, 1984.331, 1941.15, 1919.366, 
    1913.775, 1903.468, 1914.012, 1913.148, 1923.379, 1920.075, 1944.787, 
    1931.57, 1969.715, 1984.171, 2026.74, 2054.212, 2082.899, 2095.76, 
    2099.724, 2101.388,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.536441, 4.554934, 4.551334, 4.56628, 4.557984, 4.567778, 4.540185, 
    4.55567, 4.54578, 4.538103, 4.595385, 4.566948, 4.625044, 4.606815, 
    4.652697, 4.622205, 4.658861, 4.651813, 4.673042, 4.666954, 4.694181, 
    4.675854, 4.708333, 4.689799, 4.692696, 4.67525, 4.572659, 4.591839, 
    4.571525, 4.574256, 4.57303, 4.558156, 4.550675, 4.535029, 4.537866, 
    4.549359, 4.575484, 4.566603, 4.589005, 4.588498, 4.613526, 4.60223, 
    4.644434, 4.632412, 4.667208, 4.658441, 4.666796, 4.664261, 4.666829, 
    4.653975, 4.65948, 4.64818, 4.604345, 4.617199, 4.578935, 4.556035, 
    4.540864, 4.530121, 4.531639, 4.534534, 4.549426, 4.563457, 4.574171, 
    4.581347, 4.588425, 4.609902, 4.621292, 4.646869, 4.642244, 4.650079, 
    4.657569, 4.670166, 4.66809, 4.673646, 4.64987, 4.665663, 4.639612, 
    4.646728, 4.590358, 4.568997, 4.559945, 4.552026, 4.532806, 4.546073, 
    4.540841, 4.553296, 4.561224, 4.557301, 4.581543, 4.572108, 4.621968, 
    4.600446, 4.656695, 4.643193, 4.659935, 4.651386, 4.666041, 4.652851, 
    4.675714, 4.680703, 4.677294, 4.690398, 4.65212, 4.666797, 4.557191, 
    4.557831, 4.560811, 4.547723, 4.546923, 4.534951, 4.545602, 4.550143, 
    4.561683, 4.568519, 4.575024, 4.589348, 4.605384, 4.627869, 4.644067, 
    4.654947, 4.648273, 4.654165, 4.647579, 4.644495, 4.678834, 4.659532, 
    4.688512, 4.686905, 4.673779, 4.687086, 4.55828, 4.5546, 4.541843, 
    4.551825, 4.533649, 4.543818, 4.549672, 4.572307, 4.577289, 4.581914, 
    4.591056, 4.602808, 4.623474, 4.641505, 4.658005, 4.656795, 4.65722, 
    4.660912, 4.651772, 4.662414, 4.664202, 4.659528, 4.686689, 4.678919, 
    4.686871, 4.68181, 4.555796, 4.56199, 4.558642, 4.564939, 4.560503, 
    4.580252, 4.586185, 4.614014, 4.602577, 4.620785, 4.604424, 4.60732, 
    4.621383, 4.605307, 4.640511, 4.616626, 4.661056, 4.637136, 4.662558, 
    4.657933, 4.665591, 4.672456, 4.681102, 4.697085, 4.69338, 4.706766, 
    4.571233, 4.579287, 4.578577, 4.587013, 4.59326, 4.606819, 4.628623, 
    4.620415, 4.635489, 4.638519, 4.61562, 4.629672, 4.584682, 4.591932, 
    4.587613, 4.571869, 4.622307, 4.596375, 4.644336, 4.63023, 4.671477, 
    4.650935, 4.691342, 4.70869, 4.725049, 4.744221, 4.583685, 4.578208, 
    4.588017, 4.601614, 4.614251, 4.63109, 4.632814, 4.635974, 4.644166, 
    4.651061, 4.636975, 4.652791, 4.593616, 4.624562, 4.57614, 4.590686, 
    4.600811, 4.596366, 4.619477, 4.624936, 4.647163, 4.635663, 4.704406, 
    4.673909, 4.758848, 4.735012, 4.576296, 4.583666, 4.609381, 4.597133, 
    4.632215, 4.640878, 4.647928, 4.656952, 4.657926, 4.663279, 4.65451, 
    4.662932, 4.631125, 4.645321, 4.606435, 4.61588, 4.611533, 4.606769, 
    4.621483, 4.637197, 4.637531, 4.642578, 4.656824, 4.632357, 4.708355, 
    4.661327, 4.591712, 4.60595, 4.607984, 4.602463, 4.640009, 4.626381, 
    4.663148, 4.653192, 4.669512, 4.661397, 4.660204, 4.649798, 4.643327, 
    4.627006, 4.613754, 4.603263, 4.605701, 4.61723, 4.638159, 4.658015, 
    4.653661, 4.66827, 4.629665, 4.645828, 4.639577, 4.655887, 4.620197, 
    4.650584, 4.612452, 4.615787, 4.626111, 4.646927, 4.651537, 4.656468, 
    4.653425, 4.638691, 4.636279, 4.625859, 4.622986, 4.61506, 4.608506, 
    4.614495, 4.62079, 4.638696, 4.654874, 4.672554, 4.676887, 4.697619, 
    4.680741, 4.708619, 4.684915, 4.725995, 4.652346, 4.684215, 4.62658, 
    4.632766, 4.64397, 4.669733, 4.65581, 4.672094, 4.636184, 4.61763, 
    4.612834, 4.603901, 4.613039, 4.612295, 4.621049, 4.618235, 4.639291, 
    4.627973, 4.660175, 4.671965, 4.705362, 4.725915, 4.746893, 4.756175, 
    4.759001, 4.760184,
  5.625641, 5.648898, 5.64437, 5.66317, 5.652735, 5.665053, 5.63035, 
    5.649823, 5.637385, 5.627731, 5.699788, 5.664009, 5.737118, 5.714172, 
    5.771936, 5.733544, 5.7797, 5.770824, 5.797562, 5.789893, 5.824194, 
    5.801104, 5.842029, 5.818673, 5.822323, 5.800344, 5.671194, 5.695325, 
    5.669767, 5.673203, 5.67166, 5.652951, 5.643541, 5.623865, 5.627433, 
    5.641886, 5.674748, 5.663575, 5.69176, 5.691122, 5.72262, 5.708403, 
    5.761531, 5.746394, 5.790213, 5.779171, 5.789694, 5.786501, 5.789735, 
    5.773547, 5.780479, 5.766248, 5.711063, 5.727243, 5.67909, 5.650283, 
    5.631203, 5.617695, 5.619603, 5.623242, 5.64197, 5.659618, 5.673096, 
    5.682124, 5.691031, 5.718058, 5.732395, 5.764597, 5.758774, 5.76864, 
    5.778073, 5.793938, 5.791325, 5.798323, 5.768377, 5.788268, 5.755459, 
    5.76442, 5.693462, 5.666587, 5.6552, 5.645241, 5.621071, 5.637754, 
    5.631173, 5.646837, 5.656808, 5.651875, 5.682371, 5.670501, 5.733246, 
    5.706157, 5.776972, 5.759968, 5.781053, 5.770286, 5.788743, 5.77213, 
    5.800928, 5.807213, 5.802918, 5.819428, 5.771211, 5.789695, 5.651737, 
    5.652542, 5.65629, 5.639829, 5.638822, 5.623768, 5.637161, 5.642872, 
    5.657386, 5.665986, 5.674169, 5.692192, 5.712371, 5.740674, 5.761069, 
    5.77477, 5.766366, 5.773786, 5.765492, 5.761607, 5.804858, 5.780544, 
    5.817051, 5.815026, 5.79849, 5.815255, 5.653106, 5.648478, 5.632434, 
    5.644987, 5.62213, 5.634917, 5.64228, 5.670751, 5.677018, 5.682837, 
    5.694341, 5.709129, 5.735141, 5.757843, 5.778622, 5.777097, 5.777634, 
    5.782283, 5.770772, 5.784174, 5.786427, 5.78054, 5.814755, 5.804965, 
    5.814983, 5.808608, 5.649982, 5.657773, 5.653562, 5.661482, 5.655902, 
    5.680747, 5.688211, 5.723233, 5.708838, 5.731757, 5.711163, 5.714808, 
    5.73251, 5.712274, 5.756591, 5.726521, 5.782464, 5.752342, 5.784356, 
    5.778532, 5.788176, 5.796824, 5.807716, 5.827854, 5.823185, 5.840054, 
    5.6694, 5.679533, 5.678638, 5.689254, 5.697114, 5.714177, 5.741623, 
    5.73129, 5.750268, 5.754084, 5.725255, 5.742945, 5.68632, 5.695442, 
    5.690008, 5.6702, 5.733673, 5.701034, 5.761407, 5.743647, 5.795591, 
    5.769718, 5.820617, 5.842479, 5.863099, 5.88727, 5.685066, 5.678175, 
    5.690516, 5.707627, 5.723532, 5.74473, 5.746901, 5.750879, 5.761193, 
    5.769876, 5.75214, 5.772055, 5.697563, 5.736511, 5.675573, 5.693875, 
    5.706617, 5.701023, 5.73011, 5.736981, 5.764968, 5.750487, 5.837079, 
    5.798655, 5.905715, 5.875659, 5.675769, 5.685042, 5.717402, 5.701988, 
    5.746146, 5.757054, 5.765931, 5.777296, 5.778522, 5.785264, 5.77422, 
    5.784827, 5.744774, 5.762648, 5.713694, 5.725582, 5.72011, 5.714114, 
    5.732635, 5.752419, 5.75284, 5.759194, 5.777134, 5.746325, 5.842057, 
    5.782806, 5.695166, 5.713084, 5.715643, 5.708695, 5.75596, 5.738801, 
    5.7851, 5.77256, 5.793115, 5.782895, 5.781392, 5.768286, 5.760138, 
    5.739588, 5.722907, 5.709702, 5.71277, 5.727282, 5.75363, 5.778635, 
    5.773151, 5.791551, 5.742936, 5.763287, 5.755415, 5.775954, 5.731017, 
    5.769276, 5.721268, 5.725465, 5.738461, 5.76467, 5.770476, 5.776686, 
    5.772853, 5.7543, 5.751263, 5.738144, 5.734528, 5.724551, 5.716301, 
    5.723839, 5.731763, 5.754306, 5.774679, 5.796948, 5.802406, 5.828527, 
    5.807261, 5.842389, 5.81252, 5.864291, 5.771494, 5.811637, 5.739052, 
    5.74684, 5.760948, 5.793393, 5.775858, 5.796368, 5.751143, 5.727785, 
    5.721748, 5.710505, 5.722006, 5.72107, 5.732089, 5.728546, 5.755056, 
    5.740805, 5.781355, 5.796205, 5.838285, 5.86419, 5.890639, 5.902343, 
    5.905909, 5.9074,
  8.093654, 8.12784, 8.121184, 8.148828, 8.133482, 8.151597, 8.100574, 
    8.129202, 8.110916, 8.096725, 8.202695, 8.150062, 8.257644, 8.223865, 
    8.308927, 8.252381, 8.320364, 8.307286, 8.346687, 8.335384, 8.385951, 
    8.351909, 8.412253, 8.37781, 8.383192, 8.350788, 8.160628, 8.196129, 
    8.158529, 8.163583, 8.161314, 8.133801, 8.119966, 8.091043, 8.096288, 
    8.117532, 8.165856, 8.149424, 8.190882, 8.189944, 8.236299, 8.215372, 
    8.293597, 8.271303, 8.335856, 8.319585, 8.335092, 8.330386, 8.335153, 
    8.311299, 8.321513, 8.300546, 8.219289, 8.243104, 8.172242, 8.129877, 
    8.101829, 8.081975, 8.08478, 8.090128, 8.117656, 8.143604, 8.163425, 
    8.176706, 8.189809, 8.229583, 8.25069, 8.298113, 8.289536, 8.304069, 
    8.317966, 8.341347, 8.337495, 8.347809, 8.303682, 8.33299, 8.284654, 
    8.297852, 8.193387, 8.153853, 8.137108, 8.122464, 8.086937, 8.111458, 
    8.101785, 8.124811, 8.139473, 8.132218, 8.17707, 8.15961, 8.251942, 
    8.212068, 8.316345, 8.291295, 8.322357, 8.306495, 8.333691, 8.309212, 
    8.351649, 8.360914, 8.354583, 8.378922, 8.307857, 8.335093, 8.132015, 
    8.133199, 8.138709, 8.114508, 8.113029, 8.0909, 8.110586, 8.118982, 
    8.140322, 8.152968, 8.165005, 8.191518, 8.221213, 8.26288, 8.292917, 
    8.313102, 8.300719, 8.31165, 8.299432, 8.29371, 8.357443, 8.321609, 
    8.375419, 8.372434, 8.348055, 8.372769, 8.134028, 8.127224, 8.103638, 
    8.122091, 8.088493, 8.107287, 8.118111, 8.159977, 8.169195, 8.177755, 
    8.194679, 8.216442, 8.254733, 8.288164, 8.318775, 8.316529, 8.31732, 
    8.324171, 8.307211, 8.326958, 8.330277, 8.321603, 8.372033, 8.357601, 
    8.37237, 8.362969, 8.129436, 8.14089, 8.134699, 8.146345, 8.13814, 
    8.17468, 8.185661, 8.237201, 8.216014, 8.24975, 8.219435, 8.224801, 
    8.250858, 8.22107, 8.286321, 8.242043, 8.324437, 8.280063, 8.327225, 
    8.318643, 8.332854, 8.3456, 8.361655, 8.391347, 8.384463, 8.40934, 
    8.15799, 8.172894, 8.171578, 8.187195, 8.198761, 8.223871, 8.264277, 
    8.249063, 8.277008, 8.282628, 8.240178, 8.266223, 8.182878, 8.196301, 
    8.188305, 8.159166, 8.25257, 8.204529, 8.293415, 8.267258, 8.343782, 
    8.305657, 8.380676, 8.412917, 8.443339, 8.479013, 8.181034, 8.170897, 
    8.189054, 8.214231, 8.237641, 8.268851, 8.272049, 8.277908, 8.293099, 
    8.305891, 8.279764, 8.3091, 8.199421, 8.25675, 8.167069, 8.193995, 
    8.212744, 8.204513, 8.247325, 8.257442, 8.29866, 8.277331, 8.404953, 
    8.348298, 8.506248, 8.461874, 8.167358, 8.180999, 8.228618, 8.205932, 
    8.270937, 8.287003, 8.300078, 8.316822, 8.318629, 8.328564, 8.312289, 
    8.32792, 8.268918, 8.295242, 8.22316, 8.24066, 8.232605, 8.223779, 
    8.251043, 8.280176, 8.280795, 8.290155, 8.316584, 8.271201, 8.412295, 
    8.324941, 8.195893, 8.222262, 8.226029, 8.215803, 8.285391, 8.260122, 
    8.328321, 8.309844, 8.340134, 8.325072, 8.322858, 8.303548, 8.291545, 
    8.26128, 8.236721, 8.217285, 8.221801, 8.243162, 8.28196, 8.318795, 
    8.310716, 8.337829, 8.26621, 8.296183, 8.284589, 8.314846, 8.24866, 
    8.305006, 8.234308, 8.240487, 8.259622, 8.298222, 8.306775, 8.315923, 
    8.310277, 8.282946, 8.278473, 8.259155, 8.25383, 8.239141, 8.226997, 
    8.238092, 8.249759, 8.282955, 8.312965, 8.345782, 8.353827, 8.392341, 
    8.360985, 8.412785, 8.368737, 8.445098, 8.308275, 8.367436, 8.260491, 
    8.271959, 8.292738, 8.340544, 8.314703, 8.344928, 8.278297, 8.243901, 
    8.235016, 8.218467, 8.235394, 8.234016, 8.250239, 8.245023, 8.28406, 
    8.263072, 8.322803, 8.344687, 8.406732, 8.44495, 8.483987, 8.501268, 
    8.506534, 8.508736,
  12.66504, 12.72051, 12.70971, 12.75458, 12.72967, 12.75908, 12.67627, 
    12.72272, 12.69304, 12.67002, 12.84208, 12.75658, 12.93144, 12.8765, 
    13.01492, 12.92288, 13.03355, 13.01225, 13.07645, 13.05803, 13.14047, 
    13.08496, 13.18338, 13.12719, 13.13597, 13.08313, 12.77374, 12.83141, 
    12.77033, 12.77854, 12.77485, 12.73018, 12.70773, 12.66081, 12.66931, 
    12.70378, 12.78223, 12.75555, 12.82289, 12.82136, 12.89672, 12.86269, 
    12.98996, 12.95367, 13.05879, 13.03228, 13.05755, 13.04988, 13.05765, 
    13.01879, 13.03542, 13.00127, 12.86906, 12.90779, 12.7926, 12.72381, 
    12.6783, 12.6461, 12.65065, 12.65932, 12.70398, 12.7461, 12.77828, 
    12.79986, 12.82114, 12.8858, 12.92013, 12.99731, 12.98335, 13.00701, 
    13.02965, 13.06774, 13.06146, 13.07827, 13.00638, 13.05412, 12.9754, 
    12.99689, 12.82696, 12.76274, 12.73555, 12.71178, 12.65415, 12.69392, 
    12.67823, 12.71559, 12.73939, 12.72761, 12.80045, 12.77209, 12.92216, 
    12.85732, 13.02701, 12.98621, 13.0368, 13.01096, 13.05526, 13.01539, 
    13.08453, 13.09964, 13.08932, 13.129, 13.01318, 13.05755, 12.72729, 
    12.72921, 12.73815, 12.69887, 12.69647, 12.66058, 12.69251, 12.70613, 
    12.74077, 12.7613, 12.78085, 12.82392, 12.87219, 12.93996, 12.98885, 
    13.02172, 13.00156, 13.01936, 12.99946, 12.99014, 13.09398, 13.03558, 
    13.12329, 13.11842, 13.07868, 13.11897, 12.73055, 12.71951, 12.68124, 
    12.71118, 12.65667, 12.68716, 12.70472, 12.77268, 12.78765, 12.80156, 
    12.82906, 12.86443, 12.92671, 12.98111, 13.03096, 13.02731, 13.02859, 
    13.03975, 13.01213, 13.0443, 13.0497, 13.03557, 13.11777, 13.09424, 
    13.11832, 13.10299, 12.7231, 12.74169, 12.73164, 12.75055, 12.73723, 
    12.79656, 12.8144, 12.89819, 12.86373, 12.9186, 12.8693, 12.87802, 
    12.9204, 12.87195, 12.97811, 12.90606, 13.04019, 12.96793, 13.04473, 
    13.03075, 13.0539, 13.07467, 13.10085, 13.14927, 13.13804, 13.17863, 
    12.76946, 12.79366, 12.79152, 12.8169, 12.83569, 12.87651, 12.94223, 
    12.91748, 12.96295, 12.9721, 12.90303, 12.9454, 12.80988, 12.83169, 
    12.8187, 12.77137, 12.92319, 12.84507, 12.98966, 12.94708, 13.07171, 
    13.0096, 13.13186, 13.18447, 13.23413, 13.29242, 12.80689, 12.79042, 
    12.81991, 12.86084, 12.8989, 12.94968, 12.95488, 12.96442, 12.98915, 
    13.00998, 12.96744, 13.0152, 12.83676, 12.92999, 12.7842, 12.82794, 
    12.85842, 12.84504, 12.91465, 12.93111, 12.9982, 12.96348, 13.17147, 
    13.07907, 13.33694, 13.26441, 12.78467, 12.80683, 12.88423, 12.84735, 
    12.95307, 12.97922, 13.00051, 13.02778, 13.03073, 13.04691, 13.0204, 
    13.04586, 12.94979, 12.99264, 12.87535, 12.90381, 12.89071, 12.87636, 
    12.9207, 12.96811, 12.96912, 12.98435, 13.02739, 12.9535, 13.18345, 
    13.04101, 12.83103, 12.87389, 12.88002, 12.86339, 12.9766, 12.93547, 
    13.04652, 13.01642, 13.06577, 13.04122, 13.03761, 13.00616, 12.98662, 
    12.93736, 12.8974, 12.8658, 12.87314, 12.90788, 12.97101, 13.031, 
    13.01784, 13.06201, 12.94538, 12.99417, 12.97529, 13.02456, 12.91683, 
    13.00854, 12.89348, 12.90353, 12.93466, 12.99749, 13.01142, 13.02632, 
    13.01712, 12.97262, 12.96534, 12.9339, 12.92524, 12.90134, 12.88159, 
    12.89964, 12.91861, 12.97263, 13.0215, 13.07497, 13.08809, 13.15089, 
    13.09975, 13.18425, 13.11239, 13.23701, 13.01386, 13.11027, 12.93608, 
    12.95474, 12.98856, 13.06643, 13.02433, 13.07358, 12.96505, 12.90908, 
    12.89463, 12.86772, 12.89525, 12.89301, 12.91939, 12.91091, 12.97443, 
    12.94027, 13.03753, 13.07319, 13.17437, 13.23676, 13.30054, 13.3288, 
    13.3374, 13.34101,
  20.59954, 20.69561, 20.67689, 20.75467, 20.71148, 20.76247, 20.61897, 
    20.69943, 20.64802, 20.60816, 20.90657, 20.75814, 21.06198, 20.96639, 
    21.20745, 21.04708, 21.23996, 21.2028, 21.31484, 21.28267, 21.42674, 
    21.3297, 21.50184, 21.40351, 21.41887, 21.32651, 20.78791, 20.88803, 
    20.782, 20.79624, 20.78984, 20.71237, 20.67346, 20.59221, 20.60693, 
    20.66662, 20.80264, 20.75635, 20.87322, 20.87057, 21.00156, 20.94239, 
    21.16393, 21.10069, 21.28401, 21.23774, 21.28184, 21.26846, 21.28201, 
    21.2142, 21.24322, 21.18365, 20.95345, 21.02082, 20.82064, 20.70133, 
    20.62249, 20.56676, 20.57463, 20.58964, 20.66697, 20.73996, 20.79579, 
    20.83323, 20.8702, 20.98256, 21.04229, 21.17675, 21.1524, 21.19366, 
    21.23314, 21.29964, 21.28868, 21.31803, 21.19256, 21.27586, 21.13855, 
    21.17601, 20.88029, 20.76882, 20.72168, 20.68049, 20.58068, 20.64955, 
    20.62237, 20.68709, 20.72833, 20.70792, 20.83426, 20.78504, 21.04584, 
    20.93305, 21.22853, 21.1574, 21.24562, 21.20055, 21.27785, 21.20827, 
    21.32897, 21.35536, 21.33732, 21.40669, 21.20442, 21.28184, 20.70735, 
    20.71068, 20.72619, 20.65812, 20.65396, 20.59181, 20.6471, 20.6707, 
    20.73072, 20.76633, 20.80024, 20.87502, 20.9589, 21.07682, 21.162, 
    21.21932, 21.18415, 21.21519, 21.18049, 21.16425, 21.34547, 21.2435, 
    21.3967, 21.38819, 21.31873, 21.38914, 20.71301, 20.69387, 20.62757, 
    20.67944, 20.58505, 20.63783, 20.66825, 20.78607, 20.81205, 20.83619, 
    20.88394, 20.94541, 21.05374, 21.14851, 21.23544, 21.22906, 21.23131, 
    21.25078, 21.20258, 21.25871, 21.26814, 21.24348, 21.38704, 21.34592, 
    21.388, 21.36121, 20.70009, 20.73232, 20.7149, 20.74768, 20.72458, 
    20.82752, 20.85849, 21.00411, 20.9442, 21.03963, 20.95387, 20.96904, 
    21.04277, 20.95849, 21.14328, 21.01781, 21.25154, 21.12553, 21.25946, 
    21.23507, 21.27547, 21.31174, 21.35747, 21.44214, 21.42249, 21.49352, 
    20.78048, 20.82248, 20.81877, 20.86282, 20.89546, 20.96641, 21.08078, 
    21.03769, 21.11687, 21.1328, 21.01254, 21.08629, 20.85064, 20.88852, 
    20.86595, 20.78379, 21.04762, 20.91175, 21.16341, 21.08922, 21.30657, 
    21.19817, 21.41169, 21.50374, 21.59075, 21.69298, 20.84544, 20.81685, 
    20.86806, 20.93916, 21.00536, 21.09374, 21.1028, 21.11942, 21.16252, 
    21.19884, 21.12468, 21.20795, 20.89733, 21.05945, 20.80606, 20.88201, 
    20.93496, 20.91171, 21.03276, 21.06142, 21.1783, 21.11778, 21.48098, 
    21.31942, 21.77116, 21.64383, 20.80688, 20.84534, 20.97983, 20.91571, 
    21.09965, 21.14521, 21.18233, 21.22989, 21.23503, 21.26327, 21.21701, 
    21.26144, 21.09393, 21.1686, 20.9644, 21.0139, 20.99111, 20.96615, 
    21.04329, 21.12585, 21.12761, 21.15416, 21.22921, 21.1004, 21.50196, 
    21.25297, 20.88737, 20.96186, 20.97251, 20.94361, 21.14064, 21.06901, 
    21.26258, 21.21006, 21.29619, 21.25334, 21.24705, 21.19218, 21.1581, 
    21.07229, 21.00275, 20.94779, 20.96056, 21.02098, 21.13091, 21.2355, 
    21.21254, 21.28963, 21.08626, 21.17127, 21.13837, 21.22427, 21.03654, 
    21.19632, 20.99593, 21.01341, 21.06759, 21.17706, 21.20135, 21.22733, 
    21.21129, 21.13371, 21.12102, 21.06627, 21.05118, 21.0096, 20.97525, 
    21.00664, 21.03966, 21.13373, 21.21893, 21.31226, 21.33517, 21.44497, 
    21.35555, 21.50336, 21.37765, 21.59578, 21.2056, 21.37394, 21.07005, 
    21.10255, 21.16149, 21.29735, 21.22387, 21.30983, 21.12052, 21.02307, 
    20.99793, 20.95113, 20.999, 20.9951, 21.04102, 21.02625, 21.13687, 
    21.07736, 21.24689, 21.30914, 21.48606, 21.59536, 21.70724, 21.75686, 
    21.77199, 21.77831,
  34.64163, 34.8224, 34.78714, 34.93374, 34.8523, 34.94846, 34.67816, 
    34.82961, 34.73281, 34.65783, 35.22083, 34.9403, 35.51565, 35.33417, 
    35.79265, 35.48733, 35.85468, 35.78377, 35.99778, 35.93627, 36.21213, 
    36.02621, 36.35634, 36.16759, 36.19703, 36.02011, 34.99647, 35.18573, 
    34.98531, 35.01219, 35.00012, 34.85399, 34.78069, 34.62785, 34.65553, 
    34.76781, 35.02429, 34.9369, 35.15771, 35.1527, 35.40089, 35.28867, 
    35.70966, 35.58926, 35.93884, 35.85044, 35.93468, 35.9091, 35.93501, 
    35.80551, 35.86091, 35.74726, 35.30965, 35.43745, 35.0583, 34.83319, 
    34.68478, 34.58004, 34.59482, 34.62303, 34.76847, 34.90601, 35.01135, 
    35.08208, 35.15198, 35.36484, 35.47823, 35.7341, 35.6877, 35.76633, 
    35.84167, 35.9687, 35.94775, 36.00388, 35.76424, 35.92325, 35.66132, 
    35.73268, 35.17108, 34.96045, 34.87153, 34.79392, 34.60619, 34.73568, 
    34.68455, 34.80635, 34.88408, 34.8456, 35.08402, 34.99105, 35.48497, 
    35.27098, 35.83287, 35.69722, 35.8655, 35.77948, 35.92706, 35.7942, 
    36.0248, 36.07532, 36.04079, 36.17368, 35.78685, 35.93468, 34.84452, 
    34.8508, 34.88002, 34.75181, 34.74398, 34.6271, 34.73107, 34.77549, 
    34.88858, 34.95574, 35.01976, 35.16111, 35.31997, 35.54385, 35.70599, 
    35.81528, 35.7482, 35.80742, 35.74123, 35.71027, 36.05639, 35.86143, 
    36.15452, 36.13821, 36.00522, 36.14004, 34.8552, 34.81913, 34.69434, 
    34.79195, 34.61441, 34.71363, 34.77087, 34.993, 35.04207, 35.08768, 
    35.17799, 35.2944, 35.49998, 35.68029, 35.84606, 35.83387, 35.83816, 
    35.87534, 35.78336, 35.89048, 35.90851, 35.8614, 36.13602, 36.05725, 
    36.13786, 36.08653, 34.83085, 34.89159, 34.85875, 34.92056, 34.877, 
    35.07129, 35.12984, 35.40573, 35.29211, 35.47318, 35.31043, 35.3392, 
    35.47914, 35.31919, 35.67033, 35.43174, 35.87679, 35.63653, 35.89193, 
    35.84534, 35.92252, 35.99186, 36.07936, 36.24167, 36.20399, 36.34034, 
    34.98244, 35.06177, 35.05476, 35.13803, 35.1998, 35.33421, 35.55138, 
    35.46948, 35.62004, 35.65038, 35.42173, 35.56187, 35.115, 35.18665, 
    35.14395, 34.98869, 35.48835, 35.23064, 35.70868, 35.56744, 35.98196, 
    35.77494, 36.18327, 36.35999, 36.52742, 36.72464, 35.10516, 35.05113, 
    35.14795, 35.28256, 35.4081, 35.57604, 35.59328, 35.6249, 35.70697, 
    35.77621, 35.63491, 35.79359, 35.20332, 35.51084, 35.03075, 35.17433, 
    35.2746, 35.23055, 35.46014, 35.51457, 35.73705, 35.62178, 36.31626, 
    36.00655, 36.87584, 36.62977, 35.03229, 35.10497, 35.35966, 35.23814, 
    35.58728, 35.67401, 35.74473, 35.83546, 35.84526, 35.8992, 35.81088, 
    35.8957, 35.5764, 35.71856, 35.3304, 35.42431, 35.38106, 35.33371, 
    35.48014, 35.63713, 35.64048, 35.69105, 35.83416, 35.58871, 36.35656, 
    35.87952, 35.18447, 35.32558, 35.34578, 35.29098, 35.6653, 35.529, 
    35.89788, 35.79763, 35.9621, 35.88023, 35.86821, 35.76352, 35.69856, 
    35.53524, 35.40316, 35.29892, 35.32311, 35.43776, 35.64677, 35.84616, 
    35.80235, 35.94957, 35.5618, 35.72365, 35.66097, 35.82474, 35.46732, 
    35.77141, 35.3902, 35.42338, 35.5263, 35.73468, 35.78099, 35.83058, 
    35.79997, 35.6521, 35.62794, 35.52379, 35.49512, 35.41615, 35.35098, 
    35.41052, 35.47322, 35.65215, 35.81455, 35.99285, 36.03667, 36.24712, 
    36.0757, 36.35925, 36.11801, 36.53712, 35.78912, 36.11091, 35.53099, 
    35.5928, 35.70501, 35.96433, 35.82397, 35.98819, 35.627, 35.44173, 
    35.394, 35.30524, 35.39603, 35.38864, 35.47581, 35.44776, 35.65811, 
    35.54489, 35.86792, 35.98689, 36.32602, 36.5363, 36.75221, 36.84815, 
    36.87743, 36.88968,
  60.67863, 61.07135, 60.99461, 61.31424, 61.13651, 61.34641, 60.75784, 
    61.08706, 60.87648, 60.71376, 61.94413, 61.32857, 62.59651, 62.19426, 
    63.21471, 62.5336, 63.35386, 63.19481, 63.67589, 63.5373, 64.16094, 
    63.74006, 64.48912, 64.05989, 64.12666, 63.72628, 61.45144, 61.86684, 
    61.42701, 61.48586, 61.45943, 61.14019, 60.98057, 60.6488, 60.70876, 
    60.95255, 61.51235, 61.32116, 61.80519, 61.79418, 62.34188, 62.09374, 
    63.02896, 62.76028, 63.54308, 63.34436, 63.53372, 63.47617, 63.53447, 
    63.24354, 63.36786, 63.11306, 62.14007, 62.4229, 61.58688, 61.09486, 
    60.77221, 60.5453, 60.57728, 60.63834, 60.95398, 61.25367, 61.48402, 
    61.63907, 61.79259, 62.26209, 62.51339, 63.0836, 62.97988, 63.15576, 
    63.32466, 63.61035, 63.56314, 63.68966, 63.15108, 63.508, 62.92097, 
    63.08044, 61.83461, 61.37262, 61.17844, 61.00935, 60.60189, 60.88271, 
    60.77171, 61.03641, 61.20581, 61.12191, 61.64332, 61.43957, 62.52835, 
    62.0547, 63.30491, 63.00114, 63.37816, 63.1852, 63.51657, 63.21818, 
    63.73687, 63.85098, 63.77296, 64.07369, 63.20173, 63.53373, 61.11956, 
    61.13323, 61.19697, 60.91776, 60.90075, 60.64716, 60.87269, 60.96924, 
    61.21564, 61.36234, 61.50242, 61.81266, 62.16286, 62.65922, 63.02074, 
    63.26545, 63.11516, 63.24781, 63.09957, 63.03032, 63.80819, 63.36903, 
    64.03026, 63.9933, 63.69268, 63.99746, 61.14283, 61.06424, 60.79295, 
    61.00505, 60.61967, 60.83482, 60.95921, 61.44385, 61.55131, 61.65134, 
    61.8498, 62.1064, 62.5617, 62.96332, 63.33451, 63.30716, 63.31678, 
    63.40028, 63.19389, 63.43429, 63.47484, 63.36896, 63.98835, 63.81014, 
    63.99251, 63.87634, 61.08976, 61.22222, 61.15057, 61.28544, 61.19038, 
    61.61537, 61.74393, 62.35262, 62.10133, 62.50217, 62.1418, 62.20536, 
    62.5154, 62.16116, 62.94107, 62.41025, 63.40353, 62.86564, 63.43755, 
    63.33289, 63.50635, 63.66254, 63.86012, 64.22806, 64.14246, 64.45264, 
    61.42073, 61.5945, 61.57913, 61.76192, 61.8978, 62.19434, 62.67596, 
    62.49397, 62.82887, 62.89655, 62.38805, 62.6993, 61.71132, 61.86886, 
    61.77494, 61.43441, 62.53585, 61.96574, 63.02676, 62.71171, 63.64022, 
    63.17503, 64.09545, 64.49744, 64.88042, 65.33417, 61.68972, 61.57118, 
    61.78372, 62.08025, 62.35786, 62.73084, 62.76924, 62.83971, 63.02295, 
    63.17787, 62.86205, 63.21682, 61.90557, 62.58582, 61.5265, 61.84175, 
    62.06268, 61.96555, 62.47323, 62.59411, 63.09022, 62.83276, 64.39777, 
    63.69567, 65.68402, 65.11553, 61.52988, 61.6893, 62.25063, 61.98228, 
    62.75588, 62.9493, 63.1074, 63.31071, 63.33273, 63.4539, 63.25558, 
    63.44603, 62.73164, 63.04886, 62.18592, 62.39378, 62.29797, 62.19324, 
    62.51762, 62.867, 62.87447, 62.98737, 63.30781, 62.75906, 64.48964, 
    63.40967, 61.86407, 62.17528, 62.21993, 62.09884, 62.92986, 62.62619, 
    63.45094, 63.22586, 63.59548, 63.41127, 63.38426, 63.14944, 63.00415, 
    62.64006, 62.34691, 62.11637, 62.16982, 62.42359, 62.88849, 63.33474, 
    63.23645, 63.56723, 62.69914, 63.06023, 62.92019, 63.28667, 62.48916, 
    63.16713, 62.31822, 62.39172, 62.62019, 63.08491, 63.1886, 63.29978, 
    63.23112, 62.90038, 62.8465, 62.6146, 62.5509, 62.3757, 62.23141, 
    62.36323, 62.50227, 62.90049, 63.26381, 63.66477, 63.76367, 64.24043, 
    63.85184, 64.49577, 63.94757, 64.90266, 63.2068, 63.9315, 62.63061, 
    62.76817, 63.01857, 63.60049, 63.28493, 63.65427, 62.84439, 62.4324, 
    62.32663, 62.13035, 62.33114, 62.31475, 62.50801, 62.44577, 62.9138, 
    62.66153, 63.38359, 63.65133, 64.42001, 64.90079, 65.39783, 65.61983, 
    65.68771, 65.71613,
  116.3177, 117.5456, 117.3041, 118.3152, 117.7513, 118.4177, 116.5638, 
    117.5952, 116.9339, 116.4268, 120.3482, 118.3608, 122.5137, 121.171, 
    124.6258, 122.3021, 125.1096, 124.5568, 126.2418, 125.7524, 127.9808, 
    126.4695, 129.1813, 127.6151, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9487, 118.3372, 119.895, 119.8592, 121.661, 120.8393, 
    123.9848, 123.0674, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7258, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9053, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3958, 122.2342, 124.1728, 123.8164, 124.4217, 
    125.0078, 126.0099, 125.8434, 126.2906, 124.4056, 125.6494, 123.6147, 
    124.1619, 119.9907, 118.5013, 117.8839, 117.3505, 116.0801, 116.9533, 
    116.607, 117.4356, 117.9707, 117.7052, 119.3704, 118.7153, 122.2845, 
    120.7108, 124.9391, 123.8893, 125.1945, 124.5236, 125.6795, 124.6378, 
    126.4581, 126.8648, 126.5865, 127.6649, 124.5808, 125.7399, 117.6978, 
    117.741, 117.9427, 117.063, 117.0098, 116.2202, 116.922, 117.2245, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9566, 
    124.8018, 124.2816, 124.7406, 124.2278, 123.9895, 126.712, 125.1626, 
    127.5082, 127.3751, 126.3013, 127.39, 117.7713, 117.5232, 116.6731, 
    117.337, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.881, 122.3965, 123.7596, 125.0421, 124.9469, 124.9804, 
    125.2718, 124.5536, 125.3908, 125.5329, 125.1623, 127.3573, 126.719, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9218, 
    119.2802, 119.696, 121.6967, 120.8643, 122.1966, 120.9977, 121.2078, 
    122.241, 121.0616, 123.6834, 121.889, 125.2831, 123.4258, 125.4022, 
    125.0365, 125.6436, 126.1945, 126.8974, 128.2247, 127.9138, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1968, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8149, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3097, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4884, 127.7436, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7949, 121.7142, 122.9675, 123.0978, 123.3374, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.014, 
    120.7371, 120.4183, 122.0996, 122.5056, 124.1956, 123.3137, 128.8452, 
    126.3119, 133.7281, 131.5293, 119.005, 119.5191, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2548, 124.9593, 125.0359, 125.4595, 124.7676, 
    125.4319, 122.9702, 124.0532, 121.1435, 121.834, 121.5149, 121.1677, 
    122.2484, 123.4304, 123.4559, 123.842, 124.9492, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1083, 121.256, 120.8561, 123.6451, 122.6137, 
    125.4491, 124.6644, 125.9575, 125.3102, 125.2158, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.043, 
    124.7011, 125.8578, 122.8602, 124.0923, 123.612, 124.8756, 122.153, 
    124.4611, 121.5822, 121.8271, 122.5935, 124.1773, 124.5353, 124.9212, 
    124.6827, 123.5443, 123.3605, 122.5747, 122.3602, 121.7737, 121.294, 
    121.7321, 122.197, 123.5447, 124.7961, 126.2024, 126.5535, 128.2698, 
    126.8678, 129.2059, 127.2107, 130.7229, 124.5984, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9752, 124.8696, 126.1652, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5902, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6129, 133.4765, 
    133.7426, 133.8544,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02029252, -0.01996136, -0.02002529, -0.0197615, -0.01990738, 
    -0.01973531, -0.02022492, -0.01994832, -0.02012443, -0.02026249, 
    -0.01926015, -0.01974982, -0.01876547, -0.01906761, -0.01831844, 
    -0.01881213, -0.01822061, -0.01833252, -0.017998, -0.01809316, 
    -0.01767244, -0.01795427, -0.01745858, -0.01773932, -0.01769507, 
    -0.01796365, -0.01965025, -0.01932038, -0.01966997, -0.01962252, 
    -0.0196438, -0.01990434, -0.02003702, -0.02031809, -0.02026676, 
    -0.02006048, -0.01960122, -0.01975586, -0.01936868, -0.01937734, 
    -0.01895567, -0.01914455, -0.01845061, -0.01864504, -0.01808918, 
    -0.01822726, -0.01809563, -0.01813544, -0.01809511, -0.01829809, 
    -0.01821082, -0.01839055, -0.01910901, -0.01889476, -0.01954154, 
    -0.01994185, -0.0202127, -0.02040726, -0.02037963, -0.02032707, 
    -0.02005928, -0.019811, -0.01962399, -0.01949996, -0.01937858, 
    -0.01901602, -0.01882716, -0.01841154, -0.01848584, -0.01836019, 
    -0.01824106, -0.01804288, -0.01807534, -0.0179886, -0.01836351, 
    -0.0181134, -0.0185283, -0.0184138, -0.0193456, -0.01971402, -0.01987278, 
    -0.02001298, -0.02035842, -0.02011918, -0.02021312, -0.01999042, 
    -0.01985027, -0.01991946, -0.01949658, -0.01965982, -0.01881603, 
    -0.01917459, -0.01825491, -0.01847056, -0.01820363, -0.01833932, 
    -0.01810748, -0.01831599, -0.01795644, -0.01787915, -0.01793193, 
    -0.01773016, -0.01832762, -0.01809562, -0.01992139, -0.01991009, 
    -0.01985753, -0.02008968, -0.02010399, -0.0203195, -0.02012762, 
    -0.0200465, -0.01984219, -0.01972236, -0.01960919, -0.01936282, 
    -0.01909158, -0.01871918, -0.0184565, -0.01828265, -0.01838905, 
    -0.01829508, -0.01840016, -0.01844964, -0.01790806, -0.01821, 
    -0.01775902, -0.01778366, -0.01798654, -0.01778089, -0.01990216, 
    -0.01996727, -0.02019508, -0.02001656, -0.02034312, -0.02015961, 
    -0.0200549, -0.01965637, -0.01956998, -0.01949021, -0.01933371, 
    -0.01913483, -0.01879126, -0.01849775, -0.01823416, -0.01825333, 
    -0.01824658, -0.0181882, -0.01833317, -0.01816452, -0.01813637, 
    -0.01821005, -0.01778697, -0.01790674, -0.01778419, -0.01786207, 
    -0.01994608, -0.01983678, -0.01989576, -0.01978501, -0.01986296, 
    -0.01951882, -0.0194169, -0.01894758, -0.01913872, -0.01883551, 
    -0.01910769, -0.01905915, -0.01882566, -0.01909288, -0.01851378, 
    -0.01890424, -0.01818593, -0.01856833, -0.01816225, -0.01823529, 
    -0.01811454, -0.01800713, -0.01787299, -0.01762829, -0.01768463, 
    -0.0174821, -0.01967505, -0.01953546, -0.01954773, -0.01940272, 
    -0.01929621, -0.01906755, -0.01870686, -0.01884163, -0.01859504, 
    -0.01854595, -0.01892091, -0.01868971, -0.01944266, -0.0193188, 
    -0.01939246, -0.01966398, -0.01881045, -0.01924337, -0.01845219, 
    -0.01868061, -0.0180224, -0.01834652, -0.01771573, -0.01745322, 
    -0.01721011, -0.01693054, -0.01945976, -0.01955409, -0.01938556, 
    -0.01915492, -0.01894363, -0.01866658, -0.0186385, -0.01858716, 
    -0.01845492, -0.01834451, -0.01857094, -0.01831695, -0.01929016, 
    -0.01877338, -0.01958986, -0.01934001, -0.01916844, -0.01924352, 
    -0.0188571, -0.01876725, -0.01840682, -0.01859221, -0.0175176, 
    -0.0179845, -0.01672105, -0.01706412, -0.01958716, -0.01946009, 
    -0.01902472, -0.01923055, -0.01864826, -0.01850786, -0.01839458, 
    -0.01825083, -0.0182354, -0.01815089, -0.0182896, -0.01815636, -0.018666, 
    -0.01843636, -0.01907397, -0.01891661, -0.01898883, -0.01906838, 
    -0.01882401, -0.01856734, -0.01856194, -0.01848046, -0.01825287, 
    -0.01864594, -0.01745824, -0.01818165, -0.01932255, -0.01908209, 
    -0.01904806, -0.01914063, -0.01852188, -0.01874354, -0.01815295, 
    -0.01831056, -0.0180531, -0.01818054, -0.01819937, -0.01836468, 
    -0.0184684, -0.01873331, -0.01895188, -0.01912718, -0.01908626, 
    -0.01889424, -0.01855178, -0.01823399, -0.01830309, -0.01807253, 
    -0.01868983, -0.01842823, -0.01852885, -0.01826772, -0.01884522, 
    -0.01835212, -0.01897353, -0.01891815, -0.01874797, -0.01841061, 
    -0.01833691, -0.01825851, -0.01830685, -0.01854318, -0.01858222, 
    -0.01875209, -0.01879927, -0.0189302, -0.01903932, -0.01893958, 
    -0.01883544, -0.01854309, -0.01828381, -0.0180056, -0.01793823, 
    -0.01762017, -0.01787857, -0.01745429, -0.01781423, -0.01719618, 
    -0.01832403, -0.01782501, -0.01874027, -0.01863928, -0.01845806, 
    -0.01804965, -0.01826894, -0.01801278, -0.01858376, -0.01888764, 
    -0.01896717, -0.01911647, -0.01896377, -0.01897615, -0.01883117, 
    -0.01887763, -0.01853347, -0.01871749, -0.01819983, -0.01801479, 
    -0.01750319, -0.01719736, -0.01689203, -0.0167591, -0.01671887, 
    -0.01670208,
  -0.05426379, -0.05321441, -0.05341675, -0.05258257, -0.05304364, 
    -0.05249986, -0.05404934, -0.05317315, -0.05373077, -0.0541685, 
    -0.05100255, -0.05254569, -0.04945065, -0.05039767, -0.0480544, 
    -0.04959671, -0.04774964, -0.04809828, -0.04705726, -0.04735304, 
    -0.04604734, -0.04692141, -0.04538573, -0.04625455, -0.04611744, 
    -0.04695052, -0.05223133, -0.051192, -0.05229358, -0.05214384, -0.052211, 
    -0.05303403, -0.0534539, -0.05434496, -0.05418205, -0.05352819, 
    -0.05207666, -0.05256475, -0.05134399, -0.05137123, -0.05004649, 
    -0.05063926, -0.0484666, -0.04907392, -0.04734065, -0.04777034, 
    -0.04736073, -0.04748455, -0.04735912, -0.04799099, -0.04771917, 
    -0.04827922, -0.05052766, -0.04985555, -0.05188849, -0.05315268, 
    -0.05401057, -0.0546281, -0.05454034, -0.05437345, -0.05352439, 
    -0.05273894, -0.0521485, -0.05175743, -0.05137514, -0.05023577, 
    -0.04964379, -0.04834472, -0.04857656, -0.04818456, -0.04781332, 
    -0.04719672, -0.04729764, -0.04702803, -0.04819492, -0.047416, 
    -0.04870912, -0.04835176, -0.05127136, -0.05243262, -0.05293425, 
    -0.05337778, -0.05447297, -0.05371413, -0.05401192, -0.05330637, 
    -0.05286306, -0.05308184, -0.05174678, -0.05226154, -0.04960894, 
    -0.05073364, -0.04785646, -0.04852889, -0.04769678, -0.0481195, 
    -0.04739757, -0.04804678, -0.04692814, -0.0466882, -0.04685202, 
    -0.04622615, -0.04808303, -0.0473607, -0.05308797, -0.05305222, 
    -0.05288602, -0.05362068, -0.05366599, -0.05434942, -0.05374089, 
    -0.05348391, -0.05283751, -0.05245898, -0.05210182, -0.05132554, 
    -0.05047292, -0.0493058, -0.04848499, -0.04794288, -0.04827455, 
    -0.0479816, -0.0483092, -0.04846357, -0.04677793, -0.04771662, 
    -0.04631562, -0.046392, -0.04702163, -0.04638339, -0.05302713, 
    -0.05323311, -0.05395472, -0.05338913, -0.0544244, -0.05384227, 
    -0.05351051, -0.05225065, -0.05197815, -0.0517267, -0.05123393, 
    -0.05060874, -0.04953137, -0.04861375, -0.04779183, -0.04785156, 
    -0.04783052, -0.04764874, -0.04810032, -0.04757503, -0.04748743, 
    -0.04771678, -0.04640224, -0.04677384, -0.04639363, -0.04663518, 
    -0.05316608, -0.05282044, -0.05300691, -0.05265682, -0.05290318, 
    -0.05181687, -0.05149578, -0.05002112, -0.05062094, -0.04966995, 
    -0.0505235, -0.05037111, -0.0496391, -0.050477, -0.04866381, -0.04988529, 
    -0.04764168, -0.04883418, -0.04756798, -0.04779536, -0.04741956, 
    -0.04708561, -0.04666908, -0.04591065, -0.04608512, -0.04545843, 
    -0.0523096, -0.05186933, -0.051908, -0.05145113, -0.05111596, 
    -0.05039748, -0.04926725, -0.04968911, -0.04891762, -0.04876425, 
    -0.04993753, -0.0492136, -0.05157691, -0.05118703, -0.05141884, 
    -0.05227469, -0.04959146, -0.0509498, -0.04847154, -0.04918513, 
    -0.04713306, -0.04814195, -0.04618145, -0.04536917, -0.04461884, 
    -0.04375831, -0.05163077, -0.05192804, -0.0513971, -0.05067182, 
    -0.05000874, -0.04914127, -0.04905346, -0.048893, -0.04848006, 
    -0.04813568, -0.04884233, -0.04804976, -0.05109692, -0.04947541, 
    -0.05204083, -0.05125377, -0.05071431, -0.05095028, -0.04973758, 
    -0.04945621, -0.04832999, -0.04890879, -0.04556818, -0.0470153, 
    -0.04311513, -0.04416917, -0.05203231, -0.05163182, -0.05026307, 
    -0.05090949, -0.04908397, -0.0486453, -0.0482918, -0.04784377, 
    -0.04779572, -0.04753263, -0.04796454, -0.04754964, -0.04913944, 
    -0.04842215, -0.05041764, -0.04992404, -0.0501505, -0.05040011, 
    -0.04963394, -0.0488311, -0.0488142, -0.04855976, -0.04785011, 
    -0.04907672, -0.04538468, -0.04762835, -0.05119881, -0.05044314, 
    -0.05033631, -0.05062695, -0.04868908, -0.049382, -0.04753904, 
    -0.04802985, -0.04722847, -0.0476249, -0.04768351, -0.04819854, 
    -0.04852214, -0.04934999, -0.05003461, -0.0505847, -0.05045623, 
    -0.04985394, -0.04878246, -0.04779132, -0.04800658, -0.04728888, 
    -0.04921398, -0.04839677, -0.04871087, -0.04789638, -0.04970035, 
    -0.0481594, -0.05010249, -0.04992888, -0.04939587, -0.0483418, 
    -0.04811199, -0.04786769, -0.0480183, -0.0487556, -0.04887758, 
    -0.04940877, -0.04955646, -0.04996664, -0.05030889, -0.04999606, 
    -0.04966972, -0.04875533, -0.0479465, -0.04708086, -0.04687159, 
    -0.04588552, -0.04668639, -0.04537248, -0.04648679, -0.04457592, 
    -0.04807183, -0.04652021, -0.04937179, -0.0490559, -0.04848985, 
    -0.04721776, -0.04790018, -0.04710316, -0.04888237, -0.04983324, 
    -0.05008257, -0.05055105, -0.05007191, -0.05011071, -0.04965634, 
    -0.04980188, -0.04872528, -0.04930049, -0.04768496, -0.04710943, 
    -0.04552364, -0.04457953, -0.04363998, -0.04323184, -0.04310844, 
    -0.04305696,
  -0.07890929, -0.07725387, -0.07757289, -0.07625824, -0.07698469, 
    -0.07612797, -0.0785708, -0.07718883, -0.07806816, -0.07875887, 
    -0.07377228, -0.07620016, -0.07133588, -0.07282201, -0.06914855, 
    -0.07156496, -0.0686717, -0.06921722, -0.06758921, -0.0680515, 
    -0.06601233, -0.06737695, -0.06498064, -0.06633567, -0.0661217, 
    -0.06742244, -0.07570515, -0.07407007, -0.07580315, -0.07556741, 
    -0.07567313, -0.07696956, -0.07763146, -0.07903743, -0.07878026, 
    -0.07774863, -0.07546166, -0.07623018, -0.07430902, -0.07435185, 
    -0.07227068, -0.07320144, -0.06979382, -0.07074527, -0.06803215, 
    -0.0687041, -0.06806353, -0.06825712, -0.06806101, -0.06904931, 
    -0.06862404, -0.06950043, -0.07302615, -0.07197104, -0.07516553, 
    -0.07715657, -0.07850962, -0.07948453, -0.07934594, -0.07908241, 
    -0.07774263, -0.07650457, -0.07557476, -0.07495931, -0.07435801, 
    -0.07256781, -0.07163882, -0.06960297, -0.06996602, -0.06935225, 
    -0.06877133, -0.06780717, -0.06796491, -0.06754355, -0.06936847, 
    -0.06814995, -0.07017367, -0.06961401, -0.07419483, -0.07602207, 
    -0.0768123, -0.07751144, -0.07923955, -0.0780419, -0.07851176, 
    -0.07739885, -0.07670012, -0.0770449, -0.07494255, -0.07575271, 
    -0.07158414, -0.07334971, -0.06883882, -0.06989136, -0.06858902, 
    -0.06925042, -0.06812113, -0.06913661, -0.06738747, -0.06701268, 
    -0.06726855, -0.06629134, -0.06919335, -0.06806348, -0.07705456, 
    -0.07699821, -0.0767363, -0.07789449, -0.07796597, -0.07904446, 
    -0.07808412, -0.0776788, -0.07665987, -0.07606359, -0.07550126, 
    -0.07428001, -0.07294019, -0.07110875, -0.06982262, -0.06897403, 
    -0.06949313, -0.06903462, -0.06954737, -0.06978907, -0.06715282, 
    -0.06862006, -0.06643098, -0.0665502, -0.06753355, -0.06653676, 
    -0.07695867, -0.07728335, -0.0784215, -0.07752933, -0.07916285, 
    -0.07824406, -0.07772073, -0.07573555, -0.07530662, -0.07491096, 
    -0.07413598, -0.0731535, -0.07146247, -0.07002427, -0.06873771, 
    -0.06883115, -0.06879823, -0.06851388, -0.06922041, -0.06839861, 
    -0.06826163, -0.0686203, -0.06656619, -0.06714643, -0.06655274, 
    -0.06692988, -0.07717767, -0.07663297, -0.0769268, -0.0763752, 
    -0.07676333, -0.07505284, -0.07454773, -0.07223085, -0.07317267, 
    -0.07167985, -0.07301962, -0.0727803, -0.07163145, -0.07294659, 
    -0.07010268, -0.0720177, -0.06850285, -0.07036958, -0.06838759, 
    -0.06874322, -0.0681555, -0.06763351, -0.06698282, -0.06579909, 
    -0.06607127, -0.06509395, -0.07582837, -0.07513537, -0.07519623, 
    -0.0744775, -0.07395053, -0.07282171, -0.07104832, -0.0717099, 
    -0.07050031, -0.07026002, -0.07209968, -0.07096421, -0.07467533, 
    -0.07406225, -0.07442673, -0.0757734, -0.07155673, -0.07368937, 
    -0.06980155, -0.07091958, -0.06770767, -0.06928556, -0.06622158, 
    -0.06495484, -0.06378614, -0.06244756, -0.07476005, -0.07522776, 
    -0.07439254, -0.0732526, -0.07221144, -0.07085083, -0.07071319, 
    -0.07046175, -0.06981489, -0.06927574, -0.07038234, -0.06914128, 
    -0.0739206, -0.07137471, -0.07540528, -0.07416717, -0.07331934, 
    -0.07369012, -0.07178595, -0.0713446, -0.06957991, -0.07048648, 
    -0.06526504, -0.06752365, -0.06144832, -0.06308643, -0.07539187, 
    -0.0747617, -0.07261066, -0.07362602, -0.07076102, -0.07007368, 
    -0.06952012, -0.06881896, -0.06874379, -0.06833231, -0.06900793, 
    -0.0683589, -0.07084797, -0.06972422, -0.07285337, -0.0720785, 
    -0.07243394, -0.07282583, -0.07162336, -0.07036475, -0.07033828, 
    -0.06993972, -0.06882888, -0.07074965, -0.06497901, -0.06848201, 
    -0.07408077, -0.07289341, -0.07272565, -0.07318211, -0.07014227, 
    -0.07122824, -0.06834233, -0.06911013, -0.06785679, -0.06847659, 
    -0.06856827, -0.06937414, -0.06988078, -0.07117804, -0.07225204, 
    -0.07311574, -0.07291397, -0.07196851, -0.07028855, -0.0687369, 
    -0.06907371, -0.0679512, -0.0709648, -0.06968448, -0.0701764, 
    -0.06890127, -0.07172753, -0.06931288, -0.07235859, -0.0720861, 
    -0.07124998, -0.0695984, -0.06923866, -0.06885639, -0.06909205, 
    -0.07024647, -0.07043758, -0.07127022, -0.07150183, -0.07214535, 
    -0.0726826, -0.07219153, -0.0716795, -0.07024605, -0.06897969, 
    -0.06762609, -0.06729913, -0.0657599, -0.06700986, -0.06496, -0.06669819, 
    -0.06371935, -0.06917582, -0.06675036, -0.07121223, -0.07071703, 
    -0.06983023, -0.06784004, -0.06890722, -0.06766095, -0.07044509, 
    -0.07193603, -0.07232731, -0.0730629, -0.07231058, -0.07237148, 
    -0.07165849, -0.07188682, -0.07019898, -0.07110044, -0.06857054, 
    -0.06767074, -0.06519561, -0.06372496, -0.06226364, -0.06162957, 
    -0.06143793, -0.061358,
  -0.08616409, -0.08425445, -0.08462235, -0.08310658, -0.08394406, 
    -0.08295643, -0.08577351, -0.08417945, -0.08519361, -0.08599051, 
    -0.08024279, -0.08303963, -0.07743932, -0.07914896, -0.0749253, 
    -0.07770278, -0.0743776, -0.07500418, -0.07313477, -0.07366545, 
    -0.0713256, -0.07289115, -0.07014277, -0.07169645, -0.07145105, 
    -0.07294336, -0.08246914, -0.08058567, -0.08258208, -0.08231043, 
    -0.08243226, -0.0839266, -0.0846899, -0.08631197, -0.0860152, 
    -0.08482504, -0.08218858, -0.08307423, -0.08086082, -0.08091015, 
    -0.07851456, -0.07958565, -0.07566666, -0.07676022, -0.07364323, 
    -0.0744148, -0.07367926, -0.07390153, -0.07367637, -0.07481129, 
    -0.07432287, -0.07532955, -0.07938389, -0.07816985, -0.08184738, 
    -0.08414225, -0.08570292, -0.08682799, -0.08666803, -0.08636389, 
    -0.08481812, -0.08339052, -0.08231889, -0.08160982, -0.08091724, 
    -0.07885645, -0.07778772, -0.07544737, -0.07586454, -0.07515931, 
    -0.07449201, -0.07338496, -0.07356604, -0.07308237, -0.07517795, 
    -0.07377847, -0.07610317, -0.07546004, -0.08072933, -0.08283439, 
    -0.0837453, -0.08455148, -0.08654524, -0.08516333, -0.08570538, 
    -0.08442163, -0.08361597, -0.08401348, -0.08159052, -0.08252395, 
    -0.07772484, -0.07975632, -0.07456953, -0.07577874, -0.07428265, 
    -0.07504231, -0.07374538, -0.07491158, -0.07290322, -0.07247313, 
    -0.07276675, -0.0716456, -0.07497676, -0.0736792, -0.08402462, 
    -0.08395965, -0.08365767, -0.0849933, -0.08507573, -0.08632009, 
    -0.08521203, -0.0847445, -0.08356956, -0.08288223, -0.08223421, 
    -0.08082741, -0.07928496, -0.07717814, -0.07569975, -0.07472483, 
    -0.07532116, -0.07479443, -0.07538348, -0.0756612, -0.07263394, 
    -0.0743183, -0.07180577, -0.07194254, -0.07307088, -0.07192712, 
    -0.08391406, -0.08428844, -0.08560124, -0.08457211, -0.08645672, 
    -0.08539654, -0.08479287, -0.08250419, -0.08200995, -0.08155413, 
    -0.08066156, -0.07953046, -0.07758491, -0.07593148, -0.07445341, 
    -0.07456072, -0.07452291, -0.07419635, -0.07500784, -0.07406399, 
    -0.0739067, -0.07431857, -0.07196087, -0.07262661, -0.07194545, 
    -0.07237813, -0.08416658, -0.08353855, -0.08387731, -0.0832414, 
    -0.08368884, -0.08171756, -0.08113575, -0.07846875, -0.07955254, 
    -0.0778349, -0.07937638, -0.07910096, -0.07777925, -0.07929233, 
    -0.07602159, -0.07822353, -0.07418369, -0.07632836, -0.07405134, 
    -0.07445973, -0.07378485, -0.07318562, -0.07243887, -0.07108106, 
    -0.0713932, -0.07027265, -0.08261115, -0.08181264, -0.08188275, 
    -0.08105486, -0.08044801, -0.07914861, -0.07710864, -0.07786947, 
    -0.07647863, -0.07620243, -0.07831784, -0.07701194, -0.08128271, 
    -0.08057666, -0.08099638, -0.0825478, -0.07769331, -0.08014733, 
    -0.07567553, -0.07696062, -0.07327075, -0.07508269, -0.07156559, 
    -0.0701132, -0.06877412, -0.0672415, -0.08138029, -0.08191908, -0.080957, 
    -0.07964454, -0.0784464, -0.07688159, -0.07672334, -0.0764343, 
    -0.07569087, -0.07507141, -0.07634302, -0.07491694, -0.08041356, 
    -0.07748398, -0.08212361, -0.08069747, -0.07972136, -0.08014819, 
    -0.07795694, -0.07744934, -0.07542087, -0.07646272, -0.07046876, 
    -0.07305952, -0.06609818, -0.06797283, -0.08210815, -0.0813822, 
    -0.07890575, -0.08007439, -0.07677832, -0.07598826, -0.07535218, 
    -0.07454673, -0.07446038, -0.07398786, -0.07476376, -0.07401839, 
    -0.07687829, -0.07558668, -0.07918505, -0.07829347, -0.07870241, 
    -0.07915335, -0.07776993, -0.07632281, -0.07629238, -0.07583431, 
    -0.07455812, -0.07676526, -0.07014091, -0.07415976, -0.08059797, 
    -0.07923113, -0.07903807, -0.07956339, -0.07606709, -0.07731554, 
    -0.07399936, -0.07488116, -0.07344192, -0.07415354, -0.07425882, 
    -0.07518446, -0.07576659, -0.07725781, -0.07849312, -0.079487, 
    -0.07925478, -0.07816694, -0.07623523, -0.07445248, -0.07483932, 
    -0.07355031, -0.07701262, -0.07554101, -0.07610632, -0.07464126, 
    -0.07788975, -0.07511408, -0.0786157, -0.07830222, -0.07734054, 
    -0.07544211, -0.07502881, -0.07458971, -0.07486039, -0.07618686, 
    -0.07640652, -0.07736381, -0.07763016, -0.07837038, -0.07898852, 
    -0.07842351, -0.0778345, -0.07618637, -0.07473133, -0.0731771, 
    -0.07280184, -0.07103613, -0.07246991, -0.07011912, -0.07211231, 
    -0.06869762, -0.07495663, -0.07217216, -0.07729713, -0.07672776, 
    -0.07570849, -0.07342269, -0.07464808, -0.07321712, -0.07641515, 
    -0.07812958, -0.07857972, -0.07942618, -0.07856047, -0.07863053, 
    -0.07781034, -0.07807297, -0.07613226, -0.07716858, -0.07426142, 
    -0.07322835, -0.07038917, -0.06870405, -0.067031, -0.06630552, 
    -0.06608631, -0.06599487,
  -0.06725447, -0.06570853, -0.06600637, -0.06477926, -0.06545725, 
    -0.0646577, -0.06693828, -0.06564782, -0.06646883, -0.06711395, 
    -0.06246073, -0.06472506, -0.06019095, -0.06157513, -0.05815549, 
    -0.06040426, -0.05771205, -0.05821935, -0.05670581, -0.05713546, 
    -0.05524106, -0.05650856, -0.05428343, -0.0555413, -0.05534261, 
    -0.05655083, -0.06426319, -0.06273833, -0.06435462, -0.0641347, 
    -0.06423333, -0.06544312, -0.06606106, -0.06737418, -0.06713394, 
    -0.06617046, -0.06403605, -0.06475306, -0.06296109, -0.06300103, 
    -0.0610615, -0.06192869, -0.05875572, -0.05964112, -0.05711747, 
    -0.05774217, -0.05714664, -0.0573266, -0.0571443, -0.05806318, 
    -0.05766774, -0.05848278, -0.06176534, -0.06078242, -0.06375982, 
    -0.0656177, -0.06688114, -0.06779191, -0.06766242, -0.06741621, 
    -0.06616486, -0.06500912, -0.06414154, -0.06356748, -0.06300677, 
    -0.06133831, -0.06047302, -0.05857818, -0.05891594, -0.05834495, 
    -0.05780468, -0.05690836, -0.05705497, -0.05666338, -0.05836004, 
    -0.05722697, -0.05910914, -0.05858844, -0.06285464, -0.06455889, 
    -0.06529635, -0.06594899, -0.06756301, -0.06644432, -0.06688313, 
    -0.06584388, -0.06519163, -0.06551345, -0.06355186, -0.06430756, 
    -0.06042211, -0.06206687, -0.05786745, -0.05884647, -0.05763517, 
    -0.05825023, -0.05720018, -0.05814438, -0.05651834, -0.05617012, 
    -0.05640785, -0.05550013, -0.05819715, -0.0571466, -0.06552247, 
    -0.06546987, -0.06522541, -0.06630667, -0.06637341, -0.06738075, 
    -0.06648374, -0.06610525, -0.06515406, -0.06459762, -0.06407299, 
    -0.06293404, -0.06168524, -0.05997949, -0.05878251, -0.05799318, 
    -0.05847599, -0.05804953, -0.05852645, -0.05875131, -0.05630032, 
    -0.05766403, -0.0556298, -0.05574054, -0.05665408, -0.05572805, 
    -0.06543297, -0.06573606, -0.06679882, -0.0659657, -0.06749135, 
    -0.06663311, -0.06614441, -0.06429157, -0.06389143, -0.0635224, 
    -0.06279976, -0.06188401, -0.06030882, -0.05897014, -0.05777342, 
    -0.0578603, -0.0578297, -0.0575653, -0.05822232, -0.05745814, 
    -0.05733079, -0.05766425, -0.05575538, -0.05629438, -0.05574289, 
    -0.0560932, -0.06563739, -0.06512896, -0.06540322, -0.0648884, 
    -0.06525064, -0.06365471, -0.06318367, -0.06102441, -0.06190188, 
    -0.06051123, -0.06175925, -0.06153627, -0.06046617, -0.06169121, 
    -0.05904309, -0.06082587, -0.05755505, -0.05929147, -0.05744789, 
    -0.05777854, -0.05723213, -0.05674697, -0.05614239, -0.05504308, 
    -0.05529578, -0.05438858, -0.06437816, -0.06373169, -0.06378846, 
    -0.06311819, -0.06262688, -0.06157485, -0.05992322, -0.06053921, 
    -0.05941314, -0.05918951, -0.06090222, -0.05984493, -0.06330266, 
    -0.06273104, -0.06307084, -0.06432687, -0.06039659, -0.06238344, 
    -0.05876291, -0.05980338, -0.05681589, -0.05828292, -0.05543535, 
    -0.05425949, -0.05317539, -0.05193465, -0.06338166, -0.06381787, 
    -0.06303896, -0.06197637, -0.06100632, -0.05973938, -0.05961126, 
    -0.05937724, -0.05877532, -0.05827378, -0.05930334, -0.05814872, 
    -0.06259898, -0.06022711, -0.06398346, -0.06282885, -0.06203856, 
    -0.06238414, -0.06061003, -0.06019906, -0.05855672, -0.05940025, 
    -0.05454735, -0.05664488, -0.05100911, -0.05252669, -0.06397094, 
    -0.0633832, -0.06137822, -0.06232439, -0.05965578, -0.05901611, 
    -0.05850111, -0.05784898, -0.05777907, -0.05739649, -0.0580247, 
    -0.05742122, -0.05973672, -0.05869097, -0.06160435, -0.06088251, 
    -0.06121359, -0.06157869, -0.06045862, -0.05928697, -0.05926234, 
    -0.05889146, -0.05785821, -0.0596452, -0.05428193, -0.05753568, 
    -0.06274829, -0.06164166, -0.06148535, -0.06191067, -0.05907993, 
    -0.06009073, -0.05740581, -0.05811975, -0.05695448, -0.05753064, 
    -0.05761588, -0.05836531, -0.05883664, -0.06004399, -0.06104414, 
    -0.06184882, -0.06166081, -0.06078006, -0.05921606, -0.05777267, 
    -0.05808588, -0.05704224, -0.05984547, -0.058654, -0.0591117, 
    -0.05792552, -0.06055563, -0.05830834, -0.06114339, -0.06088958, 
    -0.06011097, -0.05857392, -0.0582393, -0.05788378, -0.05810294, 
    -0.0591769, -0.05935475, -0.06012981, -0.06034546, -0.06094477, 
    -0.06144524, -0.06098778, -0.0605109, -0.0591765, -0.05799844, 
    -0.05674008, -0.05643625, -0.0550067, -0.05616751, -0.05426429, 
    -0.055878, -0.05311346, -0.05818085, -0.05592645, -0.06007582, 
    -0.05961483, -0.0587896, -0.05693892, -0.05793104, -0.05677248, 
    -0.05936174, -0.06074981, -0.06111425, -0.06179958, -0.06109867, 
    -0.0611554, -0.06049134, -0.06070397, -0.0591327, -0.05997174, 
    -0.05761798, -0.05678158, -0.05448292, -0.05311866, -0.05176425, 
    -0.05117695, -0.0509995, -0.05092549,
  -0.06388928, -0.06219715, -0.0625229, -0.06118153, -0.0619224, -0.06104876, 
    -0.06354293, -0.06213076, -0.06302895, -0.06373534, -0.05865277, 
    -0.06112232, -0.05618465, -0.05768888, -0.05397796, -0.05641627, 
    -0.05349807, -0.05404709, -0.05241031, -0.05287457, -0.05082989, 
    -0.05219728, -0.0497986, -0.05115354, -0.05093935, -0.05224293, 
    -0.06061802, -0.05895514, -0.06071783, -0.06047777, -0.06058542, 
    -0.06190696, -0.06258274, -0.06402045, -0.06375724, -0.06270243, 
    -0.06037011, -0.06115292, -0.05919786, -0.05924137, -0.05713037, 
    -0.05807355, -0.05462801, -0.05558793, -0.05285512, -0.05353065, 
    -0.05288665, -0.0530812, -0.05288412, -0.05387804, -0.05345013, 
    -0.05433235, -0.05789581, -0.05682706, -0.06006872, -0.06209783, 
    -0.06348035, -0.06447828, -0.06433633, -0.0640665, -0.0626963, 
    -0.06143264, -0.06048524, -0.05985893, -0.05924763, -0.05743131, 
    -0.05649096, -0.05443567, -0.05480162, -0.05418308, -0.05359829, 
    -0.05262914, -0.05278758, -0.05236448, -0.05419942, -0.05297349, 
    -0.05501103, -0.05444678, -0.05908186, -0.06094085, -0.06174652, 
    -0.06246014, -0.06422738, -0.06300212, -0.06348255, -0.06234517, 
    -0.06163208, -0.06198385, -0.05984189, -0.06066645, -0.05643566, 
    -0.05822394, -0.0536662, -0.05472634, -0.0534149, -0.05408052, 
    -0.05294453, -0.05396593, -0.05220784, -0.0518319, -0.05208853, 
    -0.05110915, -0.05402305, -0.05288661, -0.06199371, -0.0619362, 
    -0.06166898, -0.06285147, -0.06292451, -0.06402764, -0.06304528, 
    -0.06263109, -0.06159102, -0.06098315, -0.06041043, -0.05916838, 
    -0.05780866, -0.0559551, -0.05465704, -0.05380227, -0.05432499, 
    -0.05386326, -0.05437963, -0.05462323, -0.05197244, -0.05344613, 
    -0.05124898, -0.0513684, -0.05235443, -0.05135494, -0.06189585, 
    -0.06222724, -0.06339023, -0.06247842, -0.06414884, -0.06320879, 
    -0.06267393, -0.06064899, -0.0602123, -0.05980976, -0.05902207, 
    -0.05802493, -0.05631263, -0.05486036, -0.05356447, -0.05365847, 
    -0.05362536, -0.05333933, -0.0540503, -0.05322343, -0.05308574, 
    -0.05344636, -0.05138442, -0.05196603, -0.05137095, -0.05174889, 
    -0.06211936, -0.06156359, -0.06186333, -0.06130075, -0.06169656, 
    -0.05995407, -0.05944045, -0.05709006, -0.05804438, -0.05653245, 
    -0.05788918, -0.05764661, -0.05648351, -0.05781515, -0.05493944, 
    -0.05687429, -0.05332824, -0.05520871, -0.05321235, -0.05357001, 
    -0.05297907, -0.05245478, -0.05180197, -0.05061655, -0.05088887, 
    -0.04991176, -0.06074352, -0.06003804, -0.06009996, -0.05936906, 
    -0.05883372, -0.05768857, -0.05589403, -0.05656285, -0.05534064, 
    -0.05509815, -0.05695726, -0.05580906, -0.05957016, -0.05894719, 
    -0.05931746, -0.06068753, -0.05640794, -0.0585686, -0.0546358, 
    -0.05576398, -0.05252923, -0.05411591, -0.05103932, -0.04977284, 
    -0.04860735, -0.04727606, -0.05965629, -0.06013205, -0.05928272, 
    -0.05812544, -0.05707039, -0.05569454, -0.05555554, -0.05530172, 
    -0.05464925, -0.05410602, -0.05522158, -0.05397063, -0.05880334, 
    -0.05622391, -0.06031271, -0.05905375, -0.05819313, -0.05856935, 
    -0.05663978, -0.05619346, -0.05441243, -0.05532667, -0.05008267, 
    -0.0523445, -0.04628484, -0.04791096, -0.06029906, -0.05965798, 
    -0.05747471, -0.05850429, -0.05560384, -0.05491019, -0.05435219, 
    -0.05364623, -0.05357058, -0.05315677, -0.05383638, -0.05318351, 
    -0.05569165, -0.05455786, -0.05772066, -0.05693582, -0.0572957, 
    -0.05769275, -0.05647531, -0.05520383, -0.05517712, -0.0547751, 
    -0.05365622, -0.05559236, -0.04979699, -0.0533073, -0.05896598, 
    -0.05776125, -0.05759122, -0.05805394, -0.05497937, -0.05607585, 
    -0.05316685, -0.05393926, -0.05267898, -0.05330184, -0.05339404, 
    -0.05420513, -0.05471568, -0.05602511, -0.0571115, -0.05798664, 
    -0.05778208, -0.0568245, -0.05512695, -0.05356366, -0.0539026, 
    -0.05277381, -0.05580966, -0.05451781, -0.0550138, -0.05372904, 
    -0.05658068, -0.05414344, -0.05721938, -0.05694352, -0.05609782, 
    -0.05443106, -0.05406868, -0.05368388, -0.05392106, -0.05508449, 
    -0.05527733, -0.05611828, -0.05635242, -0.05700349, -0.0575476, 
    -0.05705024, -0.0565321, -0.05508406, -0.05380796, -0.05244733, 
    -0.0521192, -0.05057735, -0.05182908, -0.04977801, -0.05151669, 
    -0.04854084, -0.05400541, -0.05156896, -0.05605966, -0.05555942, 
    -0.05466472, -0.05266216, -0.05373502, -0.05248233, -0.05528491, 
    -0.05679163, -0.05718771, -0.05793306, -0.05717077, -0.05723244, 
    -0.05651085, -0.05674183, -0.05503657, -0.05594669, -0.05339631, 
    -0.05249216, -0.0500133, -0.04854642, -0.04709344, -0.04646447, 
    -0.04627455, -0.04619535,
  -0.04035026, -0.03907193, -0.03931788, -0.03830562, -0.03886456, 
    -0.03820549, -0.04008846, -0.03902182, -0.03970009, -0.04023389, 
    -0.03640087, -0.03826097, -0.03454665, -0.03567613, -0.03289328, 
    -0.03472044, -0.03253432, -0.03294501, -0.03172149, -0.03206827, 
    -0.03054266, -0.03156244, -0.02977487, -0.03078386, -0.03062422, 
    -0.03159652, -0.03788075, -0.03662837, -0.03795599, -0.03777504, 
    -0.03785618, -0.0388529, -0.03936306, -0.04044943, -0.04025044, 
    -0.03945345, -0.03769391, -0.03828404, -0.03681104, -0.0368438, 
    -0.03525654, -0.03596527, -0.03337988, -0.03409912, -0.03205374, 
    -0.03255868, -0.03207729, -0.03222268, -0.0320754, -0.03281852, 
    -0.03249847, -0.03315851, -0.03583166, -0.03502879, -0.03746682, 
    -0.03899696, -0.04004116, -0.04079566, -0.0406883, -0.04048425, 
    -0.03944882, -0.03849502, -0.03778067, -0.03730879, -0.0368485, 
    -0.0354826, -0.03477649, -0.03323586, -0.03350989, -0.03304678, 
    -0.03260927, -0.03188492, -0.03200327, -0.03168726, -0.03305901, 
    -0.03214218, -0.03366677, -0.03324417, -0.03672373, -0.03812413, 
    -0.03873183, -0.03927049, -0.0406059, -0.03967981, -0.04004281, 
    -0.03918368, -0.03864548, -0.03891093, -0.03729596, -0.03791726, 
    -0.03473499, -0.03607835, -0.03266006, -0.03345351, -0.03247213, 
    -0.03297002, -0.03212054, -0.03288428, -0.03157032, -0.03128976, 
    -0.03148126, -0.03075077, -0.03292702, -0.03207726, -0.03891837, 
    -0.03887497, -0.03867333, -0.03956602, -0.03962119, -0.04045487, 
    -0.03971241, -0.03939957, -0.0386145, -0.03815602, -0.03772429, 
    -0.03678885, -0.03576615, -0.03437445, -0.03340161, -0.03276184, 
    -0.033153, -0.03280746, -0.0331939, -0.03337629, -0.03139462, 
    -0.03249548, -0.030855, -0.03094404, -0.03167976, -0.030934, -0.03884452, 
    -0.03909465, -0.03997305, -0.03928429, -0.04054652, -0.03983595, 
    -0.03943193, -0.03790409, -0.037575, -0.03727176, -0.03667873, 
    -0.03592872, -0.03464267, -0.03355389, -0.03258397, -0.03265428, 
    -0.03262951, -0.03241563, -0.03294741, -0.03232898, -0.03222606, 
    -0.03249566, -0.03095598, -0.03138984, -0.03094594, -0.03122782, 
    -0.03901321, -0.03859381, -0.03881998, -0.03839554, -0.03869413, 
    -0.03738046, -0.03699366, -0.03522626, -0.03594334, -0.03480763, 
    -0.03582668, -0.03564437, -0.0347709, -0.03577103, -0.03361313, 
    -0.03506424, -0.03240734, -0.03381488, -0.0323207, -0.03258811, 
    -0.03214635, -0.03175469, -0.03126742, -0.03038373, -0.0305866, 
    -0.02985905, -0.03797536, -0.03744371, -0.03749036, -0.03693992, 
    -0.03653701, -0.0356759, -0.03432865, -0.03483044, -0.03391375, 
    -0.03373204, -0.03512654, -0.03426493, -0.03709132, -0.03662238, 
    -0.03690107, -0.03793315, -0.03471419, -0.03633755, -0.03338571, 
    -0.03423112, -0.03181029, -0.03299651, -0.03069872, -0.0297557, 
    -0.02888947, -0.02790199, -0.03715618, -0.03751453, -0.03687492, 
    -0.03600429, -0.0352115, -0.03417906, -0.03407484, -0.03388458, 
    -0.03339577, -0.03298911, -0.03382453, -0.03288779, -0.03651415, 
    -0.0345761, -0.03765066, -0.03670258, -0.03605518, -0.03633812, 
    -0.03488819, -0.03455326, -0.03321846, -0.03390329, -0.02998624, 
    -0.03167235, -0.02716819, -0.02837265, -0.03764037, -0.03715745, 
    -0.03551521, -0.03628918, -0.03411105, -0.03359121, -0.03317336, 
    -0.03264511, -0.03258854, -0.03227916, -0.03278736, -0.03229914, 
    -0.03417689, -0.03332734, -0.03570002, -0.03511045, -0.03538072, 
    -0.03567904, -0.03476474, -0.03381122, -0.03379121, -0.03349003, 
    -0.03265259, -0.03410244, -0.02977367, -0.03239168, -0.03663653, 
    -0.03573052, -0.03560275, -0.03595053, -0.03364304, -0.03446503, 
    -0.03228669, -0.03286433, -0.03192214, -0.0323876, -0.03245653, 
    -0.03306328, -0.03344553, -0.03442697, -0.03524237, -0.03589994, 
    -0.03574618, -0.03502686, -0.03375361, -0.03258337, -0.0328369, 
    -0.03199298, -0.03426538, -0.03329735, -0.03366884, -0.03270706, 
    -0.03484383, -0.03301711, -0.0353234, -0.03511622, -0.0344815, 
    -0.03323241, -0.03296117, -0.03267328, -0.03285071, -0.0337218, 
    -0.0338663, -0.03449685, -0.03467252, -0.03516125, -0.03556997, 
    -0.03519636, -0.03480737, -0.03372148, -0.0327661, -0.03174913, 
    -0.03150415, -0.03035454, -0.03128765, -0.02975954, -0.03105462, 
    -0.02884008, -0.03291382, -0.03109361, -0.03445289, -0.03407775, 
    -0.03340736, -0.03190958, -0.03271153, -0.03177527, -0.03387198, 
    -0.03500219, -0.03529961, -0.03585966, -0.03528689, -0.0353332, 
    -0.03479142, -0.0349648, -0.0336859, -0.03436815, -0.03245823, 
    -0.03178261, -0.02993461, -0.02884423, -0.0277667, -0.02730108, 
    -0.02716058, -0.02710201,
  -0.01970495, -0.01870051, -0.01889313, -0.01810234, -0.01853834, 
    -0.01802441, -0.01949858, -0.0186613, -0.01919307, -0.01961318, 
    -0.01662921, -0.01806758, -0.01521542, -0.01607413, -0.01397334, 
    -0.01534703, -0.01370616, -0.01401192, -0.01310461, -0.01336065, 
    -0.01224113, -0.01298748, -0.01168475, -0.01241692, -0.01230052, 
    -0.01301256, -0.01777202, -0.01680409, -0.01783044, -0.01768999, 
    -0.01775294, -0.01852923, -0.01892855, -0.0197832, -0.01962623, 
    -0.01899944, -0.01762707, -0.01808554, -0.01694472, -0.01696996, 
    -0.0157542, -0.01629521, -0.01433697, -0.01487742, -0.01334991, 
    -0.01372427, -0.01336733, -0.01347495, -0.01336593, -0.01391762, 
    -0.01367953, -0.01417134, -0.01619298, -0.015581, -0.01745114, 
    -0.01864185, -0.01946134, -0.02005678, -0.01997189, -0.01981069, 
    -0.0189958, -0.0182499, -0.01769435, -0.01732889, -0.01697359, 
    -0.01592643, -0.01538952, -0.01422918, -0.01443441, -0.01408788, 
    -0.01376187, -0.01322517, -0.01331259, -0.01307939, -0.01409701, 
    -0.01341534, -0.01455213, -0.0142354, -0.01687748, -0.01796112, 
    -0.01843466, -0.01885599, -0.01990677, -0.01917714, -0.01946264, 
    -0.01878799, -0.01836725, -0.01857458, -0.01731896, -0.01780037, 
    -0.01535806, -0.01638181, -0.01379965, -0.01439214, -0.01365996, 
    -0.01403059, -0.01339933, -0.01396663, -0.01299328, -0.01278711, 
    -0.01292777, -0.01239277, -0.01399851, -0.01336731, -0.0185804, 
    -0.01854647, -0.01838898, -0.01908778, -0.01913109, -0.0197875, 
    -0.01920276, -0.01895718, -0.01834308, -0.01798592, -0.01765062, 
    -0.01692763, -0.01614291, -0.01508522, -0.01435326, -0.0138754, 
    -0.01416723, -0.01390938, -0.01419781, -0.01433429, -0.0128641, 
    -0.0136773, -0.01246885, -0.01253391, -0.01307387, -0.01252657, 
    -0.01852268, -0.01871829, -0.01940772, -0.0188668, -0.01985986, 
    -0.01929986, -0.01898255, -0.01779014, -0.01753491, -0.01730026, 
    -0.01684284, -0.01626723, -0.01528811, -0.01446741, -0.01374306, 
    -0.01379535, -0.01377692, -0.01361802, -0.01401371, -0.01355374, 
    -0.01347746, -0.01367744, -0.01254264, -0.01286059, -0.0125353, 
    -0.01274168, -0.01865457, -0.01832694, -0.0185035, -0.01817236, 
    -0.01840522, -0.01738431, -0.01708551, -0.01573116, -0.01627842, 
    -0.01541313, -0.01618917, -0.01604987, -0.01538528, -0.01614664, 
    -0.01451186, -0.01560794, -0.01361187, -0.01466342, -0.0135476, 
    -0.01374614, -0.01341843, -0.01312909, -0.01277073, -0.01212556, 
    -0.01227312, -0.01174552, -0.01784549, -0.01743326, -0.01746936, 
    -0.01704406, -0.01673382, -0.01607395, -0.01505062, -0.01543043, 
    -0.0147378, -0.01460116, -0.0156553, -0.0150025, -0.01716087, 
    -0.01679948, -0.0170141, -0.01781271, -0.01534229, -0.01658059, 
    -0.01434134, -0.01497698, -0.0131701, -0.01405035, -0.01235481, 
    -0.01167093, -0.01104941, -0.0103492, -0.01721095, -0.01748808, 
    -0.01699394, -0.01632508, -0.01571992, -0.0149377, -0.01485912, 
    -0.01471585, -0.01434888, -0.01404483, -0.01467068, -0.01396925, 
    -0.01671625, -0.01523771, -0.01759354, -0.0168612, -0.01636406, 
    -0.01658103, -0.01547424, -0.01522042, -0.01421617, -0.01472993, 
    -0.01183743, -0.0130684, -0.009834954, -0.01068181, -0.01758556, 
    -0.01721193, -0.0159513, -0.01654346, -0.01488641, -0.01449542, 
    -0.01418244, -0.01378853, -0.01374646, -0.0135168, -0.01389441, 
    -0.01353162, -0.01493606, -0.01429764, -0.01609237, -0.01564307, 
    -0.01584878, -0.01607635, -0.01538061, -0.01466068, -0.01464563, 
    -0.01441952, -0.01379409, -0.01487993, -0.01168389, -0.01360025, 
    -0.01681037, -0.01611568, -0.0160181, -0.01628392, -0.01453432, 
    -0.01515368, -0.01352238, -0.01395176, -0.01325265, -0.01359722, 
    -0.01364838, -0.0141002, -0.01438616, -0.0151249, -0.01574342, 
    -0.01624521, -0.01612764, -0.01557954, -0.01461737, -0.01374261, 
    -0.01393132, -0.01330499, -0.01500284, -0.01427519, -0.01455369, 
    -0.01383462, -0.01544059, -0.01406573, -0.01580511, -0.01564746, 
    -0.01516614, -0.0142266, -0.01402398, -0.01380948, -0.01394161, 
    -0.01459347, -0.0147021, -0.01517775, -0.01531073, -0.0156817, 
    -0.01599308, -0.01570841, -0.01541293, -0.01459322, -0.01387857, 
    -0.01312499, -0.0129446, -0.01210436, -0.01278557, -0.0116737, 
    -0.0126148, -0.01101418, -0.01398866, -0.01264334, -0.0151445, 
    -0.01486131, -0.01435756, -0.01324338, -0.01383795, -0.01314426, 
    -0.01470637, -0.0155608, -0.01578699, -0.0162144, -0.01577731, 
    -0.01581258, -0.01540083, -0.0155324, -0.0145665, -0.01508045, 
    -0.01364965, -0.01314967, -0.01180011, -0.01101713, -0.01025399, 
    -0.009927681, -0.009829648, -0.009788837,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  362.8776, 364.6899, 364.337, 365.8023, 364.9889, 365.9492, 363.2444, 
    364.7621, 363.7927, 363.0403, 368.6572, 365.8677, 371.5505, 369.7754, 
    374.2446, 371.2741, 374.8453, 374.1583, 376.2275, 375.634, 378.3688, 
    376.5017, 379.7498, 377.9411, 378.2238, 376.4429, 366.4277, 368.3092, 
    366.3165, 366.5844, 366.4641, 365.0058, 364.2726, 362.7391, 363.0171, 
    364.1434, 366.7048, 365.8338, 368.0309, 367.9811, 370.4288, 369.3284, 
    373.4393, 372.268, 375.6588, 374.8042, 375.6186, 375.3715, 375.6219, 
    374.3691, 374.9055, 373.8042, 369.5349, 370.7865, 367.0432, 364.798, 
    363.3109, 362.2583, 362.407, 362.6906, 364.1501, 365.5254, 366.5759, 
    367.2797, 367.974, 370.0762, 371.1852, 373.6765, 373.2259, 373.9893, 
    374.7193, 375.9471, 375.7448, 376.2865, 373.969, 375.5083, 372.9694, 
    373.6627, 368.164, 366.0686, 365.1813, 364.4049, 362.5213, 363.8215, 
    363.3086, 364.5293, 365.3064, 364.9219, 367.299, 366.3737, 371.2509, 
    369.1534, 374.6341, 373.3183, 374.9499, 374.1167, 375.5451, 374.2594, 
    376.4881, 377.0536, 376.6422, 377.9995, 374.1882, 375.6187, 364.9112, 
    364.9738, 365.266, 363.9831, 363.9047, 362.7315, 363.7752, 364.2203, 
    365.3514, 366.0217, 366.6596, 368.0646, 369.6361, 371.8256, 373.4035, 
    374.4637, 373.8133, 374.3875, 373.7457, 373.4451, 376.8712, 374.9106, 
    377.8154, 377.6586, 376.2994, 377.6763, 365.0179, 364.6571, 363.4068, 
    364.3851, 362.6039, 363.6003, 364.1742, 366.3932, 366.8817, 367.3353, 
    368.2321, 369.3851, 371.3975, 373.1539, 374.7617, 374.6437, 374.6853, 
    375.0451, 374.1543, 375.1915, 375.3658, 374.9102, 377.6376, 376.8795, 
    377.6553, 377.1615, 364.7744, 365.3815, 365.0534, 365.6707, 365.2358, 
    367.1725, 367.7544, 370.4764, 369.3625, 371.1357, 369.5426, 369.8246, 
    371.1942, 369.6285, 373.0571, 370.7308, 375.0591, 372.7285, 375.2055, 
    374.7547, 375.5011, 376.1705, 377.0925, 378.652, 378.2905, 379.5967, 
    366.2878, 367.0778, 367.008, 367.8355, 368.4484, 369.7757, 371.899, 
    371.0995, 372.5677, 372.863, 370.6326, 372.0013, 367.6068, 368.3181, 
    367.8944, 366.3503, 371.2839, 368.7541, 373.4297, 372.0555, 376.075, 
    374.0728, 378.0916, 379.7848, 381.3816, 383.2541, 367.5091, 366.9719, 
    367.934, 369.2681, 370.4994, 372.1393, 372.3072, 372.6151, 373.4131, 
    374.085, 372.7127, 374.2535, 368.4836, 371.5035, 366.7691, 368.1959, 
    369.1893, 368.7531, 371.0082, 371.5398, 373.7053, 372.5847, 379.3666, 
    376.3123, 384.683, 382.3546, 366.7843, 367.5071, 370.0252, 368.8283, 
    372.2488, 373.0928, 373.7796, 374.6591, 374.754, 375.2758, 374.4211, 
    375.2419, 372.1428, 373.5257, 369.7383, 370.658, 370.2346, 369.7708, 
    371.2036, 372.7343, 372.7667, 373.2585, 374.6471, 372.2627, 379.7524, 
    375.086, 368.2964, 369.6913, 369.8891, 369.3513, 373.0081, 371.6807, 
    375.2631, 374.2926, 375.8834, 375.0924, 374.9761, 373.9619, 373.3314, 
    371.7415, 370.451, 369.4296, 369.6669, 370.7895, 372.828, 374.7628, 
    374.3385, 375.7624, 372.0004, 373.5751, 372.9661, 374.5553, 371.0784, 
    374.0389, 370.3242, 370.6488, 371.6543, 373.6823, 374.1314, 374.612, 
    374.3153, 372.8798, 372.6447, 371.6298, 371.35, 370.5781, 369.94, 
    370.5231, 371.1361, 372.8802, 374.4566, 376.1801, 376.6025, 378.7044, 
    377.0575, 379.7781, 377.465, 381.4742, 374.2104, 377.3964, 371.7, 
    372.3025, 373.3942, 375.9051, 374.5479, 376.1353, 372.6355, 370.8284, 
    370.3614, 369.4917, 370.3813, 370.3089, 371.1613, 370.8872, 372.9382, 
    371.8356, 374.9733, 376.1227, 379.4598, 381.4662, 383.5149, 384.4217, 
    384.6979, 384.8134 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.215665e-08, 6.243071e-08, 6.237744e-08, 6.25985e-08, 6.247588e-08, 
    6.262062e-08, 6.221222e-08, 6.244159e-08, 6.229516e-08, 6.218133e-08, 
    6.302749e-08, 6.260836e-08, 6.346296e-08, 6.319562e-08, 6.386725e-08, 
    6.342135e-08, 6.395716e-08, 6.38544e-08, 6.416374e-08, 6.407512e-08, 
    6.447078e-08, 6.420464e-08, 6.467591e-08, 6.440724e-08, 6.444926e-08, 
    6.419586e-08, 6.269272e-08, 6.29753e-08, 6.267597e-08, 6.271627e-08, 
    6.269819e-08, 6.247841e-08, 6.236764e-08, 6.213571e-08, 6.217782e-08, 
    6.234817e-08, 6.273439e-08, 6.260329e-08, 6.293373e-08, 6.292627e-08, 
    6.329415e-08, 6.312828e-08, 6.374665e-08, 6.357089e-08, 6.407881e-08, 
    6.395107e-08, 6.407281e-08, 6.40359e-08, 6.407329e-08, 6.388595e-08, 
    6.396621e-08, 6.380137e-08, 6.315934e-08, 6.334801e-08, 6.27853e-08, 
    6.244696e-08, 6.222228e-08, 6.206283e-08, 6.208537e-08, 6.212834e-08, 
    6.234917e-08, 6.255681e-08, 6.271505e-08, 6.28209e-08, 6.29252e-08, 
    6.324087e-08, 6.3408e-08, 6.378219e-08, 6.371467e-08, 6.382906e-08, 
    6.393837e-08, 6.412186e-08, 6.409167e-08, 6.41725e-08, 6.382605e-08, 
    6.40563e-08, 6.36762e-08, 6.378016e-08, 6.29535e-08, 6.263866e-08, 
    6.25048e-08, 6.238768e-08, 6.21027e-08, 6.22995e-08, 6.222191e-08, 
    6.24065e-08, 6.252378e-08, 6.246577e-08, 6.282379e-08, 6.26846e-08, 
    6.34179e-08, 6.310203e-08, 6.392562e-08, 6.372853e-08, 6.397286e-08, 
    6.384818e-08, 6.40618e-08, 6.386955e-08, 6.42026e-08, 6.427513e-08, 
    6.422556e-08, 6.441596e-08, 6.385889e-08, 6.407281e-08, 6.246415e-08, 
    6.247361e-08, 6.251769e-08, 6.232393e-08, 6.231208e-08, 6.213455e-08, 
    6.229253e-08, 6.23598e-08, 6.253058e-08, 6.263159e-08, 6.272763e-08, 
    6.293877e-08, 6.317458e-08, 6.350436e-08, 6.37413e-08, 6.390013e-08, 
    6.380274e-08, 6.388873e-08, 6.37926e-08, 6.374756e-08, 6.424796e-08, 
    6.396696e-08, 6.438858e-08, 6.436525e-08, 6.417443e-08, 6.436788e-08, 
    6.248025e-08, 6.242581e-08, 6.223679e-08, 6.238472e-08, 6.211522e-08, 
    6.226607e-08, 6.23528e-08, 6.26875e-08, 6.276105e-08, 6.282924e-08, 
    6.296392e-08, 6.313677e-08, 6.343999e-08, 6.370384e-08, 6.394473e-08, 
    6.392708e-08, 6.393329e-08, 6.398709e-08, 6.385381e-08, 6.400898e-08, 
    6.403502e-08, 6.396693e-08, 6.436213e-08, 6.424923e-08, 6.436476e-08, 
    6.429125e-08, 6.244351e-08, 6.253511e-08, 6.248561e-08, 6.257869e-08, 
    6.251312e-08, 6.28047e-08, 6.289213e-08, 6.330126e-08, 6.313336e-08, 
    6.340058e-08, 6.316051e-08, 6.320305e-08, 6.340928e-08, 6.317349e-08, 
    6.368928e-08, 6.333956e-08, 6.398919e-08, 6.363992e-08, 6.401108e-08, 
    6.394369e-08, 6.405527e-08, 6.41552e-08, 6.428095e-08, 6.451294e-08, 
    6.445922e-08, 6.465324e-08, 6.267168e-08, 6.279049e-08, 6.278004e-08, 
    6.290439e-08, 6.299635e-08, 6.319569e-08, 6.351541e-08, 6.339518e-08, 
    6.361591e-08, 6.366022e-08, 6.332489e-08, 6.353077e-08, 6.287001e-08, 
    6.297676e-08, 6.291321e-08, 6.268105e-08, 6.342287e-08, 6.304215e-08, 
    6.374522e-08, 6.353896e-08, 6.414095e-08, 6.384155e-08, 6.442965e-08, 
    6.468104e-08, 6.491769e-08, 6.519421e-08, 6.285535e-08, 6.277462e-08, 
    6.291918e-08, 6.311918e-08, 6.330479e-08, 6.355153e-08, 6.357678e-08, 
    6.362301e-08, 6.374275e-08, 6.384343e-08, 6.363761e-08, 6.386867e-08, 
    6.300149e-08, 6.345593e-08, 6.274409e-08, 6.295841e-08, 6.31074e-08, 
    6.304205e-08, 6.338144e-08, 6.346144e-08, 6.37865e-08, 6.361847e-08, 
    6.461898e-08, 6.41763e-08, 6.540478e-08, 6.506145e-08, 6.27464e-08, 
    6.285507e-08, 6.323329e-08, 6.305333e-08, 6.356801e-08, 6.36947e-08, 
    6.37977e-08, 6.392935e-08, 6.394357e-08, 6.402158e-08, 6.389375e-08, 
    6.401653e-08, 6.355206e-08, 6.375961e-08, 6.319006e-08, 6.332868e-08, 
    6.326491e-08, 6.319497e-08, 6.341085e-08, 6.364085e-08, 6.364578e-08, 
    6.371953e-08, 6.392733e-08, 6.35701e-08, 6.467609e-08, 6.399301e-08, 
    6.297358e-08, 6.318288e-08, 6.321279e-08, 6.313171e-08, 6.368199e-08, 
    6.34826e-08, 6.401968e-08, 6.387452e-08, 6.411236e-08, 6.399417e-08, 
    6.397678e-08, 6.3825e-08, 6.373049e-08, 6.349174e-08, 6.329749e-08, 
    6.314347e-08, 6.317929e-08, 6.334847e-08, 6.365492e-08, 6.394485e-08, 
    6.388134e-08, 6.409429e-08, 6.353069e-08, 6.3767e-08, 6.367566e-08, 
    6.391384e-08, 6.339199e-08, 6.383632e-08, 6.327841e-08, 6.332733e-08, 
    6.347864e-08, 6.378302e-08, 6.385039e-08, 6.392229e-08, 6.387792e-08, 
    6.366271e-08, 6.362745e-08, 6.347497e-08, 6.343286e-08, 6.331668e-08, 
    6.322048e-08, 6.330837e-08, 6.340066e-08, 6.36628e-08, 6.389904e-08, 
    6.415662e-08, 6.421966e-08, 6.452062e-08, 6.427562e-08, 6.46799e-08, 
    6.433616e-08, 6.493121e-08, 6.38621e-08, 6.432608e-08, 6.348553e-08, 
    6.357608e-08, 6.373985e-08, 6.411551e-08, 6.391272e-08, 6.414989e-08, 
    6.362608e-08, 6.335431e-08, 6.328401e-08, 6.315283e-08, 6.328701e-08, 
    6.32761e-08, 6.340449e-08, 6.336324e-08, 6.367151e-08, 6.350592e-08, 
    6.397634e-08, 6.414802e-08, 6.46329e-08, 6.493014e-08, 6.523275e-08, 
    6.536635e-08, 6.540701e-08, 6.542402e-08 ;

 SOM_C_LEACHED =
  4.637716e-20, 4.137485e-20, 6.259535e-20, 3.229206e-21, -1.287217e-20, 
    -4.70693e-20, -4.575063e-20, -2.816551e-20, 1.398816e-20, -1.723467e-20, 
    1.040991e-20, 5.730806e-20, -1.980563e-20, -6.343835e-20, 7.899905e-21, 
    1.4597e-21, -6.344179e-20, -3.782745e-20, -3.094175e-20, -7.924673e-21, 
    -3.650978e-20, 8.57836e-21, -1.340286e-20, -3.788312e-20, -2.252079e-20, 
    -1.091026e-20, -2.243247e-20, -6.220446e-21, -3.000862e-20, 2.378762e-20, 
    3.569608e-20, -9.239765e-21, 3.785788e-20, 5.212655e-20, 3.99342e-20, 
    -1.207149e-20, -3.200146e-20, 8.916069e-20, -2.210676e-20, 2.378463e-20, 
    -5.885021e-20, -5.423331e-20, -1.794397e-20, 4.685951e-20, -3.813626e-20, 
    -5.1504e-20, 1.790727e-20, -2.153045e-20, -9.219673e-21, 1.041947e-20, 
    6.08221e-20, 1.253181e-20, 5.036005e-20, 3.658301e-21, -4.853224e-20, 
    -2.710538e-21, -7.488792e-21, -2.781595e-20, -3.206252e-20, 
    -4.054071e-20, 3.01545e-20, 1.629331e-20, 2.021857e-21, -4.9593e-20, 
    -1.414181e-20, -3.380079e-20, 3.733464e-20, -2.003137e-20, -3.552552e-20, 
    -1.845279e-20, 2.135445e-21, -2.71762e-20, 4.053589e-20, -5.237327e-20, 
    1.539941e-20, -3.643517e-20, 3.559425e-20, 1.212204e-21, -4.912852e-20, 
    2.567346e-20, -2.983981e-21, 2.62718e-20, 5.851384e-20, -7.723097e-21, 
    9.718362e-21, -1.239772e-20, -8.760194e-21, -2.728304e-21, -7.526749e-21, 
    5.172011e-21, -7.787248e-20, -2.548168e-20, -2.471879e-20, -6.7779e-20, 
    -3.272846e-20, -4.166866e-21, 2.391761e-20, 2.198153e-20, 2.288198e-20, 
    2.182572e-20, -5.20742e-20, -6.065187e-20, 5.913406e-20, 4.155478e-20, 
    1.56447e-20, 2.181947e-21, -3.609389e-20, 2.526981e-20, 1.374941e-21, 
    -5.640375e-21, -7.144833e-20, 6.400481e-20, 1.047396e-20, -1.563948e-20, 
    -5.777509e-20, 5.643668e-20, -9.063895e-20, -3.332686e-20, -6.86473e-20, 
    1.107293e-20, 3.982177e-20, -2.090471e-20, 1.585812e-20, 4.225139e-21, 
    5.081836e-20, 4.350069e-20, 2.98101e-20, -2.049261e-21, -7.501045e-21, 
    -2.817188e-20, 1.100023e-20, 1.342651e-20, 2.937745e-20, 9.500316e-21, 
    -5.723583e-20, -2.726154e-20, 5.168169e-20, 1.668064e-20, -6.85465e-20, 
    -5.319771e-20, -5.430901e-20, 9.229484e-21, -3.272549e-20, 1.233774e-20, 
    1.838073e-20, -7.417804e-21, 4.839371e-20, 6.924538e-20, 2.157056e-20, 
    3.438323e-20, -3.231847e-21, 5.098525e-20, -4.89727e-20, -4.700003e-20, 
    9.702879e-21, -4.838593e-20, -3.668966e-21, 2.811181e-20, 3.445815e-20, 
    -1.2415e-20, 1.961794e-20, 2.779139e-20, -1.950131e-21, 1.224316e-20, 
    -4.962014e-20, -4.872029e-20, -2.190811e-20, -5.149682e-20, 
    -3.239292e-20, 5.220554e-20, 1.975159e-20, 4.401601e-20, 6.204473e-21, 
    4.510334e-20, -2.603975e-20, 4.701292e-20, -4.058502e-20, 3.853116e-21, 
    -4.061195e-20, -5.829568e-20, 1.2652e-20, -1.964719e-20, 3.40394e-20, 
    -3.587039e-20, -7.883704e-21, -1.09835e-20, -6.946229e-20, -3.081778e-20, 
    9.896509e-21, 9.263961e-21, -7.658822e-20, -4.687032e-21, 3.982734e-20, 
    2.887988e-20, -3.722346e-20, 4.902603e-20, -7.925353e-20, 4.578273e-20, 
    5.000093e-20, -5.048492e-20, 6.269955e-21, -6.188715e-21, -5.947435e-21, 
    -1.731662e-20, -3.266364e-20, -7.823433e-20, 3.65433e-20, 4.516911e-20, 
    2.565852e-20, 4.696913e-21, 1.054521e-20, -1.002386e-20, -3.098232e-20, 
    -2.580254e-20, -6.965363e-21, 3.555911e-20, -5.053511e-20, 5.667517e-20, 
    9.547614e-21, -1.05797e-20, 1.348096e-20, 3.420306e-21, 5.197794e-20, 
    1.49175e-20, -3.990803e-21, 4.572413e-20, -5.283185e-20, 1.248763e-20, 
    -1.002644e-20, 2.820163e-20, 4.162735e-22, -5.19617e-20, 3.705988e-20, 
    -4.660786e-21, -8.840195e-21, 3.591234e-20, -6.836814e-20, 1.552236e-20, 
    -4.584798e-21, -4.385222e-20, 1.946718e-20, 4.581469e-21, -4.829237e-20, 
    -3.752838e-20, 9.864438e-21, -2.200965e-20, 7.186333e-20, 3.997198e-20, 
    -1.009455e-20, -1.680472e-20, 9.145836e-21, 5.675389e-22, 1.435039e-20, 
    2.268989e-21, -3.584102e-21, 1.355803e-20, -1.285554e-20, -5.074569e-21, 
    4.963886e-21, -3.125011e-20, -2.024924e-20, 2.03307e-20, 3.094801e-20, 
    6.643309e-21, 3.614683e-20, -3.05171e-20, 2.961425e-20, 1.205157e-20, 
    -4.634866e-20, -2.965929e-20, -6.024884e-20, 2.838408e-20, -9.824155e-21, 
    -4.467088e-20, -3.026784e-20, 4.286536e-20, 1.030543e-19, 1.06414e-21, 
    7.543212e-20, -3.306886e-20, -5.903253e-21, 6.230429e-21, 3.667636e-20, 
    8.229998e-20, -2.9476e-20, -7.632953e-20, -5.034803e-21, -7.819015e-20, 
    -7.584592e-20, 7.597962e-21, 9.018868e-21, 5.378397e-20, -3.332394e-20, 
    1.435867e-21, 3.484641e-20, 6.603802e-21, -1.521094e-20, 2.50243e-20, 
    -2.827697e-20, -5.777932e-20, -2.726014e-20, -1.68563e-20, 3.071168e-20, 
    2.923012e-20, -1.029323e-20, 2.948629e-20, -5.882507e-20, -9.340193e-20, 
    -1.131196e-20, 4.048028e-20, 2.038157e-20, -4.258683e-20, 7.549497e-20, 
    2.26419e-20, -3.373283e-21, 2.020068e-20, 4.451566e-20, -5.661312e-20, 
    -1.438079e-20, 7.878849e-20, 6.667848e-21, 9.928643e-21, -2.710514e-20, 
    -2.868057e-20, -1.809289e-20, 1.823801e-20, -5.086903e-20, -3.934143e-21, 
    -4.79334e-20, 1.490389e-20, 4.215482e-20, 4.93121e-21, 6.504998e-20, 
    4.388574e-20, 2.005735e-20, -9.858027e-21, 3.475128e-20, -4.785571e-21 ;

 SR =
  6.215762e-08, 6.243169e-08, 6.237841e-08, 6.259947e-08, 6.247685e-08, 
    6.26216e-08, 6.221319e-08, 6.244257e-08, 6.229614e-08, 6.21823e-08, 
    6.302847e-08, 6.260934e-08, 6.346394e-08, 6.319659e-08, 6.386823e-08, 
    6.342233e-08, 6.395815e-08, 6.385538e-08, 6.416472e-08, 6.40761e-08, 
    6.447177e-08, 6.420563e-08, 6.46769e-08, 6.440823e-08, 6.445025e-08, 
    6.419685e-08, 6.269369e-08, 6.297628e-08, 6.267695e-08, 6.271725e-08, 
    6.269916e-08, 6.247938e-08, 6.236861e-08, 6.213668e-08, 6.217878e-08, 
    6.234914e-08, 6.273537e-08, 6.260426e-08, 6.29347e-08, 6.292724e-08, 
    6.329513e-08, 6.312926e-08, 6.374764e-08, 6.357188e-08, 6.40798e-08, 
    6.395206e-08, 6.40738e-08, 6.403688e-08, 6.407428e-08, 6.388693e-08, 
    6.39672e-08, 6.380235e-08, 6.316031e-08, 6.334899e-08, 6.278628e-08, 
    6.244793e-08, 6.222324e-08, 6.20638e-08, 6.208634e-08, 6.212931e-08, 
    6.235014e-08, 6.255778e-08, 6.271602e-08, 6.282187e-08, 6.292617e-08, 
    6.324185e-08, 6.340898e-08, 6.378317e-08, 6.371565e-08, 6.383004e-08, 
    6.393935e-08, 6.412285e-08, 6.409265e-08, 6.417349e-08, 6.382704e-08, 
    6.405729e-08, 6.367719e-08, 6.378114e-08, 6.295448e-08, 6.263964e-08, 
    6.250578e-08, 6.238865e-08, 6.210367e-08, 6.230047e-08, 6.222289e-08, 
    6.240747e-08, 6.252476e-08, 6.246675e-08, 6.282476e-08, 6.268557e-08, 
    6.341888e-08, 6.310301e-08, 6.39266e-08, 6.372951e-08, 6.397384e-08, 
    6.384917e-08, 6.406279e-08, 6.387053e-08, 6.420358e-08, 6.427612e-08, 
    6.422655e-08, 6.441695e-08, 6.385987e-08, 6.40738e-08, 6.246512e-08, 
    6.247458e-08, 6.251866e-08, 6.232491e-08, 6.231306e-08, 6.213552e-08, 
    6.229349e-08, 6.236077e-08, 6.253156e-08, 6.263257e-08, 6.27286e-08, 
    6.293975e-08, 6.317556e-08, 6.350534e-08, 6.374228e-08, 6.390112e-08, 
    6.380372e-08, 6.388971e-08, 6.379359e-08, 6.374854e-08, 6.424895e-08, 
    6.396795e-08, 6.438957e-08, 6.436624e-08, 6.417542e-08, 6.436887e-08, 
    6.248122e-08, 6.242679e-08, 6.223777e-08, 6.238569e-08, 6.211619e-08, 
    6.226703e-08, 6.235377e-08, 6.268847e-08, 6.276202e-08, 6.283021e-08, 
    6.296489e-08, 6.313774e-08, 6.344097e-08, 6.370482e-08, 6.394571e-08, 
    6.392806e-08, 6.393427e-08, 6.398808e-08, 6.385479e-08, 6.400997e-08, 
    6.403601e-08, 6.396792e-08, 6.436311e-08, 6.425022e-08, 6.436574e-08, 
    6.429224e-08, 6.244449e-08, 6.253608e-08, 6.248658e-08, 6.257967e-08, 
    6.251409e-08, 6.280568e-08, 6.289311e-08, 6.330224e-08, 6.313434e-08, 
    6.340156e-08, 6.316149e-08, 6.320403e-08, 6.341026e-08, 6.317446e-08, 
    6.369027e-08, 6.334054e-08, 6.399017e-08, 6.36409e-08, 6.401206e-08, 
    6.394467e-08, 6.405626e-08, 6.415619e-08, 6.428195e-08, 6.451393e-08, 
    6.446022e-08, 6.465423e-08, 6.267265e-08, 6.279146e-08, 6.278102e-08, 
    6.290536e-08, 6.299733e-08, 6.319667e-08, 6.35164e-08, 6.339616e-08, 
    6.361689e-08, 6.366121e-08, 6.332587e-08, 6.353175e-08, 6.2871e-08, 
    6.297773e-08, 6.291419e-08, 6.268202e-08, 6.342385e-08, 6.304312e-08, 
    6.37462e-08, 6.353994e-08, 6.414194e-08, 6.384253e-08, 6.443064e-08, 
    6.468203e-08, 6.491868e-08, 6.51952e-08, 6.285632e-08, 6.277559e-08, 
    6.292016e-08, 6.312016e-08, 6.330577e-08, 6.355251e-08, 6.357777e-08, 
    6.362399e-08, 6.374373e-08, 6.384442e-08, 6.363859e-08, 6.386966e-08, 
    6.300247e-08, 6.345691e-08, 6.274506e-08, 6.295939e-08, 6.310837e-08, 
    6.304303e-08, 6.338242e-08, 6.346242e-08, 6.378748e-08, 6.361945e-08, 
    6.461998e-08, 6.417729e-08, 6.540579e-08, 6.506244e-08, 6.274738e-08, 
    6.285605e-08, 6.323427e-08, 6.305431e-08, 6.356899e-08, 6.369568e-08, 
    6.379868e-08, 6.393034e-08, 6.394456e-08, 6.402257e-08, 6.389474e-08, 
    6.401752e-08, 6.355304e-08, 6.37606e-08, 6.319105e-08, 6.332966e-08, 
    6.326589e-08, 6.319594e-08, 6.341183e-08, 6.364183e-08, 6.364677e-08, 
    6.372051e-08, 6.392831e-08, 6.357108e-08, 6.467708e-08, 6.399399e-08, 
    6.297455e-08, 6.318386e-08, 6.321378e-08, 6.313269e-08, 6.368298e-08, 
    6.348358e-08, 6.402067e-08, 6.387551e-08, 6.411335e-08, 6.399516e-08, 
    6.397777e-08, 6.382598e-08, 6.373148e-08, 6.349272e-08, 6.329847e-08, 
    6.314445e-08, 6.318027e-08, 6.334945e-08, 6.365591e-08, 6.394584e-08, 
    6.388233e-08, 6.409527e-08, 6.353167e-08, 6.376798e-08, 6.367664e-08, 
    6.391483e-08, 6.339297e-08, 6.383731e-08, 6.327939e-08, 6.332831e-08, 
    6.347963e-08, 6.378401e-08, 6.385137e-08, 6.392327e-08, 6.387891e-08, 
    6.366369e-08, 6.362843e-08, 6.347595e-08, 6.343384e-08, 6.331766e-08, 
    6.322146e-08, 6.330935e-08, 6.340164e-08, 6.366378e-08, 6.390003e-08, 
    6.415761e-08, 6.422066e-08, 6.452161e-08, 6.427662e-08, 6.468089e-08, 
    6.433715e-08, 6.493221e-08, 6.386308e-08, 6.432707e-08, 6.348652e-08, 
    6.357706e-08, 6.374083e-08, 6.41165e-08, 6.39137e-08, 6.415087e-08, 
    6.362706e-08, 6.335529e-08, 6.328499e-08, 6.315381e-08, 6.328799e-08, 
    6.327708e-08, 6.340547e-08, 6.336422e-08, 6.367249e-08, 6.35069e-08, 
    6.397733e-08, 6.414901e-08, 6.463389e-08, 6.493114e-08, 6.523376e-08, 
    6.536735e-08, 6.540802e-08, 6.542501e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.3407073, -0.340712, -0.3407111, -0.3407148, -0.3407128, -0.3407151, 
    -0.3407083, -0.3407121, -0.3407097, -0.3407078, -0.3407218, -0.3407149, 
    -0.3407294, -0.3407249, -0.3407526, -0.3407286, -0.3407542, -0.3407525, 
    -0.3407578, -0.3407563, -0.3409147, -0.3407585, -0.340919, -0.3409134, 
    -0.3409142, -0.3407584, -0.3407164, -0.3407209, -0.3407161, -0.3407168, 
    -0.3407165, -0.3407128, -0.3407108, -0.340707, -0.3407077, -0.3407106, 
    -0.3407171, -0.3407149, -0.3407205, -0.3407204, -0.3407266, -0.3407238, 
    -0.3407343, -0.3407313, -0.3407564, -0.3407542, -0.3407562, -0.3407556, 
    -0.3407563, -0.340753, -0.3407544, -0.3407352, -0.3407243, -0.3407275, 
    -0.3407179, -0.3407121, -0.3407085, -0.3407058, -0.3407062, -0.3407069, 
    -0.3407106, -0.3407141, -0.3407168, -0.3407186, -0.3407204, -0.3407255, 
    -0.3407284, -0.3407348, -0.3407338, -0.3407356, -0.3407539, -0.3407571, 
    -0.3407566, -0.3407579, -0.3407356, -0.3407559, -0.3407331, -0.3407349, 
    -0.3407205, -0.3407155, -0.3407131, -0.3407112, -0.3407065, -0.3407097, 
    -0.3407084, -0.3407116, -0.3407136, -0.3407126, -0.3407187, -0.3407163, 
    -0.3407286, -0.3407233, -0.3407537, -0.340734, -0.3407545, -0.340736, 
    -0.340756, -0.3407528, -0.3407585, -0.3409104, -0.3407588, -0.3409137, 
    -0.3407526, -0.3407562, -0.3407126, -0.3407127, -0.3407135, -0.3407102, 
    -0.34071, -0.340707, -0.3407097, -0.3407108, -0.3407137, -0.3407154, 
    -0.340717, -0.3407206, -0.3407245, -0.3407301, -0.3407342, -0.3407533, 
    -0.3407353, -0.3407531, -0.3407351, -0.3407343, -0.3409097, -0.3407544, 
    -0.3409131, -0.3409126, -0.340758, -0.3409126, -0.3407128, -0.340712, 
    -0.3407087, -0.3407112, -0.3407067, -0.3407092, -0.3407106, -0.3407163, 
    -0.3407176, -0.3407187, -0.340721, -0.3407239, -0.340729, -0.3407335, 
    -0.3407541, -0.3407538, -0.3407539, -0.3407548, -0.3407525, -0.3407552, 
    -0.3407556, -0.3407544, -0.3409125, -0.3409098, -0.3409125, -0.3409109, 
    -0.3407122, -0.3407138, -0.3407129, -0.3407145, -0.3407134, -0.3407182, 
    -0.3407197, -0.3407266, -0.3407238, -0.3407283, -0.3407243, -0.340725, 
    -0.3407284, -0.3407246, -0.3407332, -0.3407272, -0.3407548, -0.3407323, 
    -0.3407552, -0.3407541, -0.340756, -0.3407576, -0.3409106, -0.3409157, 
    -0.3409145, -0.3409186, -0.3407161, -0.340718, -0.3407179, -0.34072, 
    -0.3407215, -0.3407249, -0.3407303, -0.3407283, -0.3407321, -0.3407328, 
    -0.3407272, -0.3407306, -0.3407194, -0.3407211, -0.3407201, -0.3407162, 
    -0.3407287, -0.3407222, -0.3407342, -0.3407308, -0.3407574, -0.3407358, 
    -0.3409139, -0.340919, -0.3409241, -0.3409294, -0.3407192, -0.3407178, 
    -0.3407203, -0.3407235, -0.3407268, -0.340731, -0.3407314, -0.3407322, 
    -0.3407342, -0.3407359, -0.3407324, -0.3407528, -0.3407214, -0.3407293, 
    -0.3407173, -0.3407208, -0.3407234, -0.3407223, -0.3407281, -0.3407294, 
    -0.3407349, -0.3407321, -0.3409177, -0.3407579, -0.3409337, -0.3409268, 
    -0.3407173, -0.3407192, -0.3407255, -0.3407225, -0.3407313, -0.3407334, 
    -0.3407352, -0.3407538, -0.340754, -0.3407553, -0.3407532, -0.3407553, 
    -0.340731, -0.3407345, -0.3407249, -0.3407272, -0.3407261, -0.3407249, 
    -0.3407286, -0.3407324, -0.3407326, -0.3407338, -0.3407534, -0.3407313, 
    -0.3409187, -0.3407546, -0.3407212, -0.3407246, -0.3407252, -0.3407239, 
    -0.3407332, -0.3407298, -0.3407553, -0.3407529, -0.3407569, -0.3407549, 
    -0.3407546, -0.3407356, -0.340734, -0.3407299, -0.3407266, -0.3407241, 
    -0.3407247, -0.3407275, -0.3407327, -0.340754, -0.3407529, -0.3407566, 
    -0.3407306, -0.3407346, -0.340733, -0.3407535, -0.3407283, -0.3407355, 
    -0.3407264, -0.3407272, -0.3407297, -0.3407348, -0.3407524, -0.3407536, 
    -0.3407529, -0.3407328, -0.3407322, -0.3407297, -0.3407289, -0.340727, 
    -0.3407254, -0.3407269, -0.3407284, -0.3407328, -0.3407532, -0.3407577, 
    -0.3407588, -0.3409156, -0.3409102, -0.3409187, -0.3409114, -0.340924, 
    -0.3407525, -0.3409114, -0.3407299, -0.3407314, -0.3407341, -0.3407569, 
    -0.3407535, -0.3407575, -0.3407322, -0.3407275, -0.3407264, -0.3407242, 
    -0.3407265, -0.3407263, -0.3407285, -0.3407278, -0.340733, -0.3407302, 
    -0.3407546, -0.3407575, -0.3409182, -0.3409242, -0.3409304, -0.340933, 
    -0.3409338, -0.3409342 ;

 TAUY =
  -0.3407073, -0.340712, -0.3407111, -0.3407148, -0.3407128, -0.3407151, 
    -0.3407083, -0.3407121, -0.3407097, -0.3407078, -0.3407218, -0.3407149, 
    -0.3407294, -0.3407249, -0.3407526, -0.3407286, -0.3407542, -0.3407525, 
    -0.3407578, -0.3407563, -0.3409147, -0.3407585, -0.340919, -0.3409134, 
    -0.3409142, -0.3407584, -0.3407164, -0.3407209, -0.3407161, -0.3407168, 
    -0.3407165, -0.3407128, -0.3407108, -0.340707, -0.3407077, -0.3407106, 
    -0.3407171, -0.3407149, -0.3407205, -0.3407204, -0.3407266, -0.3407238, 
    -0.3407343, -0.3407313, -0.3407564, -0.3407542, -0.3407562, -0.3407556, 
    -0.3407563, -0.340753, -0.3407544, -0.3407352, -0.3407243, -0.3407275, 
    -0.3407179, -0.3407121, -0.3407085, -0.3407058, -0.3407062, -0.3407069, 
    -0.3407106, -0.3407141, -0.3407168, -0.3407186, -0.3407204, -0.3407255, 
    -0.3407284, -0.3407348, -0.3407338, -0.3407356, -0.3407539, -0.3407571, 
    -0.3407566, -0.3407579, -0.3407356, -0.3407559, -0.3407331, -0.3407349, 
    -0.3407205, -0.3407155, -0.3407131, -0.3407112, -0.3407065, -0.3407097, 
    -0.3407084, -0.3407116, -0.3407136, -0.3407126, -0.3407187, -0.3407163, 
    -0.3407286, -0.3407233, -0.3407537, -0.340734, -0.3407545, -0.340736, 
    -0.340756, -0.3407528, -0.3407585, -0.3409104, -0.3407588, -0.3409137, 
    -0.3407526, -0.3407562, -0.3407126, -0.3407127, -0.3407135, -0.3407102, 
    -0.34071, -0.340707, -0.3407097, -0.3407108, -0.3407137, -0.3407154, 
    -0.340717, -0.3407206, -0.3407245, -0.3407301, -0.3407342, -0.3407533, 
    -0.3407353, -0.3407531, -0.3407351, -0.3407343, -0.3409097, -0.3407544, 
    -0.3409131, -0.3409126, -0.340758, -0.3409126, -0.3407128, -0.340712, 
    -0.3407087, -0.3407112, -0.3407067, -0.3407092, -0.3407106, -0.3407163, 
    -0.3407176, -0.3407187, -0.340721, -0.3407239, -0.340729, -0.3407335, 
    -0.3407541, -0.3407538, -0.3407539, -0.3407548, -0.3407525, -0.3407552, 
    -0.3407556, -0.3407544, -0.3409125, -0.3409098, -0.3409125, -0.3409109, 
    -0.3407122, -0.3407138, -0.3407129, -0.3407145, -0.3407134, -0.3407182, 
    -0.3407197, -0.3407266, -0.3407238, -0.3407283, -0.3407243, -0.340725, 
    -0.3407284, -0.3407246, -0.3407332, -0.3407272, -0.3407548, -0.3407323, 
    -0.3407552, -0.3407541, -0.340756, -0.3407576, -0.3409106, -0.3409157, 
    -0.3409145, -0.3409186, -0.3407161, -0.340718, -0.3407179, -0.34072, 
    -0.3407215, -0.3407249, -0.3407303, -0.3407283, -0.3407321, -0.3407328, 
    -0.3407272, -0.3407306, -0.3407194, -0.3407211, -0.3407201, -0.3407162, 
    -0.3407287, -0.3407222, -0.3407342, -0.3407308, -0.3407574, -0.3407358, 
    -0.3409139, -0.340919, -0.3409241, -0.3409294, -0.3407192, -0.3407178, 
    -0.3407203, -0.3407235, -0.3407268, -0.340731, -0.3407314, -0.3407322, 
    -0.3407342, -0.3407359, -0.3407324, -0.3407528, -0.3407214, -0.3407293, 
    -0.3407173, -0.3407208, -0.3407234, -0.3407223, -0.3407281, -0.3407294, 
    -0.3407349, -0.3407321, -0.3409177, -0.3407579, -0.3409337, -0.3409268, 
    -0.3407173, -0.3407192, -0.3407255, -0.3407225, -0.3407313, -0.3407334, 
    -0.3407352, -0.3407538, -0.340754, -0.3407553, -0.3407532, -0.3407553, 
    -0.340731, -0.3407345, -0.3407249, -0.3407272, -0.3407261, -0.3407249, 
    -0.3407286, -0.3407324, -0.3407326, -0.3407338, -0.3407534, -0.3407313, 
    -0.3409187, -0.3407546, -0.3407212, -0.3407246, -0.3407252, -0.3407239, 
    -0.3407332, -0.3407298, -0.3407553, -0.3407529, -0.3407569, -0.3407549, 
    -0.3407546, -0.3407356, -0.340734, -0.3407299, -0.3407266, -0.3407241, 
    -0.3407247, -0.3407275, -0.3407327, -0.340754, -0.3407529, -0.3407566, 
    -0.3407306, -0.3407346, -0.340733, -0.3407535, -0.3407283, -0.3407355, 
    -0.3407264, -0.3407272, -0.3407297, -0.3407348, -0.3407524, -0.3407536, 
    -0.3407529, -0.3407328, -0.3407322, -0.3407297, -0.3407289, -0.340727, 
    -0.3407254, -0.3407269, -0.3407284, -0.3407328, -0.3407532, -0.3407577, 
    -0.3407588, -0.3409156, -0.3409102, -0.3409187, -0.3409114, -0.340924, 
    -0.3407525, -0.3409114, -0.3407299, -0.3407314, -0.3407341, -0.3407569, 
    -0.3407535, -0.3407575, -0.3407322, -0.3407275, -0.3407264, -0.3407242, 
    -0.3407265, -0.3407263, -0.3407285, -0.3407278, -0.340733, -0.3407302, 
    -0.3407546, -0.3407575, -0.3409182, -0.3409242, -0.3409304, -0.340933, 
    -0.3409338, -0.3409342 ;

 TBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.4824, 261.5035, 261.4994, 261.5163, 261.5069, 261.518, 261.4867, 
    261.5043, 261.4931, 261.4843, 261.5492, 261.5171, 261.5826, 261.5621, 
    261.6134, 261.5794, 261.6203, 261.6125, 261.6361, 261.6294, 261.6566, 
    261.6393, 261.6723, 261.6518, 261.655, 261.6386, 261.5236, 261.5452, 
    261.5223, 261.5254, 261.524, 261.5071, 261.4986, 261.4808, 261.4841, 
    261.4971, 261.5268, 261.5167, 261.5421, 261.5415, 261.5697, 261.5569, 
    261.6043, 261.5909, 261.6296, 261.6199, 261.6292, 261.6264, 261.6292, 
    261.6149, 261.621, 261.6085, 261.5593, 261.5738, 261.5307, 261.5047, 
    261.4875, 261.4753, 261.477, 261.4803, 261.4972, 261.5132, 261.5253, 
    261.5334, 261.5414, 261.5656, 261.5784, 261.607, 261.6019, 261.6106, 
    261.6189, 261.6329, 261.6306, 261.6368, 261.6104, 261.6279, 261.5989, 
    261.6069, 261.5435, 261.5194, 261.5091, 261.5002, 261.4783, 261.4934, 
    261.4875, 261.5016, 261.5106, 261.5062, 261.5336, 261.5229, 261.5791, 
    261.5549, 261.6179, 261.6029, 261.6216, 261.6121, 261.6284, 261.6136, 
    261.6391, 261.6417, 261.6409, 261.6525, 261.6128, 261.6292, 261.506, 
    261.5068, 261.5101, 261.4953, 261.4944, 261.4807, 261.4929, 261.498, 
    261.5111, 261.5189, 261.5262, 261.5424, 261.5605, 261.5858, 261.6039, 
    261.616, 261.6086, 261.6151, 261.6078, 261.6044, 261.6396, 261.6211, 
    261.6504, 261.6486, 261.637, 261.6488, 261.5073, 261.5031, 261.4886, 
    261.4999, 261.4793, 261.4908, 261.4975, 261.5232, 261.5288, 261.534, 
    261.5444, 261.5576, 261.5808, 261.601, 261.6194, 261.618, 261.6185, 
    261.6226, 261.6124, 261.6243, 261.6263, 261.6211, 261.6483, 261.6397, 
    261.6486, 261.6429, 261.5045, 261.5115, 261.5077, 261.5148, 261.5098, 
    261.5321, 261.5388, 261.5702, 261.5573, 261.5778, 261.5594, 261.5627, 
    261.5785, 261.5604, 261.5999, 261.5731, 261.6228, 261.5961, 261.6245, 
    261.6193, 261.6278, 261.6355, 261.6422, 261.6599, 261.6558, 261.6706, 
    261.5219, 261.5311, 261.5303, 261.5398, 261.5468, 261.5621, 261.5866, 
    261.5774, 261.5943, 261.5977, 261.572, 261.5878, 261.5372, 261.5453, 
    261.5405, 261.5227, 261.5795, 261.5504, 261.6042, 261.5884, 261.6344, 
    261.6116, 261.6535, 261.6727, 261.6908, 261.7118, 261.536, 261.5298, 
    261.5409, 261.5562, 261.5705, 261.5894, 261.5913, 261.5948, 261.604, 
    261.6117, 261.5959, 261.6136, 261.5472, 261.5821, 261.5275, 261.5439, 
    261.5554, 261.5504, 261.5764, 261.5825, 261.6074, 261.5945, 261.6679, 
    261.6371, 261.7279, 261.7017, 261.5277, 261.536, 261.565, 261.5512, 
    261.5906, 261.6003, 261.6082, 261.6182, 261.6193, 261.6253, 261.6155, 
    261.6249, 261.5894, 261.6053, 261.5617, 261.5723, 261.5674, 261.5621, 
    261.5786, 261.5962, 261.5966, 261.6022, 261.618, 261.5908, 261.6723, 
    261.623, 261.5451, 261.5611, 261.5634, 261.5572, 261.5994, 261.5841, 
    261.6251, 261.614, 261.6322, 261.6232, 261.6219, 261.6103, 261.6031, 
    261.5848, 261.5699, 261.5581, 261.5609, 261.5738, 261.5973, 261.6194, 
    261.6145, 261.6308, 261.5878, 261.6059, 261.5989, 261.617, 261.5771, 
    261.6111, 261.5685, 261.5722, 261.5838, 261.6071, 261.6122, 261.6177, 
    261.6143, 261.5979, 261.5952, 261.5835, 261.5803, 261.5714, 261.564, 
    261.5707, 261.5778, 261.5979, 261.6159, 261.6356, 261.6404, 261.6604, 
    261.6417, 261.6725, 261.6463, 261.6917, 261.613, 261.6456, 261.5843, 
    261.5912, 261.6038, 261.6324, 261.6169, 261.6351, 261.5951, 261.5742, 
    261.5689, 261.5588, 261.5691, 261.5683, 261.5781, 261.575, 261.5986, 
    261.5859, 261.6218, 261.6349, 261.669, 261.6917, 261.7148, 261.725, 
    261.7281, 261.7294 ;

 TG_R =
  261.4824, 261.5035, 261.4994, 261.5163, 261.5069, 261.518, 261.4867, 
    261.5043, 261.4931, 261.4843, 261.5492, 261.5171, 261.5826, 261.5621, 
    261.6134, 261.5794, 261.6203, 261.6125, 261.6361, 261.6294, 261.6566, 
    261.6393, 261.6723, 261.6518, 261.655, 261.6386, 261.5236, 261.5452, 
    261.5223, 261.5254, 261.524, 261.5071, 261.4986, 261.4808, 261.4841, 
    261.4971, 261.5268, 261.5167, 261.5421, 261.5415, 261.5697, 261.5569, 
    261.6043, 261.5909, 261.6296, 261.6199, 261.6292, 261.6264, 261.6292, 
    261.6149, 261.621, 261.6085, 261.5593, 261.5738, 261.5307, 261.5047, 
    261.4875, 261.4753, 261.477, 261.4803, 261.4972, 261.5132, 261.5253, 
    261.5334, 261.5414, 261.5656, 261.5784, 261.607, 261.6019, 261.6106, 
    261.6189, 261.6329, 261.6306, 261.6368, 261.6104, 261.6279, 261.5989, 
    261.6069, 261.5435, 261.5194, 261.5091, 261.5002, 261.4783, 261.4934, 
    261.4875, 261.5016, 261.5106, 261.5062, 261.5336, 261.5229, 261.5791, 
    261.5549, 261.6179, 261.6029, 261.6216, 261.6121, 261.6284, 261.6136, 
    261.6391, 261.6417, 261.6409, 261.6525, 261.6128, 261.6292, 261.506, 
    261.5068, 261.5101, 261.4953, 261.4944, 261.4807, 261.4929, 261.498, 
    261.5111, 261.5189, 261.5262, 261.5424, 261.5605, 261.5858, 261.6039, 
    261.616, 261.6086, 261.6151, 261.6078, 261.6044, 261.6396, 261.6211, 
    261.6504, 261.6486, 261.637, 261.6488, 261.5073, 261.5031, 261.4886, 
    261.4999, 261.4793, 261.4908, 261.4975, 261.5232, 261.5288, 261.534, 
    261.5444, 261.5576, 261.5808, 261.601, 261.6194, 261.618, 261.6185, 
    261.6226, 261.6124, 261.6243, 261.6263, 261.6211, 261.6483, 261.6397, 
    261.6486, 261.6429, 261.5045, 261.5115, 261.5077, 261.5148, 261.5098, 
    261.5321, 261.5388, 261.5702, 261.5573, 261.5778, 261.5594, 261.5627, 
    261.5785, 261.5604, 261.5999, 261.5731, 261.6228, 261.5961, 261.6245, 
    261.6193, 261.6278, 261.6355, 261.6422, 261.6599, 261.6558, 261.6706, 
    261.5219, 261.5311, 261.5303, 261.5398, 261.5468, 261.5621, 261.5866, 
    261.5774, 261.5943, 261.5977, 261.572, 261.5878, 261.5372, 261.5453, 
    261.5405, 261.5227, 261.5795, 261.5504, 261.6042, 261.5884, 261.6344, 
    261.6116, 261.6535, 261.6727, 261.6908, 261.7118, 261.536, 261.5298, 
    261.5409, 261.5562, 261.5705, 261.5894, 261.5913, 261.5948, 261.604, 
    261.6117, 261.5959, 261.6136, 261.5472, 261.5821, 261.5275, 261.5439, 
    261.5554, 261.5504, 261.5764, 261.5825, 261.6074, 261.5945, 261.6679, 
    261.6371, 261.7279, 261.7017, 261.5277, 261.536, 261.565, 261.5512, 
    261.5906, 261.6003, 261.6082, 261.6182, 261.6193, 261.6253, 261.6155, 
    261.6249, 261.5894, 261.6053, 261.5617, 261.5723, 261.5674, 261.5621, 
    261.5786, 261.5962, 261.5966, 261.6022, 261.618, 261.5908, 261.6723, 
    261.623, 261.5451, 261.5611, 261.5634, 261.5572, 261.5994, 261.5841, 
    261.6251, 261.614, 261.6322, 261.6232, 261.6219, 261.6103, 261.6031, 
    261.5848, 261.5699, 261.5581, 261.5609, 261.5738, 261.5973, 261.6194, 
    261.6145, 261.6308, 261.5878, 261.6059, 261.5989, 261.617, 261.5771, 
    261.6111, 261.5685, 261.5722, 261.5838, 261.6071, 261.6122, 261.6177, 
    261.6143, 261.5979, 261.5952, 261.5835, 261.5803, 261.5714, 261.564, 
    261.5707, 261.5778, 261.5979, 261.6159, 261.6356, 261.6404, 261.6604, 
    261.6417, 261.6725, 261.6463, 261.6917, 261.613, 261.6456, 261.5843, 
    261.5912, 261.6038, 261.6324, 261.6169, 261.6351, 261.5951, 261.5742, 
    261.5689, 261.5588, 261.5691, 261.5683, 261.5781, 261.575, 261.5986, 
    261.5859, 261.6218, 261.6349, 261.669, 261.6917, 261.7148, 261.725, 
    261.7281, 261.7294 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.6156, 254.6171, 254.6168, 254.618, 254.6174, 254.6182, 254.6159, 
    254.6172, 254.6164, 254.6157, 254.6204, 254.6181, 254.6229, 254.6214, 
    254.6252, 254.6227, 254.6257, 254.6251, 254.6269, 254.6264, 254.6282, 
    254.6271, 254.6294, 254.6279, 254.6281, 254.6271, 254.6186, 254.6201, 
    254.6185, 254.6187, 254.6186, 254.6174, 254.6167, 254.6155, 254.6157, 
    254.6167, 254.6188, 254.6181, 254.6199, 254.6199, 254.622, 254.621, 
    254.6245, 254.6235, 254.6264, 254.6257, 254.6264, 254.6262, 254.6264, 
    254.6253, 254.6258, 254.6248, 254.6212, 254.6223, 254.6191, 254.6172, 
    254.616, 254.6151, 254.6152, 254.6154, 254.6167, 254.6178, 254.6187, 
    254.6193, 254.6199, 254.6216, 254.6226, 254.6247, 254.6244, 254.625, 
    254.6256, 254.6267, 254.6265, 254.627, 254.625, 254.6263, 254.6241, 
    254.6247, 254.62, 254.6183, 254.6175, 254.6169, 254.6153, 254.6164, 
    254.6159, 254.617, 254.6176, 254.6173, 254.6193, 254.6185, 254.6227, 
    254.6209, 254.6255, 254.6244, 254.6258, 254.6251, 254.6263, 254.6252, 
    254.6271, 254.6272, 254.6272, 254.628, 254.6252, 254.6264, 254.6173, 
    254.6174, 254.6176, 254.6165, 254.6165, 254.6155, 254.6163, 254.6167, 
    254.6177, 254.6182, 254.6188, 254.62, 254.6213, 254.6232, 254.6245, 
    254.6254, 254.6249, 254.6254, 254.6248, 254.6245, 254.627, 254.6258, 
    254.6278, 254.6277, 254.627, 254.6277, 254.6174, 254.6171, 254.616, 
    254.6169, 254.6154, 254.6162, 254.6167, 254.6185, 254.619, 254.6194, 
    254.6201, 254.6211, 254.6228, 254.6243, 254.6257, 254.6256, 254.6256, 
    254.6259, 254.6251, 254.626, 254.6262, 254.6258, 254.6277, 254.627, 
    254.6277, 254.6273, 254.6172, 254.6177, 254.6174, 254.618, 254.6176, 
    254.6192, 254.6197, 254.622, 254.6211, 254.6226, 254.6212, 254.6215, 
    254.6226, 254.6213, 254.6242, 254.6222, 254.6259, 254.6239, 254.626, 
    254.6257, 254.6263, 254.6268, 254.6272, 254.6285, 254.6282, 254.6293, 
    254.6185, 254.6191, 254.6191, 254.6198, 254.6203, 254.6214, 254.6232, 
    254.6225, 254.6238, 254.624, 254.6221, 254.6233, 254.6196, 254.6202, 
    254.6198, 254.6185, 254.6227, 254.6205, 254.6245, 254.6234, 254.6268, 
    254.6251, 254.628, 254.6294, 254.6308, 254.6324, 254.6195, 254.619, 
    254.6199, 254.621, 254.622, 254.6234, 254.6236, 254.6238, 254.6245, 
    254.6251, 254.6239, 254.6252, 254.6203, 254.6229, 254.6189, 254.6201, 
    254.6209, 254.6205, 254.6225, 254.6229, 254.6248, 254.6238, 254.6291, 
    254.627, 254.6336, 254.6316, 254.6189, 254.6195, 254.6216, 254.6206, 
    254.6235, 254.6242, 254.6248, 254.6256, 254.6257, 254.6261, 254.6254, 
    254.6261, 254.6234, 254.6246, 254.6214, 254.6222, 254.6218, 254.6214, 
    254.6226, 254.6239, 254.624, 254.6244, 254.6255, 254.6235, 254.6294, 
    254.6259, 254.6202, 254.6213, 254.6215, 254.6211, 254.6242, 254.623, 
    254.6261, 254.6253, 254.6266, 254.6259, 254.6258, 254.625, 254.6244, 
    254.6231, 254.622, 254.6211, 254.6213, 254.6223, 254.624, 254.6257, 
    254.6253, 254.6265, 254.6233, 254.6246, 254.6241, 254.6255, 254.6225, 
    254.625, 254.6219, 254.6222, 254.623, 254.6247, 254.6251, 254.6255, 
    254.6253, 254.6241, 254.6239, 254.623, 254.6228, 254.6221, 254.6216, 
    254.6221, 254.6226, 254.6241, 254.6254, 254.6269, 254.6272, 254.6285, 
    254.6271, 254.6294, 254.6274, 254.6308, 254.6252, 254.6274, 254.6231, 
    254.6236, 254.6245, 254.6266, 254.6255, 254.6268, 254.6239, 254.6223, 
    254.6219, 254.6212, 254.6219, 254.6219, 254.6226, 254.6224, 254.6241, 
    254.6232, 254.6258, 254.6268, 254.6292, 254.6309, 254.6326, 254.6334, 
    254.6336, 254.6337 ;

 THBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24018, 18.24016, 18.24017, 18.24016, 18.24016, 18.24015, 18.24017, 
    18.24016, 18.24017, 18.24018, 18.24014, 18.24015, 18.24011, 18.24013, 
    18.2401, 18.24012, 18.24009, 18.2401, 18.24008, 18.24008, 18.24007, 
    18.24008, 18.24006, 18.24007, 18.24007, 18.24008, 18.24015, 18.24014, 
    18.24015, 18.24015, 18.24015, 18.24016, 18.24017, 18.24018, 18.24018, 
    18.24017, 18.24015, 18.24015, 18.24014, 18.24014, 18.24012, 18.24013, 
    18.2401, 18.24011, 18.24008, 18.24009, 18.24009, 18.24009, 18.24008, 
    18.24009, 18.24009, 18.2401, 18.24013, 18.24012, 18.24015, 18.24016, 
    18.24017, 18.24018, 18.24018, 18.24018, 18.24017, 18.24016, 18.24015, 
    18.24014, 18.24014, 18.24012, 18.24012, 18.2401, 18.2401, 18.2401, 
    18.24009, 18.24008, 18.24008, 18.24008, 18.2401, 18.24009, 18.2401, 
    18.2401, 18.24014, 18.24015, 18.24016, 18.24017, 18.24018, 18.24017, 
    18.24017, 18.24016, 18.24016, 18.24016, 18.24014, 18.24015, 18.24012, 
    18.24013, 18.24009, 18.2401, 18.24009, 18.2401, 18.24009, 18.2401, 
    18.24008, 18.24007, 18.24008, 18.24007, 18.2401, 18.24009, 18.24016, 
    18.24016, 18.24016, 18.24017, 18.24017, 18.24018, 18.24017, 18.24017, 
    18.24016, 18.24015, 18.24015, 18.24014, 18.24013, 18.24011, 18.2401, 
    18.24009, 18.2401, 18.24009, 18.2401, 18.2401, 18.24008, 18.24009, 
    18.24007, 18.24007, 18.24008, 18.24007, 18.24016, 18.24016, 18.24017, 
    18.24017, 18.24018, 18.24017, 18.24017, 18.24015, 18.24015, 18.24014, 
    18.24014, 18.24013, 18.24011, 18.2401, 18.24009, 18.24009, 18.24009, 
    18.24009, 18.2401, 18.24009, 18.24009, 18.24009, 18.24007, 18.24008, 
    18.24007, 18.24007, 18.24016, 18.24016, 18.24016, 18.24016, 18.24016, 
    18.24014, 18.24014, 18.24012, 18.24013, 18.24012, 18.24013, 18.24013, 
    18.24012, 18.24013, 18.2401, 18.24012, 18.24009, 18.2401, 18.24009, 
    18.24009, 18.24009, 18.24008, 18.24007, 18.24006, 18.24007, 18.24006, 
    18.24015, 18.24015, 18.24015, 18.24014, 18.24014, 18.24013, 18.24011, 
    18.24012, 18.24011, 18.2401, 18.24012, 18.24011, 18.24014, 18.24014, 
    18.24014, 18.24015, 18.24012, 18.24013, 18.2401, 18.24011, 18.24008, 
    18.2401, 18.24007, 18.24006, 18.24004, 18.24003, 18.24014, 18.24015, 
    18.24014, 18.24013, 18.24012, 18.24011, 18.24011, 18.24011, 18.2401, 
    18.2401, 18.2401, 18.2401, 18.24014, 18.24011, 18.24015, 18.24014, 
    18.24013, 18.24013, 18.24012, 18.24011, 18.2401, 18.24011, 18.24006, 
    18.24008, 18.24002, 18.24004, 18.24015, 18.24014, 18.24013, 18.24013, 
    18.24011, 18.2401, 18.2401, 18.24009, 18.24009, 18.24009, 18.24009, 
    18.24009, 18.24011, 18.2401, 18.24013, 18.24012, 18.24012, 18.24013, 
    18.24012, 18.2401, 18.2401, 18.2401, 18.24009, 18.24011, 18.24006, 
    18.24009, 18.24014, 18.24013, 18.24013, 18.24013, 18.2401, 18.24011, 
    18.24009, 18.24009, 18.24008, 18.24009, 18.24009, 18.2401, 18.2401, 
    18.24011, 18.24012, 18.24013, 18.24013, 18.24012, 18.2401, 18.24009, 
    18.24009, 18.24008, 18.24011, 18.2401, 18.2401, 18.24009, 18.24012, 
    18.2401, 18.24012, 18.24012, 18.24011, 18.2401, 18.2401, 18.24009, 
    18.24009, 18.2401, 18.24011, 18.24011, 18.24012, 18.24012, 18.24013, 
    18.24012, 18.24012, 18.2401, 18.24009, 18.24008, 18.24008, 18.24006, 
    18.24007, 18.24006, 18.24007, 18.24004, 18.2401, 18.24007, 18.24011, 
    18.24011, 18.2401, 18.24008, 18.24009, 18.24008, 18.24011, 18.24012, 
    18.24012, 18.24013, 18.24012, 18.24012, 18.24012, 18.24012, 18.2401, 
    18.24011, 18.24009, 18.24008, 18.24006, 18.24004, 18.24003, 18.24002, 
    18.24002, 18.24002 ;

 TOTCOLCH4 =
  1.442303e-05, 1.420776e-05, 1.424956e-05, 1.407628e-05, 1.417236e-05, 
    1.405896e-05, 1.437935e-05, 1.419921e-05, 1.431416e-05, 1.440364e-05, 
    1.374118e-05, 1.406856e-05, 1.340295e-05, 1.361046e-05, 1.309054e-05, 
    1.343518e-05, 1.302129e-05, 1.310048e-05, 1.286254e-05, 1.293061e-05, 
    1.262741e-05, 1.283115e-05, 1.247089e-05, 1.267605e-05, 1.264389e-05, 
    1.283788e-05, 1.400258e-05, 1.378184e-05, 1.401567e-05, 1.398415e-05, 
    1.39983e-05, 1.417037e-05, 1.425722e-05, 1.443953e-05, 1.440641e-05, 
    1.427253e-05, 1.396998e-05, 1.407256e-05, 1.381439e-05, 1.382021e-05, 
    1.353392e-05, 1.366285e-05, 1.318359e-05, 1.331944e-05, 1.292777e-05, 
    1.302602e-05, 1.293237e-05, 1.296075e-05, 1.2932e-05, 1.307617e-05, 
    1.301435e-05, 1.314138e-05, 1.363867e-05, 1.34921e-05, 1.393021e-05, 
    1.419496e-05, 1.437143e-05, 1.449689e-05, 1.447914e-05, 1.444531e-05, 
    1.427174e-05, 1.410895e-05, 1.398514e-05, 1.390243e-05, 1.382105e-05, 
    1.357522e-05, 1.344555e-05, 1.315615e-05, 1.32083e-05, 1.312e-05, 
    1.30358e-05, 1.289468e-05, 1.291789e-05, 1.285579e-05, 1.312235e-05, 
    1.294505e-05, 1.323802e-05, 1.315774e-05, 1.379883e-05, 1.404487e-05, 
    1.414962e-05, 1.424152e-05, 1.44655e-05, 1.431075e-05, 1.437171e-05, 
    1.422678e-05, 1.413482e-05, 1.418029e-05, 1.390017e-05, 1.400894e-05, 
    1.343788e-05, 1.368325e-05, 1.304561e-05, 1.319759e-05, 1.300925e-05, 
    1.310529e-05, 1.294082e-05, 1.308882e-05, 1.283271e-05, 1.277721e-05, 
    1.281509e-05, 1.26694e-05, 1.309703e-05, 1.293236e-05, 1.418156e-05, 
    1.417414e-05, 1.41396e-05, 1.429155e-05, 1.430086e-05, 1.444044e-05, 
    1.431624e-05, 1.426341e-05, 1.41295e-05, 1.40504e-05, 1.397529e-05, 
    1.381044e-05, 1.36268e-05, 1.337091e-05, 1.318773e-05, 1.306525e-05, 
    1.314033e-05, 1.307404e-05, 1.314815e-05, 1.318292e-05, 1.279804e-05, 
    1.301377e-05, 1.269035e-05, 1.27082e-05, 1.285431e-05, 1.270619e-05, 
    1.416894e-05, 1.421163e-05, 1.436003e-05, 1.424387e-05, 1.445565e-05, 
    1.433702e-05, 1.426888e-05, 1.400664e-05, 1.394918e-05, 1.389591e-05, 
    1.379085e-05, 1.365624e-05, 1.342078e-05, 1.321664e-05, 1.303091e-05, 
    1.30445e-05, 1.303971e-05, 1.299829e-05, 1.310095e-05, 1.298145e-05, 
    1.296141e-05, 1.301381e-05, 1.27106e-05, 1.279709e-05, 1.270859e-05, 
    1.276489e-05, 1.419775e-05, 1.412595e-05, 1.416474e-05, 1.409181e-05, 
    1.414317e-05, 1.391503e-05, 1.384678e-05, 1.352836e-05, 1.365888e-05, 
    1.345132e-05, 1.363777e-05, 1.360469e-05, 1.344451e-05, 1.362769e-05, 
    1.322786e-05, 1.349861e-05, 1.299668e-05, 1.326598e-05, 1.297984e-05, 
    1.303171e-05, 1.294586e-05, 1.286908e-05, 1.277277e-05, 1.259524e-05, 
    1.26363e-05, 1.248819e-05, 1.401904e-05, 1.392615e-05, 1.393434e-05, 
    1.383727e-05, 1.376556e-05, 1.361042e-05, 1.336237e-05, 1.345554e-05, 
    1.328462e-05, 1.325036e-05, 1.351008e-05, 1.335046e-05, 1.386407e-05, 
    1.378079e-05, 1.383037e-05, 1.40117e-05, 1.343403e-05, 1.372985e-05, 
    1.31847e-05, 1.334415e-05, 1.288002e-05, 1.311036e-05, 1.265892e-05, 
    1.246694e-05, 1.2287e-05, 1.20774e-05, 1.387553e-05, 1.393858e-05, 
    1.382574e-05, 1.366988e-05, 1.352566e-05, 1.333441e-05, 1.331488e-05, 
    1.327912e-05, 1.318662e-05, 1.310895e-05, 1.32678e-05, 1.30895e-05, 
    1.376145e-05, 1.340842e-05, 1.396242e-05, 1.379508e-05, 1.367907e-05, 
    1.372995e-05, 1.34662e-05, 1.340419e-05, 1.315283e-05, 1.328265e-05, 
    1.251424e-05, 1.285284e-05, 1.191848e-05, 1.21779e-05, 1.396062e-05, 
    1.387575e-05, 1.358118e-05, 1.372117e-05, 1.332167e-05, 1.322372e-05, 
    1.314422e-05, 1.304273e-05, 1.303179e-05, 1.297175e-05, 1.307017e-05, 
    1.297565e-05, 1.3334e-05, 1.31736e-05, 1.36148e-05, 1.350712e-05, 
    1.355664e-05, 1.361099e-05, 1.344339e-05, 1.326529e-05, 1.326153e-05, 
    1.320453e-05, 1.304414e-05, 1.332006e-05, 1.247062e-05, 1.299361e-05, 
    1.378332e-05, 1.362033e-05, 1.359712e-05, 1.366018e-05, 1.323353e-05, 
    1.338778e-05, 1.297322e-05, 1.308498e-05, 1.290199e-05, 1.299284e-05, 
    1.300622e-05, 1.312316e-05, 1.319608e-05, 1.338069e-05, 1.353132e-05, 
    1.365104e-05, 1.362318e-05, 1.349175e-05, 1.325442e-05, 1.303079e-05, 
    1.30797e-05, 1.291587e-05, 1.335055e-05, 1.316788e-05, 1.323841e-05, 
    1.305469e-05, 1.345801e-05, 1.311429e-05, 1.354616e-05, 1.350818e-05, 
    1.339085e-05, 1.315549e-05, 1.310359e-05, 1.304817e-05, 1.308236e-05, 
    1.324842e-05, 1.327568e-05, 1.33937e-05, 1.342631e-05, 1.351645e-05, 
    1.359116e-05, 1.352289e-05, 1.345127e-05, 1.324836e-05, 1.306607e-05, 
    1.286798e-05, 1.281962e-05, 1.25893e-05, 1.277678e-05, 1.246771e-05, 
    1.27303e-05, 1.227661e-05, 1.309448e-05, 1.27381e-05, 1.338552e-05, 
    1.331543e-05, 1.318882e-05, 1.289951e-05, 1.305555e-05, 1.287312e-05, 
    1.327675e-05, 1.34872e-05, 1.354181e-05, 1.364375e-05, 1.353948e-05, 
    1.354795e-05, 1.344833e-05, 1.348033e-05, 1.324164e-05, 1.336974e-05, 
    1.300655e-05, 1.287457e-05, 1.250368e-05, 1.227749e-05, 1.204832e-05, 
    1.194747e-05, 1.191682e-05, 1.190401e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24018, 18.24016, 18.24017, 18.24016, 18.24016, 18.24015, 18.24017, 
    18.24016, 18.24017, 18.24018, 18.24014, 18.24015, 18.24011, 18.24013, 
    18.2401, 18.24012, 18.24009, 18.2401, 18.24008, 18.24008, 18.24007, 
    18.24008, 18.24006, 18.24007, 18.24007, 18.24008, 18.24015, 18.24014, 
    18.24015, 18.24015, 18.24015, 18.24016, 18.24017, 18.24018, 18.24018, 
    18.24017, 18.24015, 18.24015, 18.24014, 18.24014, 18.24012, 18.24013, 
    18.2401, 18.24011, 18.24008, 18.24009, 18.24009, 18.24009, 18.24008, 
    18.24009, 18.24009, 18.2401, 18.24013, 18.24012, 18.24015, 18.24016, 
    18.24017, 18.24018, 18.24018, 18.24018, 18.24017, 18.24016, 18.24015, 
    18.24014, 18.24014, 18.24012, 18.24012, 18.2401, 18.2401, 18.2401, 
    18.24009, 18.24008, 18.24008, 18.24008, 18.2401, 18.24009, 18.2401, 
    18.2401, 18.24014, 18.24015, 18.24016, 18.24017, 18.24018, 18.24017, 
    18.24017, 18.24016, 18.24016, 18.24016, 18.24014, 18.24015, 18.24012, 
    18.24013, 18.24009, 18.2401, 18.24009, 18.2401, 18.24009, 18.2401, 
    18.24008, 18.24007, 18.24008, 18.24007, 18.2401, 18.24009, 18.24016, 
    18.24016, 18.24016, 18.24017, 18.24017, 18.24018, 18.24017, 18.24017, 
    18.24016, 18.24015, 18.24015, 18.24014, 18.24013, 18.24011, 18.2401, 
    18.24009, 18.2401, 18.24009, 18.2401, 18.2401, 18.24008, 18.24009, 
    18.24007, 18.24007, 18.24008, 18.24007, 18.24016, 18.24016, 18.24017, 
    18.24017, 18.24018, 18.24017, 18.24017, 18.24015, 18.24015, 18.24014, 
    18.24014, 18.24013, 18.24011, 18.2401, 18.24009, 18.24009, 18.24009, 
    18.24009, 18.2401, 18.24009, 18.24009, 18.24009, 18.24007, 18.24008, 
    18.24007, 18.24007, 18.24016, 18.24016, 18.24016, 18.24016, 18.24016, 
    18.24014, 18.24014, 18.24012, 18.24013, 18.24012, 18.24013, 18.24013, 
    18.24012, 18.24013, 18.2401, 18.24012, 18.24009, 18.2401, 18.24009, 
    18.24009, 18.24009, 18.24008, 18.24007, 18.24006, 18.24007, 18.24006, 
    18.24015, 18.24015, 18.24015, 18.24014, 18.24014, 18.24013, 18.24011, 
    18.24012, 18.24011, 18.2401, 18.24012, 18.24011, 18.24014, 18.24014, 
    18.24014, 18.24015, 18.24012, 18.24013, 18.2401, 18.24011, 18.24008, 
    18.2401, 18.24007, 18.24006, 18.24004, 18.24003, 18.24014, 18.24015, 
    18.24014, 18.24013, 18.24012, 18.24011, 18.24011, 18.24011, 18.2401, 
    18.2401, 18.2401, 18.2401, 18.24014, 18.24011, 18.24015, 18.24014, 
    18.24013, 18.24013, 18.24012, 18.24011, 18.2401, 18.24011, 18.24006, 
    18.24008, 18.24002, 18.24004, 18.24015, 18.24014, 18.24013, 18.24013, 
    18.24011, 18.2401, 18.2401, 18.24009, 18.24009, 18.24009, 18.24009, 
    18.24009, 18.24011, 18.2401, 18.24013, 18.24012, 18.24012, 18.24013, 
    18.24012, 18.2401, 18.2401, 18.2401, 18.24009, 18.24011, 18.24006, 
    18.24009, 18.24014, 18.24013, 18.24013, 18.24013, 18.2401, 18.24011, 
    18.24009, 18.24009, 18.24008, 18.24009, 18.24009, 18.2401, 18.2401, 
    18.24011, 18.24012, 18.24013, 18.24013, 18.24012, 18.2401, 18.24009, 
    18.24009, 18.24008, 18.24011, 18.2401, 18.2401, 18.24009, 18.24012, 
    18.2401, 18.24012, 18.24012, 18.24011, 18.2401, 18.2401, 18.24009, 
    18.24009, 18.2401, 18.24011, 18.24011, 18.24012, 18.24012, 18.24013, 
    18.24012, 18.24012, 18.2401, 18.24009, 18.24008, 18.24008, 18.24006, 
    18.24007, 18.24006, 18.24007, 18.24004, 18.2401, 18.24007, 18.24011, 
    18.24011, 18.2401, 18.24008, 18.24009, 18.24008, 18.24011, 18.24012, 
    18.24012, 18.24013, 18.24012, 18.24012, 18.24012, 18.24012, 18.2401, 
    18.24011, 18.24009, 18.24008, 18.24006, 18.24004, 18.24003, 18.24002, 
    18.24002, 18.24002 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.97623e-05, 5.976215e-05, 5.976218e-05, 5.976206e-05, 5.976213e-05, 
    5.976205e-05, 5.976227e-05, 5.976215e-05, 5.976223e-05, 5.976229e-05, 
    5.976183e-05, 5.976206e-05, 5.97616e-05, 5.976174e-05, 5.976138e-05, 
    5.976162e-05, 5.976133e-05, 5.976139e-05, 5.976122e-05, 5.976127e-05, 
    5.976106e-05, 5.97612e-05, 5.976095e-05, 5.976109e-05, 5.976107e-05, 
    5.97612e-05, 5.976201e-05, 5.976186e-05, 5.976202e-05, 5.9762e-05, 
    5.976201e-05, 5.976213e-05, 5.976219e-05, 5.976231e-05, 5.976229e-05, 
    5.97622e-05, 5.976199e-05, 5.976206e-05, 5.976188e-05, 5.976189e-05, 
    5.976169e-05, 5.976178e-05, 5.976145e-05, 5.976154e-05, 5.976127e-05, 
    5.976134e-05, 5.976127e-05, 5.976129e-05, 5.976127e-05, 5.976137e-05, 
    5.976133e-05, 5.976142e-05, 5.976176e-05, 5.976166e-05, 5.976196e-05, 
    5.976215e-05, 5.976227e-05, 5.976235e-05, 5.976234e-05, 5.976232e-05, 
    5.97622e-05, 5.976209e-05, 5.9762e-05, 5.976194e-05, 5.976189e-05, 
    5.976172e-05, 5.976163e-05, 5.976143e-05, 5.976146e-05, 5.97614e-05, 
    5.976134e-05, 5.976124e-05, 5.976126e-05, 5.976122e-05, 5.97614e-05, 
    5.976128e-05, 5.976148e-05, 5.976143e-05, 5.976187e-05, 5.976204e-05, 
    5.976211e-05, 5.976218e-05, 5.976233e-05, 5.976223e-05, 5.976227e-05, 
    5.976217e-05, 5.97621e-05, 5.976214e-05, 5.976194e-05, 5.976202e-05, 
    5.976162e-05, 5.976179e-05, 5.976135e-05, 5.976145e-05, 5.976132e-05, 
    5.976139e-05, 5.976127e-05, 5.976138e-05, 5.97612e-05, 5.976116e-05, 
    5.976119e-05, 5.976109e-05, 5.976138e-05, 5.976127e-05, 5.976214e-05, 
    5.976213e-05, 5.976211e-05, 5.976221e-05, 5.976222e-05, 5.976231e-05, 
    5.976223e-05, 5.976219e-05, 5.97621e-05, 5.976205e-05, 5.976199e-05, 
    5.976188e-05, 5.976175e-05, 5.976158e-05, 5.976145e-05, 5.976136e-05, 
    5.976141e-05, 5.976137e-05, 5.976142e-05, 5.976145e-05, 5.976118e-05, 
    5.976133e-05, 5.97611e-05, 5.976111e-05, 5.976122e-05, 5.976111e-05, 
    5.976213e-05, 5.976216e-05, 5.976226e-05, 5.976218e-05, 5.976233e-05, 
    5.976225e-05, 5.97622e-05, 5.976202e-05, 5.976198e-05, 5.976194e-05, 
    5.976187e-05, 5.976177e-05, 5.976161e-05, 5.976147e-05, 5.976134e-05, 
    5.976135e-05, 5.976134e-05, 5.976131e-05, 5.976139e-05, 5.97613e-05, 
    5.976129e-05, 5.976133e-05, 5.976111e-05, 5.976117e-05, 5.976111e-05, 
    5.976115e-05, 5.976215e-05, 5.97621e-05, 5.976213e-05, 5.976207e-05, 
    5.976211e-05, 5.976195e-05, 5.97619e-05, 5.976169e-05, 5.976178e-05, 
    5.976163e-05, 5.976176e-05, 5.976174e-05, 5.976163e-05, 5.976175e-05, 
    5.976147e-05, 5.976166e-05, 5.976131e-05, 5.97615e-05, 5.97613e-05, 
    5.976134e-05, 5.976128e-05, 5.976122e-05, 5.976116e-05, 5.976103e-05, 
    5.976106e-05, 5.976096e-05, 5.976202e-05, 5.976196e-05, 5.976197e-05, 
    5.97619e-05, 5.976185e-05, 5.976174e-05, 5.976157e-05, 5.976163e-05, 
    5.976151e-05, 5.976149e-05, 5.976167e-05, 5.976156e-05, 5.976192e-05, 
    5.976186e-05, 5.976189e-05, 5.976202e-05, 5.976162e-05, 5.976182e-05, 
    5.976145e-05, 5.976156e-05, 5.976123e-05, 5.976139e-05, 5.976108e-05, 
    5.976094e-05, 5.976082e-05, 5.976067e-05, 5.976193e-05, 5.976197e-05, 
    5.976189e-05, 5.976178e-05, 5.976168e-05, 5.976155e-05, 5.976154e-05, 
    5.976151e-05, 5.976145e-05, 5.976139e-05, 5.97615e-05, 5.976138e-05, 
    5.976185e-05, 5.97616e-05, 5.976198e-05, 5.976187e-05, 5.976179e-05, 
    5.976182e-05, 5.976164e-05, 5.97616e-05, 5.976142e-05, 5.976151e-05, 
    5.976098e-05, 5.976121e-05, 5.976055e-05, 5.976074e-05, 5.976198e-05, 
    5.976193e-05, 5.976172e-05, 5.976182e-05, 5.976154e-05, 5.976147e-05, 
    5.976142e-05, 5.976135e-05, 5.976134e-05, 5.97613e-05, 5.976137e-05, 
    5.97613e-05, 5.976155e-05, 5.976144e-05, 5.976174e-05, 5.976167e-05, 
    5.97617e-05, 5.976174e-05, 5.976163e-05, 5.97615e-05, 5.97615e-05, 
    5.976146e-05, 5.976135e-05, 5.976154e-05, 5.976095e-05, 5.976131e-05, 
    5.976186e-05, 5.976175e-05, 5.976173e-05, 5.976178e-05, 5.976148e-05, 
    5.976159e-05, 5.97613e-05, 5.976138e-05, 5.976125e-05, 5.976131e-05, 
    5.976132e-05, 5.97614e-05, 5.976145e-05, 5.976158e-05, 5.976169e-05, 
    5.976177e-05, 5.976175e-05, 5.976166e-05, 5.976149e-05, 5.976134e-05, 
    5.976137e-05, 5.976126e-05, 5.976156e-05, 5.976143e-05, 5.976148e-05, 
    5.976135e-05, 5.976163e-05, 5.97614e-05, 5.97617e-05, 5.976167e-05, 
    5.976159e-05, 5.976142e-05, 5.976139e-05, 5.976135e-05, 5.976137e-05, 
    5.976149e-05, 5.976151e-05, 5.976159e-05, 5.976161e-05, 5.976167e-05, 
    5.976173e-05, 5.976168e-05, 5.976163e-05, 5.976149e-05, 5.976136e-05, 
    5.976122e-05, 5.976119e-05, 5.976103e-05, 5.976116e-05, 5.976094e-05, 
    5.976113e-05, 5.976081e-05, 5.976138e-05, 5.976113e-05, 5.976158e-05, 
    5.976154e-05, 5.976145e-05, 5.976125e-05, 5.976135e-05, 5.976123e-05, 
    5.976151e-05, 5.976166e-05, 5.976169e-05, 5.976177e-05, 5.976169e-05, 
    5.97617e-05, 5.976163e-05, 5.976165e-05, 5.976149e-05, 5.976157e-05, 
    5.976132e-05, 5.976123e-05, 5.976097e-05, 5.976081e-05, 5.976065e-05, 
    5.976058e-05, 5.976055e-05, 5.976054e-05 ;

 TOTLITC_1m =
  5.97623e-05, 5.976215e-05, 5.976218e-05, 5.976206e-05, 5.976213e-05, 
    5.976205e-05, 5.976227e-05, 5.976215e-05, 5.976223e-05, 5.976229e-05, 
    5.976183e-05, 5.976206e-05, 5.97616e-05, 5.976174e-05, 5.976138e-05, 
    5.976162e-05, 5.976133e-05, 5.976139e-05, 5.976122e-05, 5.976127e-05, 
    5.976106e-05, 5.97612e-05, 5.976095e-05, 5.976109e-05, 5.976107e-05, 
    5.97612e-05, 5.976201e-05, 5.976186e-05, 5.976202e-05, 5.9762e-05, 
    5.976201e-05, 5.976213e-05, 5.976219e-05, 5.976231e-05, 5.976229e-05, 
    5.97622e-05, 5.976199e-05, 5.976206e-05, 5.976188e-05, 5.976189e-05, 
    5.976169e-05, 5.976178e-05, 5.976145e-05, 5.976154e-05, 5.976127e-05, 
    5.976134e-05, 5.976127e-05, 5.976129e-05, 5.976127e-05, 5.976137e-05, 
    5.976133e-05, 5.976142e-05, 5.976176e-05, 5.976166e-05, 5.976196e-05, 
    5.976215e-05, 5.976227e-05, 5.976235e-05, 5.976234e-05, 5.976232e-05, 
    5.97622e-05, 5.976209e-05, 5.9762e-05, 5.976194e-05, 5.976189e-05, 
    5.976172e-05, 5.976163e-05, 5.976143e-05, 5.976146e-05, 5.97614e-05, 
    5.976134e-05, 5.976124e-05, 5.976126e-05, 5.976122e-05, 5.97614e-05, 
    5.976128e-05, 5.976148e-05, 5.976143e-05, 5.976187e-05, 5.976204e-05, 
    5.976211e-05, 5.976218e-05, 5.976233e-05, 5.976223e-05, 5.976227e-05, 
    5.976217e-05, 5.97621e-05, 5.976214e-05, 5.976194e-05, 5.976202e-05, 
    5.976162e-05, 5.976179e-05, 5.976135e-05, 5.976145e-05, 5.976132e-05, 
    5.976139e-05, 5.976127e-05, 5.976138e-05, 5.97612e-05, 5.976116e-05, 
    5.976119e-05, 5.976109e-05, 5.976138e-05, 5.976127e-05, 5.976214e-05, 
    5.976213e-05, 5.976211e-05, 5.976221e-05, 5.976222e-05, 5.976231e-05, 
    5.976223e-05, 5.976219e-05, 5.97621e-05, 5.976205e-05, 5.976199e-05, 
    5.976188e-05, 5.976175e-05, 5.976158e-05, 5.976145e-05, 5.976136e-05, 
    5.976141e-05, 5.976137e-05, 5.976142e-05, 5.976145e-05, 5.976118e-05, 
    5.976133e-05, 5.97611e-05, 5.976111e-05, 5.976122e-05, 5.976111e-05, 
    5.976213e-05, 5.976216e-05, 5.976226e-05, 5.976218e-05, 5.976233e-05, 
    5.976225e-05, 5.97622e-05, 5.976202e-05, 5.976198e-05, 5.976194e-05, 
    5.976187e-05, 5.976177e-05, 5.976161e-05, 5.976147e-05, 5.976134e-05, 
    5.976135e-05, 5.976134e-05, 5.976131e-05, 5.976139e-05, 5.97613e-05, 
    5.976129e-05, 5.976133e-05, 5.976111e-05, 5.976117e-05, 5.976111e-05, 
    5.976115e-05, 5.976215e-05, 5.97621e-05, 5.976213e-05, 5.976207e-05, 
    5.976211e-05, 5.976195e-05, 5.97619e-05, 5.976169e-05, 5.976178e-05, 
    5.976163e-05, 5.976176e-05, 5.976174e-05, 5.976163e-05, 5.976175e-05, 
    5.976147e-05, 5.976166e-05, 5.976131e-05, 5.97615e-05, 5.97613e-05, 
    5.976134e-05, 5.976128e-05, 5.976122e-05, 5.976116e-05, 5.976103e-05, 
    5.976106e-05, 5.976096e-05, 5.976202e-05, 5.976196e-05, 5.976197e-05, 
    5.97619e-05, 5.976185e-05, 5.976174e-05, 5.976157e-05, 5.976163e-05, 
    5.976151e-05, 5.976149e-05, 5.976167e-05, 5.976156e-05, 5.976192e-05, 
    5.976186e-05, 5.976189e-05, 5.976202e-05, 5.976162e-05, 5.976182e-05, 
    5.976145e-05, 5.976156e-05, 5.976123e-05, 5.976139e-05, 5.976108e-05, 
    5.976094e-05, 5.976082e-05, 5.976067e-05, 5.976193e-05, 5.976197e-05, 
    5.976189e-05, 5.976178e-05, 5.976168e-05, 5.976155e-05, 5.976154e-05, 
    5.976151e-05, 5.976145e-05, 5.976139e-05, 5.97615e-05, 5.976138e-05, 
    5.976185e-05, 5.97616e-05, 5.976198e-05, 5.976187e-05, 5.976179e-05, 
    5.976182e-05, 5.976164e-05, 5.97616e-05, 5.976142e-05, 5.976151e-05, 
    5.976098e-05, 5.976121e-05, 5.976055e-05, 5.976074e-05, 5.976198e-05, 
    5.976193e-05, 5.976172e-05, 5.976182e-05, 5.976154e-05, 5.976147e-05, 
    5.976142e-05, 5.976135e-05, 5.976134e-05, 5.97613e-05, 5.976137e-05, 
    5.97613e-05, 5.976155e-05, 5.976144e-05, 5.976174e-05, 5.976167e-05, 
    5.97617e-05, 5.976174e-05, 5.976163e-05, 5.97615e-05, 5.97615e-05, 
    5.976146e-05, 5.976135e-05, 5.976154e-05, 5.976095e-05, 5.976131e-05, 
    5.976186e-05, 5.976175e-05, 5.976173e-05, 5.976178e-05, 5.976148e-05, 
    5.976159e-05, 5.97613e-05, 5.976138e-05, 5.976125e-05, 5.976131e-05, 
    5.976132e-05, 5.97614e-05, 5.976145e-05, 5.976158e-05, 5.976169e-05, 
    5.976177e-05, 5.976175e-05, 5.976166e-05, 5.976149e-05, 5.976134e-05, 
    5.976137e-05, 5.976126e-05, 5.976156e-05, 5.976143e-05, 5.976148e-05, 
    5.976135e-05, 5.976163e-05, 5.97614e-05, 5.97617e-05, 5.976167e-05, 
    5.976159e-05, 5.976142e-05, 5.976139e-05, 5.976135e-05, 5.976137e-05, 
    5.976149e-05, 5.976151e-05, 5.976159e-05, 5.976161e-05, 5.976167e-05, 
    5.976173e-05, 5.976168e-05, 5.976163e-05, 5.976149e-05, 5.976136e-05, 
    5.976122e-05, 5.976119e-05, 5.976103e-05, 5.976116e-05, 5.976094e-05, 
    5.976113e-05, 5.976081e-05, 5.976138e-05, 5.976113e-05, 5.976158e-05, 
    5.976154e-05, 5.976145e-05, 5.976125e-05, 5.976135e-05, 5.976123e-05, 
    5.976151e-05, 5.976166e-05, 5.976169e-05, 5.976177e-05, 5.976169e-05, 
    5.97617e-05, 5.976163e-05, 5.976165e-05, 5.976149e-05, 5.976157e-05, 
    5.976132e-05, 5.976123e-05, 5.976097e-05, 5.976081e-05, 5.976065e-05, 
    5.976058e-05, 5.976055e-05, 5.976054e-05 ;

 TOTLITN =
  1.375937e-06, 1.375933e-06, 1.375933e-06, 1.37593e-06, 1.375932e-06, 
    1.37593e-06, 1.375936e-06, 1.375932e-06, 1.375935e-06, 1.375936e-06, 
    1.375923e-06, 1.37593e-06, 1.375917e-06, 1.375921e-06, 1.375911e-06, 
    1.375917e-06, 1.375909e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375902e-06, 1.375906e-06, 1.375898e-06, 1.375903e-06, 1.375902e-06, 
    1.375906e-06, 1.375928e-06, 1.375924e-06, 1.375929e-06, 1.375928e-06, 
    1.375928e-06, 1.375932e-06, 1.375933e-06, 1.375937e-06, 1.375936e-06, 
    1.375934e-06, 1.375928e-06, 1.37593e-06, 1.375925e-06, 1.375925e-06, 
    1.375919e-06, 1.375922e-06, 1.375913e-06, 1.375915e-06, 1.375907e-06, 
    1.375909e-06, 1.375908e-06, 1.375908e-06, 1.375908e-06, 1.37591e-06, 
    1.375909e-06, 1.375912e-06, 1.375921e-06, 1.375919e-06, 1.375927e-06, 
    1.375932e-06, 1.375936e-06, 1.375938e-06, 1.375938e-06, 1.375937e-06, 
    1.375934e-06, 1.375931e-06, 1.375928e-06, 1.375927e-06, 1.375925e-06, 
    1.37592e-06, 1.375918e-06, 1.375912e-06, 1.375913e-06, 1.375911e-06, 
    1.37591e-06, 1.375907e-06, 1.375907e-06, 1.375906e-06, 1.375911e-06, 
    1.375908e-06, 1.375914e-06, 1.375912e-06, 1.375925e-06, 1.375929e-06, 
    1.375931e-06, 1.375933e-06, 1.375938e-06, 1.375935e-06, 1.375936e-06, 
    1.375933e-06, 1.375931e-06, 1.375932e-06, 1.375927e-06, 1.375929e-06, 
    1.375917e-06, 1.375922e-06, 1.37591e-06, 1.375913e-06, 1.375909e-06, 
    1.375911e-06, 1.375908e-06, 1.375911e-06, 1.375906e-06, 1.375905e-06, 
    1.375905e-06, 1.375902e-06, 1.375911e-06, 1.375908e-06, 1.375932e-06, 
    1.375932e-06, 1.375931e-06, 1.375934e-06, 1.375934e-06, 1.375937e-06, 
    1.375935e-06, 1.375934e-06, 1.375931e-06, 1.37593e-06, 1.375928e-06, 
    1.375925e-06, 1.375921e-06, 1.375916e-06, 1.375913e-06, 1.37591e-06, 
    1.375912e-06, 1.37591e-06, 1.375912e-06, 1.375912e-06, 1.375905e-06, 
    1.375909e-06, 1.375903e-06, 1.375903e-06, 1.375906e-06, 1.375903e-06, 
    1.375932e-06, 1.375933e-06, 1.375936e-06, 1.375933e-06, 1.375937e-06, 
    1.375935e-06, 1.375934e-06, 1.375929e-06, 1.375927e-06, 1.375926e-06, 
    1.375924e-06, 1.375922e-06, 1.375917e-06, 1.375913e-06, 1.37591e-06, 
    1.37591e-06, 1.37591e-06, 1.375909e-06, 1.375911e-06, 1.375909e-06, 
    1.375908e-06, 1.375909e-06, 1.375903e-06, 1.375905e-06, 1.375903e-06, 
    1.375904e-06, 1.375932e-06, 1.375931e-06, 1.375932e-06, 1.37593e-06, 
    1.375931e-06, 1.375927e-06, 1.375926e-06, 1.375919e-06, 1.375922e-06, 
    1.375918e-06, 1.375921e-06, 1.375921e-06, 1.375918e-06, 1.375921e-06, 
    1.375913e-06, 1.375919e-06, 1.375909e-06, 1.375914e-06, 1.375908e-06, 
    1.37591e-06, 1.375908e-06, 1.375906e-06, 1.375904e-06, 1.375901e-06, 
    1.375902e-06, 1.375899e-06, 1.375929e-06, 1.375927e-06, 1.375927e-06, 
    1.375925e-06, 1.375924e-06, 1.375921e-06, 1.375916e-06, 1.375918e-06, 
    1.375915e-06, 1.375914e-06, 1.375919e-06, 1.375916e-06, 1.375926e-06, 
    1.375924e-06, 1.375925e-06, 1.375929e-06, 1.375917e-06, 1.375923e-06, 
    1.375913e-06, 1.375916e-06, 1.375907e-06, 1.375911e-06, 1.375902e-06, 
    1.375898e-06, 1.375895e-06, 1.375891e-06, 1.375926e-06, 1.375927e-06, 
    1.375925e-06, 1.375922e-06, 1.375919e-06, 1.375916e-06, 1.375915e-06, 
    1.375914e-06, 1.375913e-06, 1.375911e-06, 1.375914e-06, 1.375911e-06, 
    1.375924e-06, 1.375917e-06, 1.375928e-06, 1.375925e-06, 1.375922e-06, 
    1.375923e-06, 1.375918e-06, 1.375917e-06, 1.375912e-06, 1.375915e-06, 
    1.375899e-06, 1.375906e-06, 1.375887e-06, 1.375893e-06, 1.375928e-06, 
    1.375926e-06, 1.37592e-06, 1.375923e-06, 1.375915e-06, 1.375913e-06, 
    1.375912e-06, 1.37591e-06, 1.37591e-06, 1.375908e-06, 1.37591e-06, 
    1.375908e-06, 1.375916e-06, 1.375912e-06, 1.375921e-06, 1.375919e-06, 
    1.37592e-06, 1.375921e-06, 1.375918e-06, 1.375914e-06, 1.375914e-06, 
    1.375913e-06, 1.37591e-06, 1.375915e-06, 1.375898e-06, 1.375909e-06, 
    1.375924e-06, 1.375921e-06, 1.375921e-06, 1.375922e-06, 1.375913e-06, 
    1.375917e-06, 1.375908e-06, 1.375911e-06, 1.375907e-06, 1.375909e-06, 
    1.375909e-06, 1.375911e-06, 1.375913e-06, 1.375916e-06, 1.375919e-06, 
    1.375922e-06, 1.375921e-06, 1.375919e-06, 1.375914e-06, 1.37591e-06, 
    1.375911e-06, 1.375907e-06, 1.375916e-06, 1.375912e-06, 1.375914e-06, 
    1.37591e-06, 1.375918e-06, 1.375911e-06, 1.37592e-06, 1.375919e-06, 
    1.375917e-06, 1.375912e-06, 1.375911e-06, 1.37591e-06, 1.375911e-06, 
    1.375914e-06, 1.375914e-06, 1.375917e-06, 1.375917e-06, 1.375919e-06, 
    1.375921e-06, 1.375919e-06, 1.375918e-06, 1.375914e-06, 1.37591e-06, 
    1.375906e-06, 1.375905e-06, 1.375901e-06, 1.375905e-06, 1.375898e-06, 
    1.375904e-06, 1.375895e-06, 1.375911e-06, 1.375904e-06, 1.375916e-06, 
    1.375915e-06, 1.375913e-06, 1.375907e-06, 1.37591e-06, 1.375906e-06, 
    1.375914e-06, 1.375918e-06, 1.37592e-06, 1.375922e-06, 1.37592e-06, 
    1.37592e-06, 1.375918e-06, 1.375918e-06, 1.375914e-06, 1.375916e-06, 
    1.375909e-06, 1.375906e-06, 1.375899e-06, 1.375895e-06, 1.37589e-06, 
    1.375888e-06, 1.375887e-06, 1.375887e-06 ;

 TOTLITN_1m =
  1.375937e-06, 1.375933e-06, 1.375933e-06, 1.37593e-06, 1.375932e-06, 
    1.37593e-06, 1.375936e-06, 1.375932e-06, 1.375935e-06, 1.375936e-06, 
    1.375923e-06, 1.37593e-06, 1.375917e-06, 1.375921e-06, 1.375911e-06, 
    1.375917e-06, 1.375909e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375902e-06, 1.375906e-06, 1.375898e-06, 1.375903e-06, 1.375902e-06, 
    1.375906e-06, 1.375928e-06, 1.375924e-06, 1.375929e-06, 1.375928e-06, 
    1.375928e-06, 1.375932e-06, 1.375933e-06, 1.375937e-06, 1.375936e-06, 
    1.375934e-06, 1.375928e-06, 1.37593e-06, 1.375925e-06, 1.375925e-06, 
    1.375919e-06, 1.375922e-06, 1.375913e-06, 1.375915e-06, 1.375907e-06, 
    1.375909e-06, 1.375908e-06, 1.375908e-06, 1.375908e-06, 1.37591e-06, 
    1.375909e-06, 1.375912e-06, 1.375921e-06, 1.375919e-06, 1.375927e-06, 
    1.375932e-06, 1.375936e-06, 1.375938e-06, 1.375938e-06, 1.375937e-06, 
    1.375934e-06, 1.375931e-06, 1.375928e-06, 1.375927e-06, 1.375925e-06, 
    1.37592e-06, 1.375918e-06, 1.375912e-06, 1.375913e-06, 1.375911e-06, 
    1.37591e-06, 1.375907e-06, 1.375907e-06, 1.375906e-06, 1.375911e-06, 
    1.375908e-06, 1.375914e-06, 1.375912e-06, 1.375925e-06, 1.375929e-06, 
    1.375931e-06, 1.375933e-06, 1.375938e-06, 1.375935e-06, 1.375936e-06, 
    1.375933e-06, 1.375931e-06, 1.375932e-06, 1.375927e-06, 1.375929e-06, 
    1.375917e-06, 1.375922e-06, 1.37591e-06, 1.375913e-06, 1.375909e-06, 
    1.375911e-06, 1.375908e-06, 1.375911e-06, 1.375906e-06, 1.375905e-06, 
    1.375905e-06, 1.375902e-06, 1.375911e-06, 1.375908e-06, 1.375932e-06, 
    1.375932e-06, 1.375931e-06, 1.375934e-06, 1.375934e-06, 1.375937e-06, 
    1.375935e-06, 1.375934e-06, 1.375931e-06, 1.37593e-06, 1.375928e-06, 
    1.375925e-06, 1.375921e-06, 1.375916e-06, 1.375913e-06, 1.37591e-06, 
    1.375912e-06, 1.37591e-06, 1.375912e-06, 1.375912e-06, 1.375905e-06, 
    1.375909e-06, 1.375903e-06, 1.375903e-06, 1.375906e-06, 1.375903e-06, 
    1.375932e-06, 1.375933e-06, 1.375936e-06, 1.375933e-06, 1.375937e-06, 
    1.375935e-06, 1.375934e-06, 1.375929e-06, 1.375927e-06, 1.375926e-06, 
    1.375924e-06, 1.375922e-06, 1.375917e-06, 1.375913e-06, 1.37591e-06, 
    1.37591e-06, 1.37591e-06, 1.375909e-06, 1.375911e-06, 1.375909e-06, 
    1.375908e-06, 1.375909e-06, 1.375903e-06, 1.375905e-06, 1.375903e-06, 
    1.375904e-06, 1.375932e-06, 1.375931e-06, 1.375932e-06, 1.37593e-06, 
    1.375931e-06, 1.375927e-06, 1.375926e-06, 1.375919e-06, 1.375922e-06, 
    1.375918e-06, 1.375921e-06, 1.375921e-06, 1.375918e-06, 1.375921e-06, 
    1.375913e-06, 1.375919e-06, 1.375909e-06, 1.375914e-06, 1.375908e-06, 
    1.37591e-06, 1.375908e-06, 1.375906e-06, 1.375904e-06, 1.375901e-06, 
    1.375902e-06, 1.375899e-06, 1.375929e-06, 1.375927e-06, 1.375927e-06, 
    1.375925e-06, 1.375924e-06, 1.375921e-06, 1.375916e-06, 1.375918e-06, 
    1.375915e-06, 1.375914e-06, 1.375919e-06, 1.375916e-06, 1.375926e-06, 
    1.375924e-06, 1.375925e-06, 1.375929e-06, 1.375917e-06, 1.375923e-06, 
    1.375913e-06, 1.375916e-06, 1.375907e-06, 1.375911e-06, 1.375902e-06, 
    1.375898e-06, 1.375895e-06, 1.375891e-06, 1.375926e-06, 1.375927e-06, 
    1.375925e-06, 1.375922e-06, 1.375919e-06, 1.375916e-06, 1.375915e-06, 
    1.375914e-06, 1.375913e-06, 1.375911e-06, 1.375914e-06, 1.375911e-06, 
    1.375924e-06, 1.375917e-06, 1.375928e-06, 1.375925e-06, 1.375922e-06, 
    1.375923e-06, 1.375918e-06, 1.375917e-06, 1.375912e-06, 1.375915e-06, 
    1.375899e-06, 1.375906e-06, 1.375887e-06, 1.375893e-06, 1.375928e-06, 
    1.375926e-06, 1.37592e-06, 1.375923e-06, 1.375915e-06, 1.375913e-06, 
    1.375912e-06, 1.37591e-06, 1.37591e-06, 1.375908e-06, 1.37591e-06, 
    1.375908e-06, 1.375916e-06, 1.375912e-06, 1.375921e-06, 1.375919e-06, 
    1.37592e-06, 1.375921e-06, 1.375918e-06, 1.375914e-06, 1.375914e-06, 
    1.375913e-06, 1.37591e-06, 1.375915e-06, 1.375898e-06, 1.375909e-06, 
    1.375924e-06, 1.375921e-06, 1.375921e-06, 1.375922e-06, 1.375913e-06, 
    1.375917e-06, 1.375908e-06, 1.375911e-06, 1.375907e-06, 1.375909e-06, 
    1.375909e-06, 1.375911e-06, 1.375913e-06, 1.375916e-06, 1.375919e-06, 
    1.375922e-06, 1.375921e-06, 1.375919e-06, 1.375914e-06, 1.37591e-06, 
    1.375911e-06, 1.375907e-06, 1.375916e-06, 1.375912e-06, 1.375914e-06, 
    1.37591e-06, 1.375918e-06, 1.375911e-06, 1.37592e-06, 1.375919e-06, 
    1.375917e-06, 1.375912e-06, 1.375911e-06, 1.37591e-06, 1.375911e-06, 
    1.375914e-06, 1.375914e-06, 1.375917e-06, 1.375917e-06, 1.375919e-06, 
    1.375921e-06, 1.375919e-06, 1.375918e-06, 1.375914e-06, 1.37591e-06, 
    1.375906e-06, 1.375905e-06, 1.375901e-06, 1.375905e-06, 1.375898e-06, 
    1.375904e-06, 1.375895e-06, 1.375911e-06, 1.375904e-06, 1.375916e-06, 
    1.375915e-06, 1.375913e-06, 1.375907e-06, 1.37591e-06, 1.375906e-06, 
    1.375914e-06, 1.375918e-06, 1.37592e-06, 1.375922e-06, 1.37592e-06, 
    1.37592e-06, 1.375918e-06, 1.375918e-06, 1.375914e-06, 1.375916e-06, 
    1.375909e-06, 1.375906e-06, 1.375899e-06, 1.375895e-06, 1.37589e-06, 
    1.375888e-06, 1.375887e-06, 1.375887e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.3448, 17.34478, 17.34479, 17.34477, 17.34478, 17.34477, 17.34479, 
    17.34478, 17.34479, 17.3448, 17.34476, 17.34477, 17.34473, 17.34475, 
    17.34471, 17.34474, 17.34471, 17.34472, 17.3447, 17.3447, 17.34468, 
    17.3447, 17.34468, 17.34469, 17.34469, 17.3447, 17.34477, 17.34476, 
    17.34477, 17.34477, 17.34477, 17.34478, 17.34479, 17.3448, 17.3448, 
    17.34479, 17.34477, 17.34477, 17.34476, 17.34476, 17.34474, 17.34475, 
    17.34472, 17.34473, 17.3447, 17.34471, 17.3447, 17.34471, 17.3447, 
    17.34471, 17.34471, 17.34472, 17.34475, 17.34474, 17.34477, 17.34478, 
    17.34479, 17.3448, 17.3448, 17.3448, 17.34479, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34472, 17.34472, 17.34472, 
    17.34471, 17.3447, 17.3447, 17.3447, 17.34472, 17.34471, 17.34472, 
    17.34472, 17.34476, 17.34477, 17.34478, 17.34479, 17.3448, 17.34479, 
    17.34479, 17.34478, 17.34478, 17.34478, 17.34476, 17.34477, 17.34474, 
    17.34475, 17.34471, 17.34472, 17.34471, 17.34472, 17.34471, 17.34471, 
    17.3447, 17.34469, 17.3447, 17.34469, 17.34472, 17.3447, 17.34478, 
    17.34478, 17.34478, 17.34479, 17.34479, 17.3448, 17.34479, 17.34479, 
    17.34478, 17.34477, 17.34477, 17.34476, 17.34475, 17.34473, 17.34472, 
    17.34471, 17.34472, 17.34471, 17.34472, 17.34472, 17.3447, 17.34471, 
    17.34469, 17.34469, 17.3447, 17.34469, 17.34478, 17.34478, 17.34479, 
    17.34479, 17.3448, 17.34479, 17.34479, 17.34477, 17.34477, 17.34476, 
    17.34476, 17.34475, 17.34473, 17.34472, 17.34471, 17.34471, 17.34471, 
    17.34471, 17.34472, 17.34471, 17.34471, 17.34471, 17.34469, 17.3447, 
    17.34469, 17.34469, 17.34478, 17.34478, 17.34478, 17.34478, 17.34478, 
    17.34476, 17.34476, 17.34474, 17.34475, 17.34474, 17.34475, 17.34475, 
    17.34474, 17.34475, 17.34472, 17.34474, 17.34471, 17.34472, 17.34471, 
    17.34471, 17.34471, 17.3447, 17.34469, 17.34468, 17.34469, 17.34468, 
    17.34477, 17.34476, 17.34477, 17.34476, 17.34476, 17.34475, 17.34473, 
    17.34474, 17.34473, 17.34472, 17.34474, 17.34473, 17.34476, 17.34476, 
    17.34476, 17.34477, 17.34474, 17.34475, 17.34472, 17.34473, 17.3447, 
    17.34472, 17.34469, 17.34468, 17.34466, 17.34465, 17.34476, 17.34477, 
    17.34476, 17.34475, 17.34474, 17.34473, 17.34473, 17.34473, 17.34472, 
    17.34472, 17.34472, 17.34471, 17.34476, 17.34473, 17.34477, 17.34476, 
    17.34475, 17.34475, 17.34474, 17.34473, 17.34472, 17.34473, 17.34468, 
    17.3447, 17.34464, 17.34466, 17.34477, 17.34476, 17.34474, 17.34475, 
    17.34473, 17.34472, 17.34472, 17.34471, 17.34471, 17.34471, 17.34471, 
    17.34471, 17.34473, 17.34472, 17.34475, 17.34474, 17.34474, 17.34475, 
    17.34474, 17.34472, 17.34472, 17.34472, 17.34471, 17.34473, 17.34468, 
    17.34471, 17.34476, 17.34475, 17.34475, 17.34475, 17.34472, 17.34473, 
    17.34471, 17.34471, 17.3447, 17.34471, 17.34471, 17.34472, 17.34472, 
    17.34473, 17.34474, 17.34475, 17.34475, 17.34474, 17.34472, 17.34471, 
    17.34471, 17.3447, 17.34473, 17.34472, 17.34472, 17.34471, 17.34474, 
    17.34472, 17.34474, 17.34474, 17.34473, 17.34472, 17.34472, 17.34471, 
    17.34471, 17.34472, 17.34472, 17.34473, 17.34473, 17.34474, 17.34475, 
    17.34474, 17.34474, 17.34472, 17.34471, 17.3447, 17.3447, 17.34468, 
    17.34469, 17.34468, 17.34469, 17.34466, 17.34472, 17.34469, 17.34473, 
    17.34473, 17.34472, 17.3447, 17.34471, 17.3447, 17.34472, 17.34474, 
    17.34474, 17.34475, 17.34474, 17.34474, 17.34474, 17.34474, 17.34472, 
    17.34473, 17.34471, 17.3447, 17.34468, 17.34466, 17.34465, 17.34464, 
    17.34464, 17.34464 ;

 TOTSOMC_1m =
  17.3448, 17.34478, 17.34479, 17.34477, 17.34478, 17.34477, 17.34479, 
    17.34478, 17.34479, 17.3448, 17.34476, 17.34477, 17.34473, 17.34475, 
    17.34471, 17.34474, 17.34471, 17.34472, 17.3447, 17.3447, 17.34468, 
    17.3447, 17.34468, 17.34469, 17.34469, 17.3447, 17.34477, 17.34476, 
    17.34477, 17.34477, 17.34477, 17.34478, 17.34479, 17.3448, 17.3448, 
    17.34479, 17.34477, 17.34477, 17.34476, 17.34476, 17.34474, 17.34475, 
    17.34472, 17.34473, 17.3447, 17.34471, 17.3447, 17.34471, 17.3447, 
    17.34471, 17.34471, 17.34472, 17.34475, 17.34474, 17.34477, 17.34478, 
    17.34479, 17.3448, 17.3448, 17.3448, 17.34479, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34472, 17.34472, 17.34472, 
    17.34471, 17.3447, 17.3447, 17.3447, 17.34472, 17.34471, 17.34472, 
    17.34472, 17.34476, 17.34477, 17.34478, 17.34479, 17.3448, 17.34479, 
    17.34479, 17.34478, 17.34478, 17.34478, 17.34476, 17.34477, 17.34474, 
    17.34475, 17.34471, 17.34472, 17.34471, 17.34472, 17.34471, 17.34471, 
    17.3447, 17.34469, 17.3447, 17.34469, 17.34472, 17.3447, 17.34478, 
    17.34478, 17.34478, 17.34479, 17.34479, 17.3448, 17.34479, 17.34479, 
    17.34478, 17.34477, 17.34477, 17.34476, 17.34475, 17.34473, 17.34472, 
    17.34471, 17.34472, 17.34471, 17.34472, 17.34472, 17.3447, 17.34471, 
    17.34469, 17.34469, 17.3447, 17.34469, 17.34478, 17.34478, 17.34479, 
    17.34479, 17.3448, 17.34479, 17.34479, 17.34477, 17.34477, 17.34476, 
    17.34476, 17.34475, 17.34473, 17.34472, 17.34471, 17.34471, 17.34471, 
    17.34471, 17.34472, 17.34471, 17.34471, 17.34471, 17.34469, 17.3447, 
    17.34469, 17.34469, 17.34478, 17.34478, 17.34478, 17.34478, 17.34478, 
    17.34476, 17.34476, 17.34474, 17.34475, 17.34474, 17.34475, 17.34475, 
    17.34474, 17.34475, 17.34472, 17.34474, 17.34471, 17.34472, 17.34471, 
    17.34471, 17.34471, 17.3447, 17.34469, 17.34468, 17.34469, 17.34468, 
    17.34477, 17.34476, 17.34477, 17.34476, 17.34476, 17.34475, 17.34473, 
    17.34474, 17.34473, 17.34472, 17.34474, 17.34473, 17.34476, 17.34476, 
    17.34476, 17.34477, 17.34474, 17.34475, 17.34472, 17.34473, 17.3447, 
    17.34472, 17.34469, 17.34468, 17.34466, 17.34465, 17.34476, 17.34477, 
    17.34476, 17.34475, 17.34474, 17.34473, 17.34473, 17.34473, 17.34472, 
    17.34472, 17.34472, 17.34471, 17.34476, 17.34473, 17.34477, 17.34476, 
    17.34475, 17.34475, 17.34474, 17.34473, 17.34472, 17.34473, 17.34468, 
    17.3447, 17.34464, 17.34466, 17.34477, 17.34476, 17.34474, 17.34475, 
    17.34473, 17.34472, 17.34472, 17.34471, 17.34471, 17.34471, 17.34471, 
    17.34471, 17.34473, 17.34472, 17.34475, 17.34474, 17.34474, 17.34475, 
    17.34474, 17.34472, 17.34472, 17.34472, 17.34471, 17.34473, 17.34468, 
    17.34471, 17.34476, 17.34475, 17.34475, 17.34475, 17.34472, 17.34473, 
    17.34471, 17.34471, 17.3447, 17.34471, 17.34471, 17.34472, 17.34472, 
    17.34473, 17.34474, 17.34475, 17.34475, 17.34474, 17.34472, 17.34471, 
    17.34471, 17.3447, 17.34473, 17.34472, 17.34472, 17.34471, 17.34474, 
    17.34472, 17.34474, 17.34474, 17.34473, 17.34472, 17.34472, 17.34471, 
    17.34471, 17.34472, 17.34472, 17.34473, 17.34473, 17.34474, 17.34475, 
    17.34474, 17.34474, 17.34472, 17.34471, 17.3447, 17.3447, 17.34468, 
    17.34469, 17.34468, 17.34469, 17.34466, 17.34472, 17.34469, 17.34473, 
    17.34473, 17.34472, 17.3447, 17.34471, 17.3447, 17.34472, 17.34474, 
    17.34474, 17.34475, 17.34474, 17.34474, 17.34474, 17.34474, 17.34472, 
    17.34473, 17.34471, 17.3447, 17.34468, 17.34466, 17.34465, 17.34464, 
    17.34464, 17.34464 ;

 TOTSOMN =
  1.773785, 1.773783, 1.773783, 1.773782, 1.773782, 1.773781, 1.773784, 
    1.773783, 1.773784, 1.773784, 1.773779, 1.773782, 1.773776, 1.773777, 
    1.773773, 1.773776, 1.773772, 1.773773, 1.773771, 1.773772, 1.773769, 
    1.773771, 1.773767, 1.773769, 1.773769, 1.773771, 1.773781, 1.773779, 
    1.773781, 1.773781, 1.773781, 1.773782, 1.773783, 1.773785, 1.773784, 
    1.773783, 1.773781, 1.773782, 1.773779, 1.773779, 1.773777, 1.773778, 
    1.773774, 1.773775, 1.773772, 1.773772, 1.773772, 1.773772, 1.773772, 
    1.773773, 1.773772, 1.773773, 1.773778, 1.773777, 1.77378, 1.773783, 
    1.773784, 1.773785, 1.773785, 1.773785, 1.773783, 1.773782, 1.773781, 
    1.77378, 1.773779, 1.773777, 1.773776, 1.773774, 1.773774, 1.773773, 
    1.773772, 1.773771, 1.773772, 1.773771, 1.773773, 1.773772, 1.773774, 
    1.773774, 1.773779, 1.773781, 1.773782, 1.773783, 1.773785, 1.773784, 
    1.773784, 1.773783, 1.773782, 1.773782, 1.77378, 1.773781, 1.773776, 
    1.773778, 1.773773, 1.773774, 1.773772, 1.773773, 1.773772, 1.773773, 
    1.773771, 1.77377, 1.773771, 1.773769, 1.773773, 1.773772, 1.773782, 
    1.773782, 1.773782, 1.773783, 1.773783, 1.773785, 1.773784, 1.773783, 
    1.773782, 1.773781, 1.773781, 1.773779, 1.773778, 1.773775, 1.773774, 
    1.773773, 1.773773, 1.773773, 1.773773, 1.773774, 1.77377, 1.773772, 
    1.773769, 1.77377, 1.773771, 1.77377, 1.773782, 1.773783, 1.773784, 
    1.773783, 1.773785, 1.773784, 1.773783, 1.773781, 1.77378, 1.77378, 
    1.773779, 1.773778, 1.773776, 1.773774, 1.773772, 1.773773, 1.773773, 
    1.773772, 1.773773, 1.773772, 1.773772, 1.773772, 1.77377, 1.77377, 
    1.77377, 1.77377, 1.773783, 1.773782, 1.773782, 1.773782, 1.773782, 
    1.77378, 1.77378, 1.773777, 1.773778, 1.773776, 1.773778, 1.773777, 
    1.773776, 1.773778, 1.773774, 1.773777, 1.773772, 1.773775, 1.773772, 
    1.773772, 1.773772, 1.773771, 1.77377, 1.773769, 1.773769, 1.773768, 
    1.773781, 1.77378, 1.77378, 1.77378, 1.773779, 1.773777, 1.773775, 
    1.773776, 1.773775, 1.773774, 1.773777, 1.773775, 1.77378, 1.773779, 
    1.773779, 1.773781, 1.773776, 1.773779, 1.773774, 1.773775, 1.773771, 
    1.773773, 1.773769, 1.773767, 1.773766, 1.773764, 1.77378, 1.77378, 
    1.773779, 1.773778, 1.773777, 1.773775, 1.773775, 1.773775, 1.773774, 
    1.773773, 1.773775, 1.773773, 1.773779, 1.773776, 1.773781, 1.773779, 
    1.773778, 1.773779, 1.773776, 1.773776, 1.773774, 1.773775, 1.773768, 
    1.773771, 1.773763, 1.773765, 1.773781, 1.77378, 1.773777, 1.773778, 
    1.773775, 1.773774, 1.773773, 1.773773, 1.773772, 1.773772, 1.773773, 
    1.773772, 1.773775, 1.773774, 1.773778, 1.773777, 1.773777, 1.773777, 
    1.773776, 1.773775, 1.773775, 1.773774, 1.773773, 1.773775, 1.773767, 
    1.773772, 1.773779, 1.773778, 1.773777, 1.773778, 1.773774, 1.773776, 
    1.773772, 1.773773, 1.773771, 1.773772, 1.773772, 1.773773, 1.773774, 
    1.773776, 1.773777, 1.773778, 1.773778, 1.773777, 1.773774, 1.773772, 
    1.773773, 1.773771, 1.773775, 1.773774, 1.773774, 1.773773, 1.773776, 
    1.773773, 1.773777, 1.773777, 1.773776, 1.773774, 1.773773, 1.773773, 
    1.773773, 1.773774, 1.773775, 1.773776, 1.773776, 1.773777, 1.773777, 
    1.773777, 1.773776, 1.773774, 1.773773, 1.773771, 1.773771, 1.773769, 
    1.77377, 1.773767, 1.77377, 1.773766, 1.773773, 1.77377, 1.773776, 
    1.773775, 1.773774, 1.773771, 1.773773, 1.773771, 1.773775, 1.773776, 
    1.773777, 1.773778, 1.773777, 1.773777, 1.773776, 1.773776, 1.773774, 
    1.773775, 1.773772, 1.773771, 1.773768, 1.773766, 1.773764, 1.773763, 
    1.773763, 1.773762 ;

 TOTSOMN_1m =
  1.773785, 1.773783, 1.773783, 1.773782, 1.773782, 1.773781, 1.773784, 
    1.773783, 1.773784, 1.773784, 1.773779, 1.773782, 1.773776, 1.773777, 
    1.773773, 1.773776, 1.773772, 1.773773, 1.773771, 1.773772, 1.773769, 
    1.773771, 1.773767, 1.773769, 1.773769, 1.773771, 1.773781, 1.773779, 
    1.773781, 1.773781, 1.773781, 1.773782, 1.773783, 1.773785, 1.773784, 
    1.773783, 1.773781, 1.773782, 1.773779, 1.773779, 1.773777, 1.773778, 
    1.773774, 1.773775, 1.773772, 1.773772, 1.773772, 1.773772, 1.773772, 
    1.773773, 1.773772, 1.773773, 1.773778, 1.773777, 1.77378, 1.773783, 
    1.773784, 1.773785, 1.773785, 1.773785, 1.773783, 1.773782, 1.773781, 
    1.77378, 1.773779, 1.773777, 1.773776, 1.773774, 1.773774, 1.773773, 
    1.773772, 1.773771, 1.773772, 1.773771, 1.773773, 1.773772, 1.773774, 
    1.773774, 1.773779, 1.773781, 1.773782, 1.773783, 1.773785, 1.773784, 
    1.773784, 1.773783, 1.773782, 1.773782, 1.77378, 1.773781, 1.773776, 
    1.773778, 1.773773, 1.773774, 1.773772, 1.773773, 1.773772, 1.773773, 
    1.773771, 1.77377, 1.773771, 1.773769, 1.773773, 1.773772, 1.773782, 
    1.773782, 1.773782, 1.773783, 1.773783, 1.773785, 1.773784, 1.773783, 
    1.773782, 1.773781, 1.773781, 1.773779, 1.773778, 1.773775, 1.773774, 
    1.773773, 1.773773, 1.773773, 1.773773, 1.773774, 1.77377, 1.773772, 
    1.773769, 1.77377, 1.773771, 1.77377, 1.773782, 1.773783, 1.773784, 
    1.773783, 1.773785, 1.773784, 1.773783, 1.773781, 1.77378, 1.77378, 
    1.773779, 1.773778, 1.773776, 1.773774, 1.773772, 1.773773, 1.773773, 
    1.773772, 1.773773, 1.773772, 1.773772, 1.773772, 1.77377, 1.77377, 
    1.77377, 1.77377, 1.773783, 1.773782, 1.773782, 1.773782, 1.773782, 
    1.77378, 1.77378, 1.773777, 1.773778, 1.773776, 1.773778, 1.773777, 
    1.773776, 1.773778, 1.773774, 1.773777, 1.773772, 1.773775, 1.773772, 
    1.773772, 1.773772, 1.773771, 1.77377, 1.773769, 1.773769, 1.773768, 
    1.773781, 1.77378, 1.77378, 1.77378, 1.773779, 1.773777, 1.773775, 
    1.773776, 1.773775, 1.773774, 1.773777, 1.773775, 1.77378, 1.773779, 
    1.773779, 1.773781, 1.773776, 1.773779, 1.773774, 1.773775, 1.773771, 
    1.773773, 1.773769, 1.773767, 1.773766, 1.773764, 1.77378, 1.77378, 
    1.773779, 1.773778, 1.773777, 1.773775, 1.773775, 1.773775, 1.773774, 
    1.773773, 1.773775, 1.773773, 1.773779, 1.773776, 1.773781, 1.773779, 
    1.773778, 1.773779, 1.773776, 1.773776, 1.773774, 1.773775, 1.773768, 
    1.773771, 1.773763, 1.773765, 1.773781, 1.77378, 1.773777, 1.773778, 
    1.773775, 1.773774, 1.773773, 1.773773, 1.773772, 1.773772, 1.773773, 
    1.773772, 1.773775, 1.773774, 1.773778, 1.773777, 1.773777, 1.773777, 
    1.773776, 1.773775, 1.773775, 1.773774, 1.773773, 1.773775, 1.773767, 
    1.773772, 1.773779, 1.773778, 1.773777, 1.773778, 1.773774, 1.773776, 
    1.773772, 1.773773, 1.773771, 1.773772, 1.773772, 1.773773, 1.773774, 
    1.773776, 1.773777, 1.773778, 1.773778, 1.773777, 1.773774, 1.773772, 
    1.773773, 1.773771, 1.773775, 1.773774, 1.773774, 1.773773, 1.773776, 
    1.773773, 1.773777, 1.773777, 1.773776, 1.773774, 1.773773, 1.773773, 
    1.773773, 1.773774, 1.773775, 1.773776, 1.773776, 1.773777, 1.773777, 
    1.773777, 1.773776, 1.773774, 1.773773, 1.773771, 1.773771, 1.773769, 
    1.77377, 1.773767, 1.77377, 1.773766, 1.773773, 1.77377, 1.773776, 
    1.773775, 1.773774, 1.773771, 1.773773, 1.773771, 1.773775, 1.773776, 
    1.773777, 1.773778, 1.773777, 1.773777, 1.773776, 1.773776, 1.773774, 
    1.773775, 1.773772, 1.773771, 1.773768, 1.773766, 1.773764, 1.773763, 
    1.773763, 1.773762 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  249.9807, 249.9809, 249.9809, 249.9811, 249.981, 249.9811, 249.9807, 
    249.9809, 249.9808, 249.9807, 249.9815, 249.9811, 249.9819, 249.9817, 
    249.9823, 249.9819, 249.9824, 249.9823, 249.9826, 249.9825, 249.9829, 
    249.9827, 249.9831, 249.9828, 249.9829, 249.9826, 249.9812, 249.9814, 
    249.9812, 249.9812, 249.9812, 249.981, 249.9809, 249.9807, 249.9807, 
    249.9809, 249.9812, 249.9811, 249.9814, 249.9814, 249.9818, 249.9816, 
    249.9822, 249.982, 249.9825, 249.9824, 249.9825, 249.9825, 249.9825, 
    249.9823, 249.9824, 249.9823, 249.9816, 249.9818, 249.9813, 249.9809, 
    249.9807, 249.9806, 249.9806, 249.9806, 249.9809, 249.981, 249.9812, 
    249.9813, 249.9814, 249.9817, 249.9819, 249.9822, 249.9822, 249.9823, 
    249.9824, 249.9826, 249.9825, 249.9826, 249.9823, 249.9825, 249.9821, 
    249.9822, 249.9814, 249.9811, 249.981, 249.9809, 249.9806, 249.9808, 
    249.9807, 249.9809, 249.981, 249.981, 249.9813, 249.9812, 249.9819, 
    249.9816, 249.9824, 249.9822, 249.9824, 249.9823, 249.9825, 249.9823, 
    249.9826, 249.9827, 249.9827, 249.9828, 249.9823, 249.9825, 249.981, 
    249.981, 249.981, 249.9808, 249.9808, 249.9807, 249.9808, 249.9809, 
    249.981, 249.9811, 249.9812, 249.9814, 249.9816, 249.982, 249.9822, 
    249.9823, 249.9823, 249.9823, 249.9822, 249.9822, 249.9827, 249.9824, 
    249.9828, 249.9828, 249.9826, 249.9828, 249.981, 249.9809, 249.9807, 
    249.9809, 249.9806, 249.9808, 249.9809, 249.9812, 249.9812, 249.9813, 
    249.9814, 249.9816, 249.9819, 249.9822, 249.9824, 249.9824, 249.9824, 
    249.9824, 249.9823, 249.9825, 249.9825, 249.9824, 249.9828, 249.9827, 
    249.9828, 249.9827, 249.9809, 249.981, 249.981, 249.9811, 249.981, 
    249.9813, 249.9814, 249.9818, 249.9816, 249.9819, 249.9816, 249.9817, 
    249.9819, 249.9816, 249.9821, 249.9818, 249.9824, 249.9821, 249.9825, 
    249.9824, 249.9825, 249.9826, 249.9827, 249.9829, 249.9829, 249.9831, 
    249.9812, 249.9813, 249.9813, 249.9814, 249.9815, 249.9817, 249.982, 
    249.9819, 249.9821, 249.9821, 249.9818, 249.982, 249.9814, 249.9814, 
    249.9814, 249.9812, 249.9819, 249.9815, 249.9822, 249.982, 249.9826, 
    249.9823, 249.9829, 249.9831, 249.9833, 249.9836, 249.9813, 249.9813, 
    249.9814, 249.9816, 249.9818, 249.982, 249.982, 249.9821, 249.9822, 
    249.9823, 249.9821, 249.9823, 249.9815, 249.9819, 249.9812, 249.9814, 
    249.9816, 249.9815, 249.9818, 249.9819, 249.9822, 249.9821, 249.983, 
    249.9826, 249.9838, 249.9835, 249.9812, 249.9813, 249.9817, 249.9815, 
    249.982, 249.9821, 249.9823, 249.9824, 249.9824, 249.9825, 249.9823, 
    249.9825, 249.982, 249.9822, 249.9817, 249.9818, 249.9817, 249.9817, 
    249.9819, 249.9821, 249.9821, 249.9822, 249.9824, 249.982, 249.9831, 
    249.9824, 249.9815, 249.9816, 249.9817, 249.9816, 249.9821, 249.9819, 
    249.9825, 249.9823, 249.9826, 249.9824, 249.9824, 249.9823, 249.9822, 
    249.9819, 249.9818, 249.9816, 249.9817, 249.9818, 249.9821, 249.9824, 
    249.9823, 249.9825, 249.982, 249.9822, 249.9821, 249.9824, 249.9819, 
    249.9823, 249.9818, 249.9818, 249.9819, 249.9822, 249.9823, 249.9824, 
    249.9823, 249.9821, 249.9821, 249.9819, 249.9819, 249.9818, 249.9817, 
    249.9818, 249.9819, 249.9821, 249.9823, 249.9826, 249.9827, 249.9829, 
    249.9827, 249.9831, 249.9827, 249.9833, 249.9823, 249.9827, 249.9819, 
    249.982, 249.9822, 249.9825, 249.9824, 249.9826, 249.9821, 249.9818, 
    249.9818, 249.9816, 249.9818, 249.9818, 249.9819, 249.9818, 249.9821, 
    249.982, 249.9824, 249.9826, 249.983, 249.9833, 249.9836, 249.9838, 
    249.9838, 249.9838 ;

 TREFMNAV_R =
  249.9807, 249.9809, 249.9809, 249.9811, 249.981, 249.9811, 249.9807, 
    249.9809, 249.9808, 249.9807, 249.9815, 249.9811, 249.9819, 249.9817, 
    249.9823, 249.9819, 249.9824, 249.9823, 249.9826, 249.9825, 249.9829, 
    249.9827, 249.9831, 249.9828, 249.9829, 249.9826, 249.9812, 249.9814, 
    249.9812, 249.9812, 249.9812, 249.981, 249.9809, 249.9807, 249.9807, 
    249.9809, 249.9812, 249.9811, 249.9814, 249.9814, 249.9818, 249.9816, 
    249.9822, 249.982, 249.9825, 249.9824, 249.9825, 249.9825, 249.9825, 
    249.9823, 249.9824, 249.9823, 249.9816, 249.9818, 249.9813, 249.9809, 
    249.9807, 249.9806, 249.9806, 249.9806, 249.9809, 249.981, 249.9812, 
    249.9813, 249.9814, 249.9817, 249.9819, 249.9822, 249.9822, 249.9823, 
    249.9824, 249.9826, 249.9825, 249.9826, 249.9823, 249.9825, 249.9821, 
    249.9822, 249.9814, 249.9811, 249.981, 249.9809, 249.9806, 249.9808, 
    249.9807, 249.9809, 249.981, 249.981, 249.9813, 249.9812, 249.9819, 
    249.9816, 249.9824, 249.9822, 249.9824, 249.9823, 249.9825, 249.9823, 
    249.9826, 249.9827, 249.9827, 249.9828, 249.9823, 249.9825, 249.981, 
    249.981, 249.981, 249.9808, 249.9808, 249.9807, 249.9808, 249.9809, 
    249.981, 249.9811, 249.9812, 249.9814, 249.9816, 249.982, 249.9822, 
    249.9823, 249.9823, 249.9823, 249.9822, 249.9822, 249.9827, 249.9824, 
    249.9828, 249.9828, 249.9826, 249.9828, 249.981, 249.9809, 249.9807, 
    249.9809, 249.9806, 249.9808, 249.9809, 249.9812, 249.9812, 249.9813, 
    249.9814, 249.9816, 249.9819, 249.9822, 249.9824, 249.9824, 249.9824, 
    249.9824, 249.9823, 249.9825, 249.9825, 249.9824, 249.9828, 249.9827, 
    249.9828, 249.9827, 249.9809, 249.981, 249.981, 249.9811, 249.981, 
    249.9813, 249.9814, 249.9818, 249.9816, 249.9819, 249.9816, 249.9817, 
    249.9819, 249.9816, 249.9821, 249.9818, 249.9824, 249.9821, 249.9825, 
    249.9824, 249.9825, 249.9826, 249.9827, 249.9829, 249.9829, 249.9831, 
    249.9812, 249.9813, 249.9813, 249.9814, 249.9815, 249.9817, 249.982, 
    249.9819, 249.9821, 249.9821, 249.9818, 249.982, 249.9814, 249.9814, 
    249.9814, 249.9812, 249.9819, 249.9815, 249.9822, 249.982, 249.9826, 
    249.9823, 249.9829, 249.9831, 249.9833, 249.9836, 249.9813, 249.9813, 
    249.9814, 249.9816, 249.9818, 249.982, 249.982, 249.9821, 249.9822, 
    249.9823, 249.9821, 249.9823, 249.9815, 249.9819, 249.9812, 249.9814, 
    249.9816, 249.9815, 249.9818, 249.9819, 249.9822, 249.9821, 249.983, 
    249.9826, 249.9838, 249.9835, 249.9812, 249.9813, 249.9817, 249.9815, 
    249.982, 249.9821, 249.9823, 249.9824, 249.9824, 249.9825, 249.9823, 
    249.9825, 249.982, 249.9822, 249.9817, 249.9818, 249.9817, 249.9817, 
    249.9819, 249.9821, 249.9821, 249.9822, 249.9824, 249.982, 249.9831, 
    249.9824, 249.9815, 249.9816, 249.9817, 249.9816, 249.9821, 249.9819, 
    249.9825, 249.9823, 249.9826, 249.9824, 249.9824, 249.9823, 249.9822, 
    249.9819, 249.9818, 249.9816, 249.9817, 249.9818, 249.9821, 249.9824, 
    249.9823, 249.9825, 249.982, 249.9822, 249.9821, 249.9824, 249.9819, 
    249.9823, 249.9818, 249.9818, 249.9819, 249.9822, 249.9823, 249.9824, 
    249.9823, 249.9821, 249.9821, 249.9819, 249.9819, 249.9818, 249.9817, 
    249.9818, 249.9819, 249.9821, 249.9823, 249.9826, 249.9827, 249.9829, 
    249.9827, 249.9831, 249.9827, 249.9833, 249.9823, 249.9827, 249.9819, 
    249.982, 249.9822, 249.9825, 249.9824, 249.9826, 249.9821, 249.9818, 
    249.9818, 249.9816, 249.9818, 249.9818, 249.9819, 249.9818, 249.9821, 
    249.982, 249.9824, 249.9826, 249.983, 249.9833, 249.9836, 249.9838, 
    249.9838, 249.9838 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  258.6014, 258.6018, 258.6017, 258.602, 258.6019, 258.6021, 258.6015, 
    258.6018, 258.6016, 258.6014, 258.6026, 258.6021, 258.6032, 258.6029, 
    258.6038, 258.6032, 258.6039, 258.6038, 258.6042, 258.6041, 258.6048, 
    258.6043, 258.6051, 258.6047, 258.6048, 258.6043, 258.6022, 258.6025, 
    258.6021, 258.6022, 258.6022, 258.6019, 258.6017, 258.6014, 258.6014, 
    258.6017, 258.6022, 258.6021, 258.6025, 258.6025, 258.603, 258.6028, 
    258.6037, 258.6034, 258.6041, 258.6039, 258.6041, 258.6041, 258.6041, 
    258.6039, 258.604, 258.6037, 258.6028, 258.6031, 258.6023, 258.6018, 
    258.6015, 258.6013, 258.6013, 258.6014, 258.6017, 258.602, 258.6022, 
    258.6024, 258.6025, 258.6029, 258.6032, 258.6037, 258.6036, 258.6038, 
    258.6039, 258.6042, 258.6042, 258.6043, 258.6038, 258.6041, 258.6036, 
    258.6037, 258.6025, 258.6021, 258.6019, 258.6017, 258.6013, 258.6016, 
    258.6015, 258.6018, 258.6019, 258.6018, 258.6024, 258.6021, 258.6032, 
    258.6028, 258.6039, 258.6036, 258.604, 258.6038, 258.6041, 258.6039, 
    258.6043, 258.6046, 258.6043, 258.6047, 258.6038, 258.6041, 258.6018, 
    258.6019, 258.6019, 258.6017, 258.6016, 258.6014, 258.6016, 258.6017, 
    258.6019, 258.6021, 258.6022, 258.6025, 258.6028, 258.6033, 258.6036, 
    258.6039, 258.6037, 258.6039, 258.6037, 258.6037, 258.6045, 258.604, 
    258.6047, 258.6047, 258.6043, 258.6047, 258.6019, 258.6018, 258.6015, 
    258.6017, 258.6013, 258.6016, 258.6017, 258.6021, 258.6023, 258.6024, 
    258.6025, 258.6028, 258.6032, 258.6036, 258.6039, 258.6039, 258.6039, 
    258.604, 258.6038, 258.604, 258.6041, 258.604, 258.6047, 258.6045, 
    258.6047, 258.6046, 258.6018, 258.602, 258.6019, 258.602, 258.6019, 
    258.6023, 258.6024, 258.603, 258.6028, 258.6031, 258.6028, 258.6029, 
    258.6032, 258.6028, 258.6036, 258.6031, 258.604, 258.6035, 258.604, 
    258.6039, 258.6041, 258.6042, 258.6046, 258.6049, 258.6048, 258.605, 
    258.6021, 258.6023, 258.6023, 258.6025, 258.6026, 258.6029, 258.6033, 
    258.6031, 258.6035, 258.6035, 258.6031, 258.6034, 258.6024, 258.6026, 
    258.6025, 258.6021, 258.6032, 258.6027, 258.6037, 258.6034, 258.6042, 
    258.6038, 258.6048, 258.6051, 258.6054, 258.6057, 258.6024, 258.6023, 
    258.6025, 258.6028, 258.603, 258.6034, 258.6034, 258.6035, 258.6037, 
    258.6038, 258.6035, 258.6038, 258.6026, 258.6032, 258.6022, 258.6025, 
    258.6028, 258.6027, 258.6031, 258.6033, 258.6037, 258.6035, 258.605, 
    258.6043, 258.606, 258.6056, 258.6022, 258.6024, 258.6029, 258.6027, 
    258.6034, 258.6036, 258.6037, 258.6039, 258.6039, 258.6041, 258.6039, 
    258.604, 258.6034, 258.6037, 258.6029, 258.6031, 258.603, 258.6029, 
    258.6032, 258.6035, 258.6035, 258.6036, 258.6039, 258.6034, 258.605, 
    258.604, 258.6026, 258.6028, 258.6029, 258.6028, 258.6036, 258.6033, 
    258.604, 258.6039, 258.6042, 258.604, 258.604, 258.6038, 258.6036, 
    258.6033, 258.603, 258.6028, 258.6028, 258.6031, 258.6035, 258.6039, 
    258.6039, 258.6042, 258.6034, 258.6037, 258.6035, 258.6039, 258.6031, 
    258.6038, 258.603, 258.6031, 258.6033, 258.6037, 258.6038, 258.6039, 
    258.6039, 258.6035, 258.6035, 258.6033, 258.6032, 258.6031, 258.6029, 
    258.603, 258.6032, 258.6035, 258.6039, 258.6042, 258.6043, 258.6049, 
    258.6046, 258.605, 258.6046, 258.6054, 258.6038, 258.6046, 258.6033, 
    258.6034, 258.6036, 258.6042, 258.6039, 258.6042, 258.6035, 258.6031, 
    258.603, 258.6028, 258.603, 258.603, 258.6032, 258.6031, 258.6035, 
    258.6033, 258.604, 258.6042, 258.605, 258.6054, 258.6058, 258.606, 
    258.606, 258.606 ;

 TREFMXAV_R =
  258.6014, 258.6018, 258.6017, 258.602, 258.6019, 258.6021, 258.6015, 
    258.6018, 258.6016, 258.6014, 258.6026, 258.6021, 258.6032, 258.6029, 
    258.6038, 258.6032, 258.6039, 258.6038, 258.6042, 258.6041, 258.6048, 
    258.6043, 258.6051, 258.6047, 258.6048, 258.6043, 258.6022, 258.6025, 
    258.6021, 258.6022, 258.6022, 258.6019, 258.6017, 258.6014, 258.6014, 
    258.6017, 258.6022, 258.6021, 258.6025, 258.6025, 258.603, 258.6028, 
    258.6037, 258.6034, 258.6041, 258.6039, 258.6041, 258.6041, 258.6041, 
    258.6039, 258.604, 258.6037, 258.6028, 258.6031, 258.6023, 258.6018, 
    258.6015, 258.6013, 258.6013, 258.6014, 258.6017, 258.602, 258.6022, 
    258.6024, 258.6025, 258.6029, 258.6032, 258.6037, 258.6036, 258.6038, 
    258.6039, 258.6042, 258.6042, 258.6043, 258.6038, 258.6041, 258.6036, 
    258.6037, 258.6025, 258.6021, 258.6019, 258.6017, 258.6013, 258.6016, 
    258.6015, 258.6018, 258.6019, 258.6018, 258.6024, 258.6021, 258.6032, 
    258.6028, 258.6039, 258.6036, 258.604, 258.6038, 258.6041, 258.6039, 
    258.6043, 258.6046, 258.6043, 258.6047, 258.6038, 258.6041, 258.6018, 
    258.6019, 258.6019, 258.6017, 258.6016, 258.6014, 258.6016, 258.6017, 
    258.6019, 258.6021, 258.6022, 258.6025, 258.6028, 258.6033, 258.6036, 
    258.6039, 258.6037, 258.6039, 258.6037, 258.6037, 258.6045, 258.604, 
    258.6047, 258.6047, 258.6043, 258.6047, 258.6019, 258.6018, 258.6015, 
    258.6017, 258.6013, 258.6016, 258.6017, 258.6021, 258.6023, 258.6024, 
    258.6025, 258.6028, 258.6032, 258.6036, 258.6039, 258.6039, 258.6039, 
    258.604, 258.6038, 258.604, 258.6041, 258.604, 258.6047, 258.6045, 
    258.6047, 258.6046, 258.6018, 258.602, 258.6019, 258.602, 258.6019, 
    258.6023, 258.6024, 258.603, 258.6028, 258.6031, 258.6028, 258.6029, 
    258.6032, 258.6028, 258.6036, 258.6031, 258.604, 258.6035, 258.604, 
    258.6039, 258.6041, 258.6042, 258.6046, 258.6049, 258.6048, 258.605, 
    258.6021, 258.6023, 258.6023, 258.6025, 258.6026, 258.6029, 258.6033, 
    258.6031, 258.6035, 258.6035, 258.6031, 258.6034, 258.6024, 258.6026, 
    258.6025, 258.6021, 258.6032, 258.6027, 258.6037, 258.6034, 258.6042, 
    258.6038, 258.6048, 258.6051, 258.6054, 258.6057, 258.6024, 258.6023, 
    258.6025, 258.6028, 258.603, 258.6034, 258.6034, 258.6035, 258.6037, 
    258.6038, 258.6035, 258.6038, 258.6026, 258.6032, 258.6022, 258.6025, 
    258.6028, 258.6027, 258.6031, 258.6033, 258.6037, 258.6035, 258.605, 
    258.6043, 258.606, 258.6056, 258.6022, 258.6024, 258.6029, 258.6027, 
    258.6034, 258.6036, 258.6037, 258.6039, 258.6039, 258.6041, 258.6039, 
    258.604, 258.6034, 258.6037, 258.6029, 258.6031, 258.603, 258.6029, 
    258.6032, 258.6035, 258.6035, 258.6036, 258.6039, 258.6034, 258.605, 
    258.604, 258.6026, 258.6028, 258.6029, 258.6028, 258.6036, 258.6033, 
    258.604, 258.6039, 258.6042, 258.604, 258.604, 258.6038, 258.6036, 
    258.6033, 258.603, 258.6028, 258.6028, 258.6031, 258.6035, 258.6039, 
    258.6039, 258.6042, 258.6034, 258.6037, 258.6035, 258.6039, 258.6031, 
    258.6038, 258.603, 258.6031, 258.6033, 258.6037, 258.6038, 258.6039, 
    258.6039, 258.6035, 258.6035, 258.6033, 258.6032, 258.6031, 258.6029, 
    258.603, 258.6032, 258.6035, 258.6039, 258.6042, 258.6043, 258.6049, 
    258.6046, 258.605, 258.6046, 258.6054, 258.6038, 258.6046, 258.6033, 
    258.6034, 258.6036, 258.6042, 258.6039, 258.6042, 258.6035, 258.6031, 
    258.603, 258.6028, 258.603, 258.603, 258.6032, 258.6031, 258.6035, 
    258.6033, 258.604, 258.6042, 258.605, 258.6054, 258.6058, 258.606, 
    258.606, 258.606 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  253.9724, 253.9726, 253.9725, 253.9727, 253.9726, 253.9727, 253.9724, 
    253.9726, 253.9725, 253.9724, 253.9729, 253.9727, 253.9732, 253.973, 
    253.9734, 253.9732, 253.9735, 253.9734, 253.9736, 253.9736, 253.9738, 
    253.9737, 253.974, 253.9738, 253.9738, 253.9737, 253.9727, 253.9729, 
    253.9727, 253.9727, 253.9727, 253.9726, 253.9725, 253.9724, 253.9724, 
    253.9725, 253.9727, 253.9727, 253.9729, 253.9729, 253.9731, 253.973, 
    253.9734, 253.9733, 253.9736, 253.9735, 253.9736, 253.9736, 253.9736, 
    253.9735, 253.9735, 253.9734, 253.973, 253.9731, 253.9728, 253.9726, 
    253.9724, 253.9723, 253.9724, 253.9724, 253.9725, 253.9726, 253.9727, 
    253.9728, 253.9729, 253.9731, 253.9732, 253.9734, 253.9734, 253.9734, 
    253.9735, 253.9736, 253.9736, 253.9736, 253.9734, 253.9736, 253.9733, 
    253.9734, 253.9729, 253.9727, 253.9726, 253.9725, 253.9724, 253.9725, 
    253.9724, 253.9725, 253.9726, 253.9726, 253.9728, 253.9727, 253.9732, 
    253.973, 253.9735, 253.9734, 253.9735, 253.9734, 253.9736, 253.9735, 
    253.9737, 253.9737, 253.9737, 253.9738, 253.9734, 253.9736, 253.9726, 
    253.9726, 253.9726, 253.9725, 253.9725, 253.9724, 253.9725, 253.9725, 
    253.9726, 253.9727, 253.9727, 253.9729, 253.973, 253.9732, 253.9734, 
    253.9735, 253.9734, 253.9735, 253.9734, 253.9734, 253.9737, 253.9735, 
    253.9738, 253.9738, 253.9736, 253.9738, 253.9726, 253.9726, 253.9724, 
    253.9725, 253.9724, 253.9725, 253.9725, 253.9727, 253.9728, 253.9728, 
    253.9729, 253.973, 253.9732, 253.9734, 253.9735, 253.9735, 253.9735, 
    253.9735, 253.9734, 253.9735, 253.9736, 253.9735, 253.9738, 253.9737, 
    253.9738, 253.9737, 253.9726, 253.9726, 253.9726, 253.9727, 253.9726, 
    253.9728, 253.9729, 253.9731, 253.973, 253.9732, 253.973, 253.973, 
    253.9732, 253.973, 253.9733, 253.9731, 253.9735, 253.9733, 253.9735, 
    253.9735, 253.9736, 253.9736, 253.9737, 253.9739, 253.9738, 253.974, 
    253.9727, 253.9728, 253.9728, 253.9729, 253.9729, 253.973, 253.9732, 
    253.9732, 253.9733, 253.9733, 253.9731, 253.9733, 253.9728, 253.9729, 
    253.9729, 253.9727, 253.9732, 253.9729, 253.9734, 253.9733, 253.9736, 
    253.9734, 253.9738, 253.974, 253.9741, 253.9743, 253.9728, 253.9728, 
    253.9729, 253.973, 253.9731, 253.9733, 253.9733, 253.9733, 253.9734, 
    253.9734, 253.9733, 253.9735, 253.9729, 253.9732, 253.9728, 253.9729, 
    253.973, 253.9729, 253.9732, 253.9732, 253.9734, 253.9733, 253.9739, 
    253.9736, 253.9744, 253.9742, 253.9728, 253.9728, 253.9731, 253.9729, 
    253.9733, 253.9733, 253.9734, 253.9735, 253.9735, 253.9736, 253.9735, 
    253.9736, 253.9733, 253.9734, 253.973, 253.9731, 253.9731, 253.973, 
    253.9732, 253.9733, 253.9733, 253.9734, 253.9735, 253.9733, 253.974, 
    253.9735, 253.9729, 253.973, 253.9731, 253.973, 253.9733, 253.9732, 
    253.9736, 253.9735, 253.9736, 253.9735, 253.9735, 253.9734, 253.9734, 
    253.9732, 253.9731, 253.973, 253.973, 253.9731, 253.9733, 253.9735, 
    253.9735, 253.9736, 253.9733, 253.9734, 253.9733, 253.9735, 253.9732, 
    253.9734, 253.9731, 253.9731, 253.9732, 253.9734, 253.9734, 253.9735, 
    253.9735, 253.9733, 253.9733, 253.9732, 253.9732, 253.9731, 253.9731, 
    253.9731, 253.9732, 253.9733, 253.9735, 253.9736, 253.9737, 253.9739, 
    253.9737, 253.974, 253.9737, 253.9741, 253.9734, 253.9737, 253.9732, 
    253.9733, 253.9734, 253.9736, 253.9735, 253.9736, 253.9733, 253.9731, 
    253.9731, 253.973, 253.9731, 253.9731, 253.9732, 253.9731, 253.9733, 
    253.9732, 253.9735, 253.9736, 253.9739, 253.9741, 253.9743, 253.9744, 
    253.9744, 253.9744 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  253.9724, 253.9726, 253.9725, 253.9727, 253.9726, 253.9727, 253.9724, 
    253.9726, 253.9725, 253.9724, 253.9729, 253.9727, 253.9732, 253.973, 
    253.9734, 253.9732, 253.9735, 253.9734, 253.9736, 253.9736, 253.9738, 
    253.9737, 253.974, 253.9738, 253.9738, 253.9737, 253.9727, 253.9729, 
    253.9727, 253.9727, 253.9727, 253.9726, 253.9725, 253.9724, 253.9724, 
    253.9725, 253.9727, 253.9727, 253.9729, 253.9729, 253.9731, 253.973, 
    253.9734, 253.9733, 253.9736, 253.9735, 253.9736, 253.9736, 253.9736, 
    253.9735, 253.9735, 253.9734, 253.973, 253.9731, 253.9728, 253.9726, 
    253.9724, 253.9723, 253.9724, 253.9724, 253.9725, 253.9726, 253.9727, 
    253.9728, 253.9729, 253.9731, 253.9732, 253.9734, 253.9734, 253.9734, 
    253.9735, 253.9736, 253.9736, 253.9736, 253.9734, 253.9736, 253.9733, 
    253.9734, 253.9729, 253.9727, 253.9726, 253.9725, 253.9724, 253.9725, 
    253.9724, 253.9725, 253.9726, 253.9726, 253.9728, 253.9727, 253.9732, 
    253.973, 253.9735, 253.9734, 253.9735, 253.9734, 253.9736, 253.9735, 
    253.9737, 253.9737, 253.9737, 253.9738, 253.9734, 253.9736, 253.9726, 
    253.9726, 253.9726, 253.9725, 253.9725, 253.9724, 253.9725, 253.9725, 
    253.9726, 253.9727, 253.9727, 253.9729, 253.973, 253.9732, 253.9734, 
    253.9735, 253.9734, 253.9735, 253.9734, 253.9734, 253.9737, 253.9735, 
    253.9738, 253.9738, 253.9736, 253.9738, 253.9726, 253.9726, 253.9724, 
    253.9725, 253.9724, 253.9725, 253.9725, 253.9727, 253.9728, 253.9728, 
    253.9729, 253.973, 253.9732, 253.9734, 253.9735, 253.9735, 253.9735, 
    253.9735, 253.9734, 253.9735, 253.9736, 253.9735, 253.9738, 253.9737, 
    253.9738, 253.9737, 253.9726, 253.9726, 253.9726, 253.9727, 253.9726, 
    253.9728, 253.9729, 253.9731, 253.973, 253.9732, 253.973, 253.973, 
    253.9732, 253.973, 253.9733, 253.9731, 253.9735, 253.9733, 253.9735, 
    253.9735, 253.9736, 253.9736, 253.9737, 253.9739, 253.9738, 253.974, 
    253.9727, 253.9728, 253.9728, 253.9729, 253.9729, 253.973, 253.9732, 
    253.9732, 253.9733, 253.9733, 253.9731, 253.9733, 253.9728, 253.9729, 
    253.9729, 253.9727, 253.9732, 253.9729, 253.9734, 253.9733, 253.9736, 
    253.9734, 253.9738, 253.974, 253.9741, 253.9743, 253.9728, 253.9728, 
    253.9729, 253.973, 253.9731, 253.9733, 253.9733, 253.9733, 253.9734, 
    253.9734, 253.9733, 253.9735, 253.9729, 253.9732, 253.9728, 253.9729, 
    253.973, 253.9729, 253.9732, 253.9732, 253.9734, 253.9733, 253.9739, 
    253.9736, 253.9744, 253.9742, 253.9728, 253.9728, 253.9731, 253.9729, 
    253.9733, 253.9733, 253.9734, 253.9735, 253.9735, 253.9736, 253.9735, 
    253.9736, 253.9733, 253.9734, 253.973, 253.9731, 253.9731, 253.973, 
    253.9732, 253.9733, 253.9733, 253.9734, 253.9735, 253.9733, 253.974, 
    253.9735, 253.9729, 253.973, 253.9731, 253.973, 253.9733, 253.9732, 
    253.9736, 253.9735, 253.9736, 253.9735, 253.9735, 253.9734, 253.9734, 
    253.9732, 253.9731, 253.973, 253.973, 253.9731, 253.9733, 253.9735, 
    253.9735, 253.9736, 253.9733, 253.9734, 253.9733, 253.9735, 253.9732, 
    253.9734, 253.9731, 253.9731, 253.9732, 253.9734, 253.9734, 253.9735, 
    253.9735, 253.9733, 253.9733, 253.9732, 253.9732, 253.9731, 253.9731, 
    253.9731, 253.9732, 253.9733, 253.9735, 253.9736, 253.9737, 253.9739, 
    253.9737, 253.974, 253.9737, 253.9741, 253.9734, 253.9737, 253.9732, 
    253.9733, 253.9734, 253.9736, 253.9735, 253.9736, 253.9733, 253.9731, 
    253.9731, 253.973, 253.9731, 253.9731, 253.9732, 253.9731, 253.9733, 
    253.9732, 253.9735, 253.9736, 253.9739, 253.9741, 253.9743, 253.9744, 
    253.9744, 253.9744 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  254.5119, 254.5134, 254.5131, 254.5143, 254.5137, 254.5145, 254.5122, 
    254.5135, 254.5127, 254.5121, 254.5166, 254.5144, 254.5191, 254.5177, 
    254.5214, 254.5189, 254.5219, 254.5213, 254.5231, 254.5226, 254.5247, 
    254.5233, 254.5259, 254.5244, 254.5246, 254.5232, 254.5149, 254.5164, 
    254.5148, 254.515, 254.5149, 254.5137, 254.5131, 254.5118, 254.5121, 
    254.513, 254.5151, 254.5144, 254.5162, 254.5162, 254.5182, 254.5173, 
    254.5207, 254.5198, 254.5226, 254.5219, 254.5226, 254.5224, 254.5226, 
    254.5215, 254.522, 254.521, 254.5175, 254.5185, 254.5154, 254.5135, 
    254.5123, 254.5114, 254.5116, 254.5118, 254.513, 254.5141, 254.515, 
    254.5156, 254.5162, 254.5179, 254.5188, 254.5209, 254.5206, 254.5212, 
    254.5218, 254.5228, 254.5227, 254.5231, 254.5212, 254.5224, 254.5203, 
    254.5209, 254.5162, 254.5146, 254.5138, 254.5132, 254.5116, 254.5127, 
    254.5123, 254.5133, 254.514, 254.5136, 254.5156, 254.5148, 254.5189, 
    254.5171, 254.5217, 254.5206, 254.522, 254.5213, 254.5225, 254.5214, 
    254.5233, 254.5237, 254.5234, 254.5245, 254.5214, 254.5225, 254.5136, 
    254.5137, 254.5139, 254.5128, 254.5128, 254.5118, 254.5127, 254.513, 
    254.514, 254.5145, 254.5151, 254.5162, 254.5175, 254.5194, 254.5207, 
    254.5216, 254.5211, 254.5215, 254.521, 254.5207, 254.5235, 254.5219, 
    254.5243, 254.5242, 254.5231, 254.5242, 254.5137, 254.5134, 254.5124, 
    254.5132, 254.5117, 254.5125, 254.513, 254.5148, 254.5153, 254.5156, 
    254.5164, 254.5173, 254.519, 254.5205, 254.5218, 254.5217, 254.5218, 
    254.5221, 254.5213, 254.5222, 254.5223, 254.522, 254.5242, 254.5236, 
    254.5242, 254.5238, 254.5135, 254.514, 254.5137, 254.5143, 254.5139, 
    254.5155, 254.5159, 254.5182, 254.5173, 254.5188, 254.5175, 254.5177, 
    254.5188, 254.5175, 254.5204, 254.5184, 254.5221, 254.5201, 254.5222, 
    254.5218, 254.5225, 254.523, 254.5237, 254.525, 254.5247, 254.5258, 
    254.5148, 254.5154, 254.5154, 254.5161, 254.5166, 254.5177, 254.5194, 
    254.5188, 254.52, 254.5202, 254.5184, 254.5195, 254.5159, 254.5164, 
    254.5161, 254.5148, 254.5189, 254.5168, 254.5207, 254.5196, 254.5229, 
    254.5212, 254.5246, 254.5259, 254.5273, 254.5288, 254.5158, 254.5154, 
    254.5161, 254.5172, 254.5183, 254.5196, 254.5198, 254.52, 254.5207, 
    254.5213, 254.5201, 254.5214, 254.5165, 254.5191, 254.5152, 254.5163, 
    254.5172, 254.5168, 254.5187, 254.5191, 254.5209, 254.52, 254.5256, 
    254.5231, 254.53, 254.5281, 254.5152, 254.5158, 254.5179, 254.5169, 
    254.5197, 254.5204, 254.521, 254.5217, 254.5218, 254.5223, 254.5216, 
    254.5222, 254.5196, 254.5208, 254.5176, 254.5184, 254.5181, 254.5177, 
    254.5189, 254.5201, 254.5202, 254.5206, 254.5216, 254.5197, 254.5258, 
    254.522, 254.5164, 254.5176, 254.5178, 254.5173, 254.5204, 254.5193, 
    254.5222, 254.5215, 254.5228, 254.5221, 254.522, 254.5212, 254.5206, 
    254.5193, 254.5182, 254.5174, 254.5176, 254.5185, 254.5202, 254.5218, 
    254.5215, 254.5227, 254.5195, 254.5208, 254.5203, 254.5217, 254.5188, 
    254.5211, 254.5181, 254.5184, 254.5192, 254.5209, 254.5213, 254.5217, 
    254.5215, 254.5202, 254.5201, 254.5192, 254.519, 254.5183, 254.5178, 
    254.5183, 254.5188, 254.5203, 254.5216, 254.523, 254.5234, 254.525, 
    254.5237, 254.5258, 254.5239, 254.5273, 254.5213, 254.5239, 254.5193, 
    254.5198, 254.5207, 254.5228, 254.5217, 254.5229, 254.5201, 254.5185, 
    254.5182, 254.5174, 254.5182, 254.5181, 254.5188, 254.5186, 254.5203, 
    254.5194, 254.522, 254.5229, 254.5257, 254.5273, 254.5291, 254.5298, 
    254.5301, 254.5302,
  255.6251, 255.6266, 255.6263, 255.6275, 255.6269, 255.6277, 255.6254, 
    255.6267, 255.6259, 255.6253, 255.6299, 255.6276, 255.6323, 255.6309, 
    255.6346, 255.6321, 255.6351, 255.6346, 255.6363, 255.6358, 255.638, 
    255.6366, 255.6392, 255.6377, 255.6379, 255.6365, 255.6281, 255.6296, 
    255.628, 255.6282, 255.6281, 255.6269, 255.6263, 255.625, 255.6252, 
    255.6262, 255.6283, 255.6276, 255.6294, 255.6294, 255.6314, 255.6305, 
    255.634, 255.633, 255.6358, 255.6351, 255.6358, 255.6356, 255.6358, 
    255.6348, 255.6352, 255.6343, 255.6307, 255.6317, 255.6286, 255.6267, 
    255.6255, 255.6246, 255.6247, 255.625, 255.6262, 255.6273, 255.6282, 
    255.6288, 255.6294, 255.6311, 255.632, 255.6341, 255.6338, 255.6344, 
    255.635, 255.6361, 255.6359, 255.6364, 255.6344, 255.6357, 255.6336, 
    255.6342, 255.6294, 255.6278, 255.627, 255.6264, 255.6248, 255.6259, 
    255.6255, 255.6265, 255.6272, 255.6268, 255.6288, 255.628, 255.6321, 
    255.6303, 255.635, 255.6339, 255.6352, 255.6345, 255.6357, 255.6347, 
    255.6365, 255.6369, 255.6367, 255.6378, 255.6346, 255.6358, 255.6268, 
    255.6269, 255.6271, 255.626, 255.626, 255.625, 255.6259, 255.6262, 
    255.6272, 255.6277, 255.6283, 255.6294, 255.6307, 255.6326, 255.6339, 
    255.6348, 255.6343, 255.6348, 255.6342, 255.634, 255.6368, 255.6352, 
    255.6376, 255.6375, 255.6364, 255.6375, 255.6269, 255.6266, 255.6256, 
    255.6264, 255.6249, 255.6257, 255.6262, 255.628, 255.6285, 255.6288, 
    255.6296, 255.6305, 255.6322, 255.6337, 255.6351, 255.635, 255.635, 
    255.6353, 255.6346, 255.6354, 255.6356, 255.6352, 255.6375, 255.6368, 
    255.6375, 255.6371, 255.6267, 255.6272, 255.6269, 255.6274, 255.6271, 
    255.6287, 255.6292, 255.6314, 255.6305, 255.632, 255.6307, 255.6309, 
    255.632, 255.6308, 255.6336, 255.6316, 255.6353, 255.6333, 255.6355, 
    255.6351, 255.6357, 255.6363, 255.637, 255.6383, 255.638, 255.6391, 
    255.628, 255.6286, 255.6286, 255.6293, 255.6298, 255.6309, 255.6327, 
    255.632, 255.6332, 255.6335, 255.6316, 255.6327, 255.6291, 255.6296, 
    255.6293, 255.628, 255.6321, 255.63, 255.634, 255.6328, 255.6362, 
    255.6345, 255.6378, 255.6392, 255.6406, 255.6422, 255.629, 255.6285, 
    255.6293, 255.6304, 255.6315, 255.6329, 255.633, 255.6333, 255.6339, 
    255.6345, 255.6333, 255.6347, 255.6297, 255.6323, 255.6284, 255.6295, 
    255.6304, 255.63, 255.6319, 255.6324, 255.6342, 255.6333, 255.6389, 
    255.6364, 255.6434, 255.6414, 255.6284, 255.629, 255.6311, 255.6301, 
    255.633, 255.6337, 255.6343, 255.635, 255.6351, 255.6355, 255.6348, 
    255.6355, 255.6329, 255.634, 255.6308, 255.6316, 255.6313, 255.6309, 
    255.6321, 255.6333, 255.6334, 255.6338, 255.6349, 255.633, 255.6391, 
    255.6353, 255.6296, 255.6308, 255.631, 255.6305, 255.6336, 255.6325, 
    255.6355, 255.6347, 255.636, 255.6354, 255.6353, 255.6344, 255.6339, 
    255.6325, 255.6314, 255.6306, 255.6308, 255.6317, 255.6334, 255.6351, 
    255.6347, 255.6359, 255.6328, 255.6341, 255.6335, 255.6349, 255.632, 
    255.6344, 255.6313, 255.6316, 255.6325, 255.6341, 255.6346, 255.6349, 
    255.6347, 255.6335, 255.6333, 255.6324, 255.6322, 255.6316, 255.631, 
    255.6315, 255.632, 255.6335, 255.6348, 255.6363, 255.6366, 255.6383, 
    255.6369, 255.6391, 255.6372, 255.6406, 255.6346, 255.6372, 255.6325, 
    255.633, 255.6339, 255.636, 255.6349, 255.6362, 255.6333, 255.6317, 
    255.6314, 255.6306, 255.6314, 255.6313, 255.632, 255.6318, 255.6335, 
    255.6326, 255.6353, 255.6362, 255.639, 255.6407, 255.6424, 255.6432, 
    255.6434, 255.6435,
  257.2191, 257.2204, 257.2202, 257.2213, 257.2206, 257.2213, 257.2194, 
    257.2205, 257.2198, 257.2192, 257.2233, 257.2213, 257.2255, 257.2242, 
    257.2276, 257.2253, 257.2281, 257.2275, 257.2291, 257.2287, 257.2307, 
    257.2293, 257.2318, 257.2304, 257.2306, 257.2293, 257.2217, 257.2231, 
    257.2216, 257.2218, 257.2217, 257.2206, 257.2201, 257.219, 257.2192, 
    257.22, 257.2219, 257.2213, 257.2229, 257.2229, 257.2247, 257.2239, 
    257.227, 257.2261, 257.2287, 257.228, 257.2287, 257.2285, 257.2287, 
    257.2277, 257.2281, 257.2273, 257.224, 257.225, 257.2222, 257.2205, 
    257.2194, 257.2186, 257.2188, 257.2189, 257.22, 257.221, 257.2218, 
    257.2224, 257.2229, 257.2244, 257.2253, 257.2272, 257.2268, 257.2274, 
    257.228, 257.2289, 257.2288, 257.2292, 257.2274, 257.2286, 257.2267, 
    257.2272, 257.2229, 257.2215, 257.2208, 257.2202, 257.2188, 257.2198, 
    257.2194, 257.2203, 257.2209, 257.2206, 257.2224, 257.2217, 257.2253, 
    257.2238, 257.2279, 257.2269, 257.2281, 257.2275, 257.2286, 257.2276, 
    257.2293, 257.2297, 257.2294, 257.2304, 257.2276, 257.2286, 257.2206, 
    257.2206, 257.2209, 257.2199, 257.2198, 257.219, 257.2198, 257.2201, 
    257.2209, 257.2214, 257.2219, 257.2229, 257.2241, 257.2258, 257.227, 
    257.2278, 257.2273, 257.2277, 257.2272, 257.227, 257.2296, 257.2281, 
    257.2303, 257.2302, 257.2292, 257.2302, 257.2207, 257.2204, 257.2195, 
    257.2202, 257.2189, 257.2196, 257.22, 257.2217, 257.2221, 257.2224, 
    257.2231, 257.2239, 257.2254, 257.2268, 257.228, 257.2279, 257.228, 
    257.2282, 257.2275, 257.2283, 257.2285, 257.2281, 257.2302, 257.2296, 
    257.2302, 257.2298, 257.2205, 257.2209, 257.2207, 257.2212, 257.2208, 
    257.2223, 257.2227, 257.2247, 257.2239, 257.2252, 257.2241, 257.2242, 
    257.2253, 257.2241, 257.2267, 257.2249, 257.2282, 257.2264, 257.2283, 
    257.228, 257.2286, 257.2291, 257.2297, 257.2309, 257.2307, 257.2316, 
    257.2216, 257.2222, 257.2222, 257.2228, 257.2232, 257.2242, 257.2258, 
    257.2252, 257.2263, 257.2266, 257.2249, 257.2259, 257.2226, 257.2231, 
    257.2228, 257.2216, 257.2253, 257.2234, 257.227, 257.226, 257.229, 
    257.2274, 257.2305, 257.2318, 257.233, 257.2344, 257.2225, 257.2221, 
    257.2228, 257.2238, 257.2248, 257.226, 257.2261, 257.2264, 257.227, 
    257.2275, 257.2264, 257.2276, 257.2232, 257.2255, 257.222, 257.223, 
    257.2238, 257.2234, 257.2252, 257.2256, 257.2272, 257.2263, 257.2314, 
    257.2292, 257.2356, 257.2337, 257.222, 257.2225, 257.2244, 257.2235, 
    257.2261, 257.2267, 257.2273, 257.2279, 257.228, 257.2284, 257.2278, 
    257.2284, 257.226, 257.2271, 257.2242, 257.2249, 257.2246, 257.2242, 
    257.2253, 257.2264, 257.2265, 257.2268, 257.2278, 257.2261, 257.2317, 
    257.2282, 257.2231, 257.2241, 257.2243, 257.2239, 257.2267, 257.2256, 
    257.2284, 257.2277, 257.2289, 257.2283, 257.2282, 257.2274, 257.2269, 
    257.2257, 257.2247, 257.224, 257.2242, 257.225, 257.2265, 257.228, 
    257.2277, 257.2288, 257.2259, 257.2271, 257.2266, 257.2278, 257.2252, 
    257.2274, 257.2246, 257.2249, 257.2256, 257.2271, 257.2275, 257.2279, 
    257.2277, 257.2266, 257.2264, 257.2256, 257.2254, 257.2248, 257.2244, 
    257.2248, 257.2253, 257.2266, 257.2278, 257.2291, 257.2294, 257.2309, 
    257.2297, 257.2317, 257.2299, 257.233, 257.2275, 257.2299, 257.2257, 
    257.2261, 257.2269, 257.2289, 257.2278, 257.229, 257.2264, 257.225, 
    257.2247, 257.224, 257.2247, 257.2246, 257.2253, 257.2251, 257.2266, 
    257.2258, 257.2281, 257.229, 257.2315, 257.2331, 257.2346, 257.2354, 
    257.2356, 257.2357,
  259.3044, 259.3054, 259.3052, 259.306, 259.3055, 259.3061, 259.3046, 
    259.3054, 259.3049, 259.3045, 259.3075, 259.306, 259.3091, 259.3081, 
    259.3106, 259.3089, 259.3109, 259.3105, 259.3117, 259.3114, 259.3128, 
    259.3119, 259.3136, 259.3126, 259.3128, 259.3118, 259.3063, 259.3073, 
    259.3062, 259.3064, 259.3063, 259.3055, 259.3051, 259.3044, 259.3045, 
    259.3051, 259.3065, 259.306, 259.3072, 259.3072, 259.3085, 259.3079, 
    259.3102, 259.3095, 259.3114, 259.3109, 259.3114, 259.3112, 259.3114, 
    259.3107, 259.3109, 259.3103, 259.308, 259.3087, 259.3066, 259.3054, 
    259.3047, 259.3041, 259.3042, 259.3043, 259.3051, 259.3058, 259.3064, 
    259.3068, 259.3072, 259.3083, 259.3089, 259.3103, 259.31, 259.3104, 
    259.3109, 259.3116, 259.3114, 259.3117, 259.3104, 259.3113, 259.3099, 
    259.3103, 259.3072, 259.3061, 259.3056, 259.3052, 259.3042, 259.3049, 
    259.3047, 259.3053, 259.3057, 259.3055, 259.3068, 259.3063, 259.3089, 
    259.3078, 259.3108, 259.3101, 259.311, 259.3105, 259.3113, 259.3106, 
    259.3119, 259.3121, 259.3119, 259.3127, 259.3105, 259.3113, 259.3055, 
    259.3055, 259.3057, 259.305, 259.305, 259.3044, 259.3049, 259.3051, 
    259.3058, 259.3061, 259.3064, 259.3072, 259.308, 259.3092, 259.3101, 
    259.3107, 259.3104, 259.3107, 259.3103, 259.3102, 259.312, 259.3109, 
    259.3126, 259.3125, 259.3117, 259.3125, 259.3056, 259.3054, 259.3047, 
    259.3052, 259.3043, 259.3048, 259.3051, 259.3063, 259.3065, 259.3068, 
    259.3073, 259.3079, 259.309, 259.31, 259.3109, 259.3108, 259.3109, 
    259.311, 259.3105, 259.3111, 259.3112, 259.311, 259.3125, 259.312, 
    259.3125, 259.3122, 259.3055, 259.3058, 259.3056, 259.3059, 259.3057, 
    259.3067, 259.307, 259.3085, 259.3079, 259.3089, 259.308, 259.3081, 
    259.3089, 259.308, 259.3099, 259.3086, 259.311, 259.3097, 259.3111, 
    259.3109, 259.3113, 259.3117, 259.3122, 259.313, 259.3128, 259.3136, 
    259.3062, 259.3067, 259.3066, 259.3071, 259.3074, 259.3081, 259.3093, 
    259.3088, 259.3097, 259.3098, 259.3086, 259.3093, 259.3069, 259.3073, 
    259.3071, 259.3063, 259.3089, 259.3076, 259.3101, 259.3094, 259.3116, 
    259.3105, 259.3127, 259.3136, 259.3146, 259.3156, 259.3069, 259.3066, 
    259.3071, 259.3078, 259.3085, 259.3094, 259.3095, 259.3097, 259.3101, 
    259.3105, 259.3097, 259.3106, 259.3074, 259.3091, 259.3065, 259.3073, 
    259.3078, 259.3076, 259.3088, 259.3091, 259.3103, 259.3097, 259.3134, 
    259.3117, 259.3165, 259.3151, 259.3065, 259.3069, 259.3083, 259.3076, 
    259.3095, 259.3099, 259.3103, 259.3108, 259.3109, 259.3112, 259.3107, 
    259.3112, 259.3094, 259.3102, 259.3081, 259.3086, 259.3084, 259.3081, 
    259.3089, 259.3097, 259.3098, 259.31, 259.3108, 259.3095, 259.3136, 
    259.311, 259.3073, 259.308, 259.3082, 259.3079, 259.3099, 259.3092, 
    259.3112, 259.3106, 259.3115, 259.3111, 259.311, 259.3104, 259.3101, 
    259.3092, 259.3085, 259.308, 259.3081, 259.3087, 259.3098, 259.3109, 
    259.3106, 259.3114, 259.3094, 259.3102, 259.3099, 259.3108, 259.3088, 
    259.3104, 259.3084, 259.3086, 259.3091, 259.3102, 259.3105, 259.3108, 
    259.3106, 259.3098, 259.3097, 259.3091, 259.309, 259.3086, 259.3082, 
    259.3085, 259.3089, 259.3098, 259.3107, 259.3117, 259.3119, 259.313, 
    259.3121, 259.3136, 259.3123, 259.3146, 259.3105, 259.3123, 259.3092, 
    259.3095, 259.3101, 259.3115, 259.3108, 259.3116, 259.3097, 259.3087, 
    259.3084, 259.308, 259.3085, 259.3084, 259.3089, 259.3087, 259.3099, 
    259.3093, 259.311, 259.3116, 259.3135, 259.3146, 259.3158, 259.3163, 
    259.3165, 259.3166,
  261.451, 261.4515, 261.4514, 261.4518, 261.4515, 261.4518, 261.4511, 
    261.4515, 261.4512, 261.4511, 261.4524, 261.4518, 261.4532, 261.4528, 
    261.4539, 261.4531, 261.4541, 261.4539, 261.4545, 261.4543, 261.455, 
    261.4546, 261.4554, 261.4549, 261.455, 261.4545, 261.4519, 261.4524, 
    261.4519, 261.4519, 261.4519, 261.4515, 261.4514, 261.451, 261.451, 
    261.4513, 261.452, 261.4518, 261.4523, 261.4523, 261.4529, 261.4526, 
    261.4537, 261.4534, 261.4543, 261.4541, 261.4543, 261.4543, 261.4543, 
    261.454, 261.4541, 261.4538, 261.4527, 261.453, 261.4521, 261.4515, 
    261.4511, 261.4509, 261.4509, 261.451, 261.4513, 261.4517, 261.4519, 
    261.4521, 261.4523, 261.4528, 261.4531, 261.4538, 261.4537, 261.4539, 
    261.4541, 261.4544, 261.4543, 261.4545, 261.4539, 261.4543, 261.4536, 
    261.4538, 261.4523, 261.4518, 261.4516, 261.4514, 261.4509, 261.4513, 
    261.4511, 261.4514, 261.4516, 261.4515, 261.4521, 261.4519, 261.4531, 
    261.4526, 261.454, 261.4537, 261.4541, 261.4539, 261.4543, 261.4539, 
    261.4546, 261.4547, 261.4546, 261.455, 261.4539, 261.4543, 261.4515, 
    261.4515, 261.4516, 261.4513, 261.4513, 261.451, 261.4512, 261.4514, 
    261.4516, 261.4518, 261.452, 261.4523, 261.4527, 261.4533, 261.4537, 
    261.454, 261.4538, 261.454, 261.4538, 261.4537, 261.4547, 261.4541, 
    261.4549, 261.4549, 261.4545, 261.4549, 261.4515, 261.4515, 261.4511, 
    261.4514, 261.451, 261.4512, 261.4513, 261.4519, 261.452, 261.4521, 
    261.4524, 261.4526, 261.4532, 261.4536, 261.4541, 261.454, 261.4541, 
    261.4542, 261.4539, 261.4542, 261.4543, 261.4541, 261.4549, 261.4547, 
    261.4549, 261.4547, 261.4515, 261.4516, 261.4516, 261.4517, 261.4516, 
    261.4521, 261.4522, 261.4529, 261.4526, 261.4531, 261.4527, 261.4528, 
    261.4531, 261.4527, 261.4536, 261.453, 261.4542, 261.4535, 261.4542, 
    261.4541, 261.4543, 261.4545, 261.4547, 261.4551, 261.455, 261.4554, 
    261.4519, 261.4521, 261.4521, 261.4522, 261.4524, 261.4528, 261.4533, 
    261.4531, 261.4535, 261.4536, 261.453, 261.4533, 261.4522, 261.4524, 
    261.4523, 261.4519, 261.4531, 261.4525, 261.4537, 261.4533, 261.4544, 
    261.4539, 261.455, 261.4554, 261.4559, 261.4565, 261.4522, 261.452, 
    261.4523, 261.4526, 261.4529, 261.4534, 261.4534, 261.4535, 261.4537, 
    261.4539, 261.4535, 261.4539, 261.4524, 261.4532, 261.452, 261.4523, 
    261.4526, 261.4525, 261.4531, 261.4532, 261.4538, 261.4535, 261.4553, 
    261.4545, 261.4569, 261.4562, 261.452, 261.4522, 261.4528, 261.4525, 
    261.4534, 261.4536, 261.4538, 261.454, 261.4541, 261.4542, 261.454, 
    261.4542, 261.4534, 261.4537, 261.4528, 261.453, 261.4529, 261.4528, 
    261.4531, 261.4535, 261.4536, 261.4537, 261.454, 261.4534, 261.4554, 
    261.4541, 261.4524, 261.4527, 261.4528, 261.4526, 261.4536, 261.4532, 
    261.4542, 261.4539, 261.4544, 261.4542, 261.4541, 261.4539, 261.4537, 
    261.4533, 261.4529, 261.4527, 261.4527, 261.453, 261.4536, 261.4541, 
    261.4539, 261.4543, 261.4533, 261.4538, 261.4536, 261.454, 261.4531, 
    261.4539, 261.4529, 261.453, 261.4532, 261.4538, 261.4539, 261.454, 
    261.4539, 261.4536, 261.4535, 261.4532, 261.4532, 261.453, 261.4528, 
    261.4529, 261.4531, 261.4536, 261.454, 261.4545, 261.4546, 261.4551, 
    261.4547, 261.4554, 261.4548, 261.4559, 261.4539, 261.4548, 261.4532, 
    261.4534, 261.4537, 261.4544, 261.454, 261.4544, 261.4535, 261.453, 
    261.4529, 261.4527, 261.4529, 261.4529, 261.4531, 261.453, 261.4536, 
    261.4533, 261.4541, 261.4544, 261.4554, 261.4559, 261.4565, 261.4568, 
    261.4569, 261.4569,
  262.7756, 262.7757, 262.7757, 262.7758, 262.7757, 262.7758, 262.7756, 
    262.7757, 262.7756, 262.7756, 262.7759, 262.7758, 262.7761, 262.776, 
    262.7763, 262.7761, 262.7763, 262.7763, 262.7764, 262.7764, 262.7766, 
    262.7764, 262.7766, 262.7765, 262.7766, 262.7764, 262.7758, 262.7759, 
    262.7758, 262.7758, 262.7758, 262.7757, 262.7757, 262.7756, 262.7756, 
    262.7757, 262.7758, 262.7758, 262.7759, 262.7759, 262.776, 262.776, 
    262.7762, 262.7762, 262.7764, 262.7763, 262.7764, 262.7763, 262.7764, 
    262.7763, 262.7763, 262.7762, 262.776, 262.7761, 262.7758, 262.7757, 
    262.7756, 262.7756, 262.7756, 262.7756, 262.7757, 262.7758, 262.7758, 
    262.7758, 262.7759, 262.776, 262.7761, 262.7762, 262.7762, 262.7762, 
    262.7763, 262.7764, 262.7764, 262.7764, 262.7762, 262.7764, 262.7762, 
    262.7762, 262.7759, 262.7758, 262.7757, 262.7757, 262.7756, 262.7756, 
    262.7756, 262.7757, 262.7757, 262.7757, 262.7758, 262.7758, 262.7761, 
    262.7759, 262.7763, 262.7762, 262.7763, 262.7763, 262.7764, 262.7763, 
    262.7764, 262.7765, 262.7764, 262.7765, 262.7763, 262.7764, 262.7757, 
    262.7757, 262.7757, 262.7757, 262.7757, 262.7756, 262.7756, 262.7757, 
    262.7757, 262.7758, 262.7758, 262.7759, 262.776, 262.7761, 262.7762, 
    262.7763, 262.7762, 262.7763, 262.7762, 262.7762, 262.7764, 262.7763, 
    262.7765, 262.7765, 262.7764, 262.7765, 262.7757, 262.7757, 262.7756, 
    262.7757, 262.7756, 262.7756, 262.7757, 262.7758, 262.7758, 262.7758, 
    262.7759, 262.776, 262.7761, 262.7762, 262.7763, 262.7763, 262.7763, 
    262.7763, 262.7763, 262.7763, 262.7763, 262.7763, 262.7765, 262.7765, 
    262.7765, 262.7765, 262.7757, 262.7757, 262.7757, 262.7758, 262.7757, 
    262.7758, 262.7759, 262.776, 262.776, 262.7761, 262.776, 262.776, 
    262.7761, 262.776, 262.7762, 262.776, 262.7763, 262.7762, 262.7763, 
    262.7763, 262.7764, 262.7764, 262.7765, 262.7766, 262.7766, 262.7766, 
    262.7758, 262.7758, 262.7758, 262.7759, 262.7759, 262.776, 262.7761, 
    262.7761, 262.7762, 262.7762, 262.776, 262.7761, 262.7758, 262.7759, 
    262.7759, 262.7758, 262.7761, 262.7759, 262.7762, 262.7761, 262.7764, 
    262.7762, 262.7765, 262.7766, 262.7768, 262.7769, 262.7758, 262.7758, 
    262.7759, 262.776, 262.776, 262.7761, 262.7762, 262.7762, 262.7762, 
    262.7763, 262.7762, 262.7763, 262.7759, 262.7761, 262.7758, 262.7759, 
    262.7759, 262.7759, 262.7761, 262.7761, 262.7762, 262.7762, 262.7766, 
    262.7764, 262.777, 262.7768, 262.7758, 262.7758, 262.776, 262.7759, 
    262.7762, 262.7762, 262.7762, 262.7763, 262.7763, 262.7763, 262.7763, 
    262.7763, 262.7761, 262.7762, 262.776, 262.776, 262.776, 262.776, 
    262.7761, 262.7762, 262.7762, 262.7762, 262.7763, 262.7762, 262.7766, 
    262.7763, 262.7759, 262.776, 262.776, 262.776, 262.7762, 262.7761, 
    262.7763, 262.7763, 262.7764, 262.7763, 262.7763, 262.7762, 262.7762, 
    262.7761, 262.776, 262.776, 262.776, 262.7761, 262.7762, 262.7763, 
    262.7763, 262.7764, 262.7761, 262.7762, 262.7762, 262.7763, 262.7761, 
    262.7762, 262.776, 262.776, 262.7761, 262.7762, 262.7763, 262.7763, 
    262.7763, 262.7762, 262.7762, 262.7761, 262.7761, 262.776, 262.776, 
    262.776, 262.7761, 262.7762, 262.7763, 262.7764, 262.7764, 262.7766, 
    262.7765, 262.7766, 262.7765, 262.7768, 262.7763, 262.7765, 262.7761, 
    262.7762, 262.7762, 262.7764, 262.7763, 262.7764, 262.7762, 262.7761, 
    262.776, 262.776, 262.776, 262.776, 262.7761, 262.7761, 262.7762, 
    262.7761, 262.7763, 262.7764, 262.7766, 262.7768, 262.7769, 262.777, 
    262.777, 262.777,
  263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1192, 263.1191, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1192, 
    263.1191, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1191, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1192, 263.1191, 263.1191, 
    263.1192, 263.1191, 263.1192, 263.1191, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1191, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1191, 263.1192, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1192, 263.1191, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1193, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1191, 263.1192, 263.1191, 263.1191, 
    263.1191, 263.1191, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1193, 263.1193, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1191, 263.1191, 263.1191, 263.1191, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1191, 263.1191, 263.1191, 263.1191, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1191, 263.1191, 263.1191, 263.1191, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1191, 263.1191, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1191, 263.1191, 
    263.1191, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1191, 
    263.1191, 263.1191, 263.1191, 263.1191, 263.1192, 263.1192, 263.1192, 
    263.1192, 263.1192, 263.1192, 263.1192, 263.1192, 263.1193, 263.1193, 
    263.1193, 263.1193,
  263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 263.1492, 
    263.1492, 263.1492,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.0843, 263.0988, 263.096, 263.1076, 263.1012, 263.1088, 263.0873, 
    263.0994, 263.0916, 263.0856, 263.1302, 263.1082, 263.153, 263.139, 
    263.174, 263.1508, 263.1787, 263.1733, 263.1894, 263.1848, 263.2047, 
    263.1915, 263.2154, 263.2015, 263.2036, 263.1911, 263.1126, 263.1274, 
    263.1118, 263.1139, 263.1129, 263.1013, 263.0955, 263.0832, 263.0854, 
    263.0945, 263.1148, 263.1079, 263.1253, 263.1249, 263.1442, 263.1355, 
    263.1678, 263.1586, 263.185, 263.1784, 263.1847, 263.1828, 263.1847, 
    263.175, 263.1792, 263.1706, 263.1371, 263.147, 263.1175, 263.0996, 
    263.0878, 263.0794, 263.0806, 263.0828, 263.0945, 263.1055, 263.1138, 
    263.1194, 263.1249, 263.1414, 263.1501, 263.1696, 263.1661, 263.172, 
    263.1777, 263.1872, 263.1857, 263.1898, 263.1719, 263.1838, 263.1641, 
    263.1695, 263.1263, 263.1098, 263.1027, 263.0965, 263.0815, 263.0919, 
    263.0878, 263.0975, 263.1037, 263.1007, 263.1195, 263.1122, 263.1506, 
    263.1342, 263.1771, 263.1668, 263.1795, 263.173, 263.1841, 263.1741, 
    263.1914, 263.1946, 263.1926, 263.2019, 263.1736, 263.1847, 263.1006, 
    263.1011, 263.1034, 263.0932, 263.0925, 263.0832, 263.0915, 263.0951, 
    263.1041, 263.1094, 263.1145, 263.1256, 263.1379, 263.1552, 263.1675, 
    263.1757, 263.1707, 263.1751, 263.1702, 263.1678, 263.1932, 263.1792, 
    263.2005, 263.1993, 263.19, 263.1994, 263.1014, 263.0986, 263.0886, 
    263.0964, 263.0822, 263.0901, 263.0947, 263.1123, 263.1162, 263.1198, 
    263.1269, 263.136, 263.1518, 263.1655, 263.178, 263.1771, 263.1775, 
    263.1802, 263.1733, 263.1814, 263.1827, 263.1792, 263.1992, 263.1933, 
    263.1993, 263.1955, 263.0995, 263.1043, 263.1017, 263.1066, 263.1031, 
    263.1185, 263.1231, 263.1446, 263.1358, 263.1497, 263.1372, 263.1394, 
    263.1501, 263.1379, 263.1648, 263.1465, 263.1804, 263.1622, 263.1815, 
    263.178, 263.1838, 263.189, 263.1949, 263.2069, 263.2042, 263.2142, 
    263.1115, 263.1178, 263.1172, 263.1238, 263.1286, 263.1391, 263.1557, 
    263.1495, 263.161, 263.1633, 263.1458, 263.1565, 263.1219, 263.1276, 
    263.1242, 263.112, 263.1509, 263.131, 263.1677, 263.157, 263.1882, 
    263.1727, 263.2026, 263.2156, 263.2278, 263.2421, 263.1212, 263.1169, 
    263.1245, 263.135, 263.1447, 263.1576, 263.1589, 263.1613, 263.1676, 
    263.1728, 263.1621, 263.1741, 263.1288, 263.1526, 263.1153, 263.1266, 
    263.1344, 263.131, 263.1488, 263.1529, 263.1698, 263.1611, 263.2124, 
    263.19, 263.2529, 263.2352, 263.1154, 263.1212, 263.141, 263.1316, 
    263.1585, 263.1651, 263.1704, 263.1772, 263.178, 263.182, 263.1754, 
    263.1818, 263.1576, 263.1684, 263.1388, 263.146, 263.1427, 263.139, 
    263.1503, 263.1622, 263.1625, 263.1664, 263.1771, 263.1586, 263.2153, 
    263.1805, 263.1274, 263.1384, 263.14, 263.1357, 263.1644, 263.154, 
    263.1819, 263.1744, 263.1867, 263.1806, 263.1797, 263.1718, 263.1669, 
    263.1545, 263.1444, 263.1364, 263.1382, 263.147, 263.163, 263.178, 
    263.1747, 263.1858, 263.1565, 263.1688, 263.1641, 263.1765, 263.1493, 
    263.1724, 263.1434, 263.1459, 263.1538, 263.1696, 263.1732, 263.1769, 
    263.1746, 263.1634, 263.1616, 263.1536, 263.1514, 263.1454, 263.1404, 
    263.1449, 263.1497, 263.1634, 263.1757, 263.189, 263.1923, 263.2073, 
    263.1946, 263.2155, 263.1977, 263.2285, 263.1737, 263.1972, 263.1542, 
    263.1589, 263.1674, 263.1869, 263.1764, 263.1887, 263.1615, 263.1473, 
    263.1437, 263.1368, 263.1438, 263.1432, 263.15, 263.1478, 263.1638, 
    263.1552, 263.1797, 263.1886, 263.2131, 263.2285, 263.2441, 263.2509, 
    263.2531, 263.2539 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9727, 253.9735, 253.9734, 253.974, 253.9737, 253.9741, 253.9729, 
    253.9736, 253.9731, 253.9728, 253.9753, 253.9741, 253.9767, 253.9759, 
    253.9779, 253.9765, 253.9782, 253.9779, 253.9789, 253.9786, 253.9798, 
    253.979, 253.9804, 253.9796, 253.9797, 253.979, 253.9743, 253.9752, 
    253.9743, 253.9744, 253.9744, 253.9737, 253.9733, 253.9727, 253.9728, 
    253.9733, 253.9745, 253.9741, 253.9751, 253.9751, 253.9762, 253.9757, 
    253.9776, 253.977, 253.9786, 253.9782, 253.9786, 253.9785, 253.9786, 
    253.978, 253.9782, 253.9777, 253.9758, 253.9763, 253.9746, 253.9736, 
    253.9729, 253.9724, 253.9725, 253.9726, 253.9733, 253.9739, 253.9744, 
    253.9747, 253.9751, 253.976, 253.9765, 253.9777, 253.9775, 253.9778, 
    253.9782, 253.9787, 253.9786, 253.9789, 253.9778, 253.9785, 253.9774, 
    253.9777, 253.9751, 253.9742, 253.9738, 253.9734, 253.9725, 253.9731, 
    253.9729, 253.9735, 253.9738, 253.9737, 253.9747, 253.9743, 253.9765, 
    253.9756, 253.9781, 253.9775, 253.9783, 253.9779, 253.9785, 253.978, 
    253.979, 253.9792, 253.979, 253.9796, 253.9779, 253.9786, 253.9736, 
    253.9737, 253.9738, 253.9732, 253.9732, 253.9727, 253.9731, 253.9733, 
    253.9739, 253.9742, 253.9745, 253.9751, 253.9758, 253.9768, 253.9776, 
    253.978, 253.9778, 253.978, 253.9777, 253.9776, 253.9791, 253.9782, 
    253.9796, 253.9795, 253.9789, 253.9795, 253.9737, 253.9735, 253.973, 
    253.9734, 253.9726, 253.9731, 253.9733, 253.9743, 253.9746, 253.9748, 
    253.9752, 253.9757, 253.9766, 253.9774, 253.9782, 253.9781, 253.9781, 
    253.9783, 253.9779, 253.9784, 253.9785, 253.9783, 253.9795, 253.9791, 
    253.9795, 253.9792, 253.9736, 253.9739, 253.9737, 253.974, 253.9738, 
    253.9747, 253.9749, 253.9762, 253.9757, 253.9765, 253.9758, 253.9759, 
    253.9765, 253.9758, 253.9774, 253.9763, 253.9783, 253.9772, 253.9784, 
    253.9782, 253.9785, 253.9788, 253.9792, 253.9799, 253.9798, 253.9804, 
    253.9743, 253.9746, 253.9746, 253.975, 253.9753, 253.9759, 253.9769, 
    253.9765, 253.9772, 253.9773, 253.9763, 253.9769, 253.9749, 253.9752, 
    253.975, 253.9743, 253.9766, 253.9754, 253.9776, 253.9769, 253.9788, 
    253.9778, 253.9797, 253.9804, 253.9812, 253.982, 253.9748, 253.9746, 
    253.975, 253.9756, 253.9762, 253.977, 253.9771, 253.9772, 253.9776, 
    253.9779, 253.9772, 253.978, 253.9753, 253.9767, 253.9745, 253.9751, 
    253.9756, 253.9754, 253.9765, 253.9767, 253.9777, 253.9772, 253.9802, 
    253.9789, 253.9827, 253.9816, 253.9745, 253.9749, 253.976, 253.9754, 
    253.977, 253.9774, 253.9777, 253.9781, 253.9782, 253.9784, 253.978, 
    253.9784, 253.977, 253.9776, 253.9759, 253.9763, 253.9761, 253.9759, 
    253.9765, 253.9772, 253.9773, 253.9775, 253.9781, 253.977, 253.9804, 
    253.9783, 253.9752, 253.9758, 253.9759, 253.9757, 253.9774, 253.9768, 
    253.9784, 253.978, 253.9787, 253.9783, 253.9783, 253.9778, 253.9775, 
    253.9768, 253.9762, 253.9757, 253.9758, 253.9763, 253.9773, 253.9782, 
    253.978, 253.9786, 253.9769, 253.9776, 253.9773, 253.9781, 253.9765, 
    253.9778, 253.9761, 253.9763, 253.9767, 253.9777, 253.9779, 253.9781, 
    253.978, 253.9773, 253.9772, 253.9767, 253.9766, 253.9763, 253.976, 
    253.9762, 253.9765, 253.9773, 253.978, 253.9788, 253.979, 253.9799, 
    253.9792, 253.9804, 253.9793, 253.9812, 253.9779, 253.9793, 253.9768, 
    253.9771, 253.9775, 253.9787, 253.9781, 253.9788, 253.9772, 253.9763, 
    253.9762, 253.9758, 253.9762, 253.9761, 253.9765, 253.9764, 253.9773, 
    253.9768, 253.9783, 253.9788, 253.9803, 253.9812, 253.9822, 253.9826, 
    253.9827, 253.9828 ;

 TWS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 T_SCALAR =
  0.1407037, 0.1407121, 0.1407105, 0.1407173, 0.1407136, 0.1407179, 
    0.1407055, 0.1407124, 0.140708, 0.1407045, 0.1407302, 0.1407176, 
    0.140744, 0.1407358, 0.1407567, 0.1407426, 0.1407595, 0.1407564, 
    0.1407662, 0.1407634, 0.1407756, 0.1407675, 0.1407822, 0.1407738, 
    0.140775, 0.1407672, 0.1407203, 0.1407285, 0.1407197, 0.1407209, 
    0.1407204, 0.1407136, 0.14071, 0.1407031, 0.1407044, 0.1407095, 
    0.1407215, 0.1407175, 0.1407278, 0.1407275, 0.1407389, 0.1407338, 
    0.140753, 0.1407476, 0.1407635, 0.1407595, 0.1407633, 0.1407622, 
    0.1407633, 0.1407574, 0.1407599, 0.1407548, 0.1407347, 0.1407405, 
    0.1407231, 0.1407124, 0.1407057, 0.1407009, 0.1407016, 0.1407028, 
    0.1407096, 0.1407161, 0.140721, 0.1407243, 0.1407275, 0.1407369, 
    0.1407423, 0.140754, 0.1407521, 0.1407555, 0.1407591, 0.1407648, 
    0.1407639, 0.1407664, 0.1407555, 0.1407627, 0.1407509, 0.1407541, 
    0.1407278, 0.1407186, 0.1407142, 0.1407108, 0.1407021, 0.1407081, 
    0.1407057, 0.1407115, 0.1407151, 0.1407133, 0.1407244, 0.14072, 
    0.1407426, 0.1407329, 0.1407587, 0.1407525, 0.1407602, 0.1407563, 
    0.1407629, 0.1407569, 0.1407674, 0.1407696, 0.140768, 0.1407742, 
    0.1407566, 0.1407632, 0.1407132, 0.1407135, 0.1407149, 0.1407088, 
    0.1407085, 0.1407031, 0.1407079, 0.14071, 0.1407153, 0.1407184, 
    0.1407214, 0.1407279, 0.1407351, 0.1407454, 0.1407529, 0.1407579, 
    0.1407549, 0.1407575, 0.1407545, 0.1407531, 0.1407688, 0.1407599, 
    0.1407733, 0.1407726, 0.1407664, 0.1407727, 0.1407137, 0.1407121, 
    0.1407062, 0.1407108, 0.1407025, 0.1407071, 0.1407097, 0.14072, 
    0.1407224, 0.1407245, 0.1407287, 0.140734, 0.1407434, 0.1407516, 
    0.1407593, 0.1407588, 0.1407589, 0.1407606, 0.1407564, 0.1407613, 
    0.140762, 0.14076, 0.1407725, 0.1407689, 0.1407726, 0.1407703, 0.1407126, 
    0.1407154, 0.1407139, 0.1407167, 0.1407147, 0.1407236, 0.1407263, 
    0.140739, 0.1407339, 0.1407421, 0.1407348, 0.140736, 0.1407422, 
    0.1407352, 0.1407511, 0.1407401, 0.1407607, 0.1407494, 0.1407613, 
    0.1407593, 0.1407628, 0.1407658, 0.1407699, 0.1407771, 0.1407755, 
    0.1407816, 0.1407197, 0.1407232, 0.140723, 0.1407268, 0.1407297, 
    0.1407359, 0.1407458, 0.1407421, 0.140749, 0.1407503, 0.1407399, 
    0.1407462, 0.1407257, 0.1407289, 0.1407271, 0.1407199, 0.1407428, 
    0.1407309, 0.140753, 0.1407465, 0.1407654, 0.1407559, 0.1407745, 
    0.1407822, 0.1407899, 0.1407984, 0.1407253, 0.1407229, 0.1407273, 
    0.1407333, 0.1407392, 0.1407469, 0.1407478, 0.1407492, 0.140753, 
    0.1407561, 0.1407495, 0.1407569, 0.1407294, 0.1407439, 0.1407218, 
    0.1407283, 0.140733, 0.1407311, 0.1407417, 0.1407442, 0.1407542, 
    0.1407491, 0.1407802, 0.1407663, 0.1408053, 0.1407943, 0.140722, 
    0.1407253, 0.140737, 0.1407314, 0.1407475, 0.1407514, 0.1407547, 
    0.1407587, 0.1407592, 0.1407616, 0.1407577, 0.1407615, 0.1407469, 
    0.1407535, 0.1407357, 0.14074, 0.1407381, 0.1407359, 0.1407426, 
    0.1407496, 0.1407499, 0.1407521, 0.1407581, 0.1407476, 0.1407817, 
    0.1407602, 0.140729, 0.1407353, 0.1407364, 0.1407339, 0.140751, 
    0.1407448, 0.1407616, 0.1407571, 0.1407645, 0.1407608, 0.1407603, 
    0.1407555, 0.1407526, 0.140745, 0.140739, 0.1407343, 0.1407354, 
    0.1407406, 0.1407501, 0.1407592, 0.1407572, 0.140764, 0.1407463, 
    0.1407536, 0.1407507, 0.1407583, 0.140742, 0.1407553, 0.1407385, 0.14074, 
    0.1407447, 0.140754, 0.1407563, 0.1407585, 0.1407572, 0.1407503, 
    0.1407493, 0.1407446, 0.1407432, 0.1407397, 0.1407367, 0.1407394, 
    0.1407422, 0.1407504, 0.1407578, 0.1407659, 0.1407679, 0.140777, 
    0.1407694, 0.1407817, 0.1407709, 0.1407899, 0.1407564, 0.140771, 
    0.1407449, 0.1407478, 0.1407527, 0.1407644, 0.1407583, 0.1407655, 
    0.1407493, 0.1407407, 0.1407387, 0.1407346, 0.1407388, 0.1407384, 
    0.1407424, 0.1407411, 0.1407507, 0.1407456, 0.1407602, 0.1407655, 
    0.1407809, 0.1407901, 0.1407999, 0.1408041, 0.1408054, 0.1408059,
  0.1471514, 0.1471603, 0.1471586, 0.1471658, 0.1471619, 0.1471665, 
    0.1471533, 0.1471606, 0.147156, 0.1471523, 0.1471795, 0.1471661, 
    0.1471942, 0.1471855, 0.1472077, 0.1471928, 0.1472108, 0.1472075, 
    0.1472179, 0.1472149, 0.147228, 0.1472193, 0.147235, 0.147226, 0.1472273, 
    0.1472189, 0.147169, 0.1471778, 0.1471684, 0.1471697, 0.1471691, 
    0.1471619, 0.1471581, 0.1471508, 0.1471522, 0.1471576, 0.1471702, 
    0.1471661, 0.147177, 0.1471767, 0.1471888, 0.1471833, 0.1472038, 
    0.147198, 0.147215, 0.1472107, 0.1472148, 0.1472136, 0.1472148, 
    0.1472085, 0.1472112, 0.1472057, 0.1471843, 0.1471905, 0.147172, 
    0.1471606, 0.1471535, 0.1471484, 0.1471491, 0.1471505, 0.1471576, 
    0.1471645, 0.1471698, 0.1471732, 0.1471767, 0.1471867, 0.1471924, 
    0.1472049, 0.1472028, 0.1472065, 0.1472103, 0.1472164, 0.1472154, 
    0.1472181, 0.1472065, 0.1472142, 0.1472016, 0.147205, 0.147177, 
    0.1471672, 0.1471626, 0.1471589, 0.1471497, 0.147156, 0.1471535, 
    0.1471596, 0.1471634, 0.1471616, 0.1471733, 0.1471687, 0.1471927, 
    0.1471824, 0.1472099, 0.1472033, 0.1472114, 0.1472073, 0.1472144, 
    0.147208, 0.1472191, 0.1472216, 0.1472199, 0.1472264, 0.1472076, 
    0.1472147, 0.1471615, 0.1471618, 0.1471633, 0.1471568, 0.1471564, 
    0.1471507, 0.1471559, 0.147158, 0.1471637, 0.147167, 0.1471701, 
    0.1471771, 0.1471847, 0.1471957, 0.1472037, 0.147209, 0.1472058, 
    0.1472086, 0.1472054, 0.147204, 0.1472207, 0.1472112, 0.1472255, 
    0.1472247, 0.1472181, 0.1472248, 0.147162, 0.1471603, 0.147154, 
    0.1471589, 0.1471501, 0.147155, 0.1471577, 0.1471687, 0.1471712, 
    0.1471734, 0.1471779, 0.1471836, 0.1471936, 0.1472024, 0.1472105, 
    0.1472099, 0.1472102, 0.1472119, 0.1472075, 0.1472127, 0.1472135, 
    0.1472112, 0.1472246, 0.1472208, 0.1472247, 0.1472222, 0.1471609, 
    0.1471638, 0.1471622, 0.1471652, 0.147163, 0.1471725, 0.1471754, 
    0.1471889, 0.1471835, 0.1471922, 0.1471844, 0.1471857, 0.1471923, 
    0.1471848, 0.1472018, 0.1471901, 0.147212, 0.1472, 0.1472127, 0.1472105, 
    0.1472142, 0.1472175, 0.1472219, 0.1472296, 0.1472278, 0.1472344, 
    0.1471683, 0.1471721, 0.1471719, 0.147176, 0.1471789, 0.1471856, 
    0.1471961, 0.1471922, 0.1471995, 0.147201, 0.1471899, 0.1471966, 
    0.1471747, 0.1471781, 0.1471762, 0.1471685, 0.1471929, 0.1471803, 
    0.1472038, 0.1471969, 0.1472171, 0.1472069, 0.1472268, 0.147235, 
    0.1472433, 0.1472525, 0.1471743, 0.1471717, 0.1471765, 0.1471829, 
    0.1471891, 0.1471973, 0.1471982, 0.1471997, 0.1472038, 0.1472071, 
    0.1472001, 0.147208, 0.1471787, 0.1471941, 0.1471706, 0.1471775, 
    0.1471825, 0.1471805, 0.1471918, 0.1471944, 0.1472051, 0.1471996, 
    0.1472329, 0.1472181, 0.1472598, 0.147248, 0.1471708, 0.1471744, 
    0.1471867, 0.1471808, 0.1471979, 0.1472021, 0.1472056, 0.1472099, 
    0.1472105, 0.147213, 0.1472088, 0.1472129, 0.1471974, 0.1472043, 
    0.1471854, 0.1471899, 0.1471879, 0.1471856, 0.1471927, 0.1472002, 
    0.1472005, 0.1472029, 0.1472093, 0.147198, 0.1472345, 0.1472116, 
    0.1471783, 0.1471849, 0.1471861, 0.1471835, 0.1472017, 0.1471951, 
    0.147213, 0.1472082, 0.1472161, 0.1472122, 0.1472116, 0.1472065, 
    0.1472033, 0.1471953, 0.1471889, 0.1471839, 0.1471851, 0.1471906, 
    0.1472007, 0.1472104, 0.1472083, 0.1472155, 0.1471967, 0.1472045, 
    0.1472014, 0.1472095, 0.147192, 0.1472063, 0.1471884, 0.14719, 0.1471949, 
    0.1472049, 0.1472074, 0.1472097, 0.1472083, 0.147201, 0.1471999, 
    0.1471948, 0.1471934, 0.1471896, 0.1471864, 0.1471893, 0.1471923, 
    0.1472011, 0.1472089, 0.1472176, 0.1472197, 0.1472295, 0.1472214, 
    0.1472346, 0.147223, 0.1472433, 0.1472074, 0.147223, 0.1471952, 
    0.1471982, 0.1472035, 0.147216, 0.1472094, 0.1472172, 0.1471998, 
    0.1471907, 0.1471885, 0.1471842, 0.1471886, 0.1471883, 0.1471925, 
    0.1471912, 0.1472013, 0.1471959, 0.1472115, 0.1472172, 0.1472336, 
    0.1472436, 0.147254, 0.1472586, 0.14726, 0.1472605,
  0.1568999, 0.1569084, 0.1569068, 0.1569135, 0.1569098, 0.1569142, 
    0.1569017, 0.1569086, 0.1569043, 0.1569008, 0.1569265, 0.1569138, 
    0.1569405, 0.1569322, 0.1569534, 0.1569391, 0.1569563, 0.1569531, 
    0.1569631, 0.1569603, 0.1569728, 0.1569644, 0.1569796, 0.1569709, 
    0.1569722, 0.1569641, 0.1569165, 0.1569249, 0.156916, 0.1569172, 
    0.1569167, 0.1569099, 0.1569063, 0.1568994, 0.1569007, 0.1569058, 
    0.1569178, 0.1569138, 0.1569241, 0.1569239, 0.1569353, 0.1569301, 
    0.1569497, 0.1569442, 0.1569604, 0.1569563, 0.1569602, 0.156959, 
    0.1569602, 0.1569541, 0.1569567, 0.1569515, 0.1569311, 0.156937, 
    0.1569194, 0.1569087, 0.156902, 0.1568971, 0.1568978, 0.1568991, 
    0.1569058, 0.1569123, 0.1569173, 0.1569206, 0.1569238, 0.1569334, 
    0.1569388, 0.1569507, 0.1569487, 0.1569523, 0.1569559, 0.1569617, 
    0.1569608, 0.1569633, 0.1569523, 0.1569596, 0.1569475, 0.1569508, 
    0.1569242, 0.1569149, 0.1569105, 0.1569071, 0.1568983, 0.1569043, 
    0.1569019, 0.1569077, 0.1569113, 0.1569096, 0.1569207, 0.1569163, 
    0.1569391, 0.1569293, 0.1569554, 0.1569491, 0.156957, 0.156953, 
    0.1569598, 0.1569537, 0.1569643, 0.1569667, 0.156965, 0.1569713, 
    0.1569533, 0.1569601, 0.1569095, 0.1569098, 0.1569111, 0.1569051, 
    0.1569047, 0.1568993, 0.1569042, 0.1569062, 0.1569116, 0.1569147, 
    0.1569176, 0.1569242, 0.1569315, 0.1569419, 0.1569495, 0.1569546, 
    0.1569515, 0.1569543, 0.1569512, 0.1569498, 0.1569658, 0.1569567, 
    0.1569704, 0.1569697, 0.1569634, 0.1569698, 0.15691, 0.1569083, 
    0.1569024, 0.156907, 0.1568988, 0.1569033, 0.1569059, 0.1569163, 
    0.1569187, 0.1569208, 0.156925, 0.1569304, 0.1569399, 0.1569483, 
    0.1569561, 0.1569555, 0.1569557, 0.1569574, 0.1569532, 0.1569581, 
    0.1569589, 0.1569568, 0.1569696, 0.1569659, 0.1569697, 0.1569673, 
    0.1569089, 0.1569117, 0.1569102, 0.156913, 0.1569109, 0.1569199, 
    0.1569226, 0.1569354, 0.1569303, 0.1569386, 0.1569312, 0.1569325, 
    0.1569387, 0.1569316, 0.1569477, 0.1569366, 0.1569575, 0.156946, 
    0.1569582, 0.156956, 0.1569596, 0.1569628, 0.1569669, 0.1569743, 
    0.1569726, 0.1569789, 0.1569159, 0.1569195, 0.1569193, 0.1569232, 
    0.156926, 0.1569323, 0.1569423, 0.1569386, 0.1569456, 0.156947, 
    0.1569364, 0.1569428, 0.156922, 0.1569252, 0.1569234, 0.1569161, 
    0.1569393, 0.1569273, 0.1569497, 0.1569431, 0.1569623, 0.1569526, 
    0.1569717, 0.1569796, 0.1569876, 0.1569964, 0.1569216, 0.1569191, 
    0.1569237, 0.1569297, 0.1569357, 0.1569435, 0.1569443, 0.1569458, 
    0.1569496, 0.1569528, 0.1569461, 0.1569536, 0.1569258, 0.1569404, 
    0.1569181, 0.1569247, 0.1569294, 0.1569274, 0.1569382, 0.1569407, 
    0.1569509, 0.1569457, 0.1569776, 0.1569633, 0.1570035, 0.1569921, 
    0.1569182, 0.1569216, 0.1569334, 0.1569278, 0.1569441, 0.156948, 
    0.1569514, 0.1569555, 0.156956, 0.1569585, 0.1569545, 0.1569584, 
    0.1569435, 0.1569501, 0.1569321, 0.1569364, 0.1569345, 0.1569323, 
    0.1569391, 0.1569462, 0.1569465, 0.1569488, 0.1569549, 0.1569441, 
    0.1569791, 0.1569571, 0.1569253, 0.1569317, 0.1569328, 0.1569303, 
    0.1569476, 0.1569413, 0.1569584, 0.1569538, 0.1569615, 0.1569577, 
    0.1569571, 0.1569522, 0.1569492, 0.1569416, 0.1569354, 0.1569307, 
    0.1569318, 0.156937, 0.1569467, 0.156956, 0.1569539, 0.1569609, 
    0.1569429, 0.1569503, 0.1569474, 0.1569551, 0.1569384, 0.1569521, 
    0.1569349, 0.1569365, 0.1569412, 0.1569507, 0.1569531, 0.1569553, 
    0.1569539, 0.156947, 0.1569459, 0.1569411, 0.1569397, 0.1569361, 
    0.1569331, 0.1569358, 0.1569387, 0.156947, 0.1569545, 0.1569628, 
    0.1569649, 0.1569743, 0.1569665, 0.1569792, 0.1569681, 0.1569876, 
    0.1569531, 0.1569681, 0.1569415, 0.1569443, 0.1569494, 0.1569613, 
    0.156955, 0.1569625, 0.1569459, 0.1569371, 0.1569351, 0.1569309, 
    0.1569352, 0.1569348, 0.1569389, 0.1569376, 0.1569473, 0.1569421, 
    0.156957, 0.1569625, 0.1569782, 0.1569878, 0.1569979, 0.1570023, 
    0.1570037, 0.1570042,
  0.1704893, 0.1704958, 0.1704945, 0.1704997, 0.1704969, 0.1705003, 
    0.1704907, 0.170496, 0.1704926, 0.17049, 0.1705098, 0.1705, 0.1705206, 
    0.1705142, 0.1705307, 0.1705196, 0.170533, 0.1705305, 0.1705383, 
    0.1705361, 0.170546, 0.1705394, 0.1705514, 0.1705445, 0.1705455, 
    0.1705391, 0.1705021, 0.1705085, 0.1705016, 0.1705026, 0.1705022, 
    0.1704969, 0.1704942, 0.1704889, 0.1704899, 0.1704938, 0.170503, 
    0.1704999, 0.1705079, 0.1705077, 0.1705166, 0.1705126, 0.1705278, 
    0.1705235, 0.1705362, 0.1705329, 0.170536, 0.1705351, 0.170536, 
    0.1705313, 0.1705333, 0.1705292, 0.1705133, 0.1705179, 0.1705042, 
    0.170496, 0.1704909, 0.1704872, 0.1704877, 0.1704887, 0.1704938, 
    0.1704988, 0.1705026, 0.1705052, 0.1705077, 0.1705151, 0.1705193, 
    0.1705286, 0.170527, 0.1705298, 0.1705326, 0.1705372, 0.1705365, 
    0.1705385, 0.1705298, 0.1705355, 0.1705261, 0.1705287, 0.170508, 
    0.1705008, 0.1704974, 0.1704948, 0.1704881, 0.1704927, 0.1704909, 
    0.1704953, 0.170498, 0.1704967, 0.1705052, 0.1705019, 0.1705195, 
    0.1705119, 0.1705323, 0.1705274, 0.1705335, 0.1705304, 0.1705357, 
    0.1705309, 0.1705393, 0.1705411, 0.1705399, 0.1705448, 0.1705306, 
    0.170536, 0.1704966, 0.1704969, 0.1704979, 0.1704932, 0.170493, 
    0.1704889, 0.1704926, 0.1704941, 0.1704982, 0.1705006, 0.1705029, 
    0.170508, 0.1705136, 0.1705217, 0.1705277, 0.1705317, 0.1705292, 
    0.1705314, 0.170529, 0.1705279, 0.1705404, 0.1705333, 0.1705441, 
    0.1705435, 0.1705385, 0.1705436, 0.170497, 0.1704957, 0.1704912, 
    0.1704948, 0.1704884, 0.1704919, 0.1704939, 0.1705019, 0.1705037, 
    0.1705053, 0.1705086, 0.1705128, 0.1705201, 0.1705267, 0.1705328, 
    0.1705324, 0.1705325, 0.1705338, 0.1705305, 0.1705344, 0.170535, 
    0.1705333, 0.1705434, 0.1705406, 0.1705435, 0.1705416, 0.1704962, 
    0.1704983, 0.1704971, 0.1704993, 0.1704978, 0.1705046, 0.1705067, 
    0.1705167, 0.1705127, 0.1705192, 0.1705134, 0.1705144, 0.1705192, 
    0.1705137, 0.1705263, 0.1705176, 0.1705339, 0.1705249, 0.1705344, 
    0.1705328, 0.1705356, 0.1705381, 0.1705413, 0.1705472, 0.1705459, 
    0.1705508, 0.1705016, 0.1705043, 0.1705042, 0.1705071, 0.1705094, 
    0.1705142, 0.170522, 0.1705191, 0.1705246, 0.1705257, 0.1705174, 
    0.1705224, 0.1705063, 0.1705088, 0.1705073, 0.1705018, 0.1705197, 
    0.1705104, 0.1705278, 0.1705226, 0.1705377, 0.1705301, 0.1705451, 
    0.1705514, 0.1705577, 0.1705648, 0.170506, 0.170504, 0.1705075, 
    0.1705122, 0.1705169, 0.1705229, 0.1705236, 0.1705247, 0.1705277, 
    0.1705302, 0.170525, 0.1705309, 0.1705092, 0.1705205, 0.1705033, 
    0.1705083, 0.170512, 0.1705105, 0.1705188, 0.1705208, 0.1705288, 
    0.1705247, 0.1705498, 0.1705385, 0.1705704, 0.1705613, 0.1705034, 
    0.170506, 0.1705151, 0.1705107, 0.1705234, 0.1705265, 0.1705291, 
    0.1705323, 0.1705328, 0.1705347, 0.1705315, 0.1705346, 0.170523, 
    0.1705281, 0.1705141, 0.1705174, 0.1705159, 0.1705142, 0.1705195, 
    0.1705251, 0.1705253, 0.1705271, 0.1705319, 0.1705234, 0.170551, 
    0.1705336, 0.1705088, 0.1705138, 0.1705146, 0.1705127, 0.1705262, 
    0.1705212, 0.1705347, 0.170531, 0.170537, 0.170534, 0.1705336, 0.1705298, 
    0.1705274, 0.1705215, 0.1705167, 0.170513, 0.1705139, 0.1705179, 
    0.1705254, 0.1705327, 0.1705311, 0.1705366, 0.1705225, 0.1705283, 
    0.170526, 0.170532, 0.170519, 0.1705297, 0.1705163, 0.1705175, 0.1705212, 
    0.1705286, 0.1705304, 0.1705322, 0.1705311, 0.1705257, 0.1705248, 
    0.1705211, 0.17052, 0.1705172, 0.1705149, 0.170517, 0.1705192, 0.1705257, 
    0.1705316, 0.1705381, 0.1705398, 0.1705472, 0.170541, 0.1705511, 
    0.1705423, 0.1705577, 0.1705305, 0.1705422, 0.1705214, 0.1705236, 
    0.1705275, 0.1705369, 0.170532, 0.1705378, 0.1705248, 0.170518, 
    0.1705164, 0.1705132, 0.1705165, 0.1705162, 0.1705194, 0.1705184, 
    0.1705259, 0.1705219, 0.1705335, 0.1705378, 0.1705503, 0.1705579, 
    0.170566, 0.1705695, 0.1705706, 0.170571,
  0.1855468, 0.18555, 0.1855494, 0.185552, 0.1855506, 0.1855523, 0.1855475, 
    0.1855502, 0.1855485, 0.1855471, 0.1855572, 0.1855522, 0.1855628, 
    0.1855594, 0.185568, 0.1855622, 0.1855693, 0.185568, 0.1855721, 
    0.1855709, 0.1855762, 0.1855727, 0.1855791, 0.1855754, 0.1855759, 
    0.1855725, 0.1855532, 0.1855565, 0.185553, 0.1855535, 0.1855533, 
    0.1855506, 0.1855492, 0.1855466, 0.1855471, 0.1855491, 0.1855537, 
    0.1855522, 0.1855562, 0.1855561, 0.1855607, 0.1855586, 0.1855665, 
    0.1855643, 0.185571, 0.1855692, 0.1855709, 0.1855704, 0.1855709, 
    0.1855684, 0.1855694, 0.1855673, 0.185559, 0.1855613, 0.1855543, 
    0.1855502, 0.1855476, 0.1855458, 0.185546, 0.1855465, 0.1855491, 
    0.1855516, 0.1855535, 0.1855548, 0.1855561, 0.1855599, 0.1855621, 
    0.185567, 0.1855661, 0.1855676, 0.1855691, 0.1855715, 0.1855711, 
    0.1855722, 0.1855676, 0.1855706, 0.1855656, 0.185567, 0.1855562, 
    0.1855526, 0.1855509, 0.1855495, 0.1855462, 0.1855485, 0.1855476, 
    0.1855498, 0.1855512, 0.1855505, 0.1855548, 0.1855531, 0.1855622, 
    0.1855582, 0.1855689, 0.1855663, 0.1855695, 0.1855679, 0.1855707, 
    0.1855682, 0.1855726, 0.1855736, 0.1855729, 0.1855756, 0.185568, 
    0.1855709, 0.1855505, 0.1855506, 0.1855511, 0.1855488, 0.1855486, 
    0.1855466, 0.1855484, 0.1855492, 0.1855513, 0.1855525, 0.1855537, 
    0.1855562, 0.1855592, 0.1855633, 0.1855665, 0.1855686, 0.1855673, 
    0.1855684, 0.1855672, 0.1855666, 0.1855732, 0.1855694, 0.1855752, 
    0.1855749, 0.1855722, 0.1855749, 0.1855507, 0.18555, 0.1855478, 
    0.1855495, 0.1855464, 0.1855481, 0.1855491, 0.1855531, 0.1855541, 
    0.1855549, 0.1855566, 0.1855587, 0.1855625, 0.1855659, 0.1855692, 
    0.1855689, 0.185569, 0.1855697, 0.185568, 0.18557, 0.1855703, 0.1855695, 
    0.1855748, 0.1855733, 0.1855749, 0.1855739, 0.1855502, 0.1855513, 
    0.1855507, 0.1855518, 0.185551, 0.1855545, 0.1855556, 0.1855607, 
    0.1855587, 0.185562, 0.185559, 0.1855595, 0.185562, 0.1855592, 0.1855657, 
    0.1855612, 0.1855697, 0.185565, 0.18557, 0.1855692, 0.1855706, 0.185572, 
    0.1855737, 0.1855769, 0.1855761, 0.1855788, 0.185553, 0.1855544, 
    0.1855543, 0.1855558, 0.1855569, 0.1855595, 0.1855635, 0.185562, 
    0.1855648, 0.1855654, 0.1855611, 0.1855637, 0.1855554, 0.1855567, 
    0.1855559, 0.1855531, 0.1855623, 0.1855575, 0.1855665, 0.1855638, 
    0.1855718, 0.1855678, 0.1855757, 0.1855791, 0.1855825, 0.1855864, 
    0.1855552, 0.1855543, 0.185556, 0.1855584, 0.1855608, 0.185564, 
    0.1855643, 0.1855649, 0.1855665, 0.1855678, 0.1855651, 0.1855682, 
    0.1855569, 0.1855627, 0.1855538, 0.1855564, 0.1855583, 0.1855575, 
    0.1855618, 0.1855628, 0.185567, 0.1855649, 0.1855782, 0.1855722, 
    0.1855895, 0.1855845, 0.1855539, 0.1855552, 0.1855599, 0.1855577, 
    0.1855642, 0.1855659, 0.1855672, 0.1855689, 0.1855692, 0.1855702, 
    0.1855685, 0.1855701, 0.185564, 0.1855667, 0.1855594, 0.1855611, 
    0.1855603, 0.1855595, 0.1855622, 0.1855651, 0.1855652, 0.1855662, 
    0.1855687, 0.1855642, 0.1855789, 0.1855696, 0.1855567, 0.1855592, 
    0.1855597, 0.1855587, 0.1855657, 0.1855631, 0.1855702, 0.1855682, 
    0.1855714, 0.1855698, 0.1855696, 0.1855676, 0.1855663, 0.1855632, 
    0.1855607, 0.1855588, 0.1855593, 0.1855614, 0.1855653, 0.1855691, 
    0.1855683, 0.1855712, 0.1855637, 0.1855668, 0.1855656, 0.1855687, 
    0.1855619, 0.1855675, 0.1855605, 0.1855611, 0.1855631, 0.1855669, 
    0.1855679, 0.1855688, 0.1855683, 0.1855654, 0.185565, 0.185563, 
    0.1855624, 0.185561, 0.1855598, 0.1855609, 0.185562, 0.1855654, 
    0.1855685, 0.185572, 0.1855729, 0.1855768, 0.1855735, 0.1855789, 
    0.1855742, 0.1855825, 0.185568, 0.1855742, 0.1855632, 0.1855643, 
    0.1855664, 0.1855714, 0.1855687, 0.1855718, 0.185565, 0.1855614, 
    0.1855606, 0.1855589, 0.1855606, 0.1855605, 0.1855621, 0.1855616, 
    0.1855656, 0.1855634, 0.1855696, 0.1855718, 0.1855785, 0.1855827, 
    0.185587, 0.185589, 0.1855896, 0.1855898,
  0.1955522, 0.1955529, 0.1955528, 0.1955534, 0.195553, 0.1955535, 0.1955523, 
    0.1955529, 0.1955525, 0.1955522, 0.1955546, 0.1955534, 0.195556, 
    0.1955552, 0.1955574, 0.1955559, 0.1955577, 0.1955574, 0.1955585, 
    0.1955581, 0.1955596, 0.1955586, 0.1955603, 0.1955594, 0.1955595, 
    0.1955586, 0.1955537, 0.1955545, 0.1955536, 0.1955537, 0.1955537, 
    0.195553, 0.1955527, 0.1955521, 0.1955522, 0.1955527, 0.1955538, 
    0.1955534, 0.1955544, 0.1955544, 0.1955555, 0.195555, 0.195557, 
    0.1955564, 0.1955582, 0.1955577, 0.1955581, 0.195558, 0.1955581, 
    0.1955575, 0.1955578, 0.1955572, 0.1955551, 0.1955557, 0.1955539, 
    0.1955529, 0.1955523, 0.1955519, 0.195552, 0.1955521, 0.1955527, 
    0.1955533, 0.1955537, 0.1955541, 0.1955544, 0.1955553, 0.1955559, 
    0.1955571, 0.1955569, 0.1955573, 0.1955577, 0.1955583, 0.1955582, 
    0.1955585, 0.1955573, 0.1955581, 0.1955568, 0.1955571, 0.1955544, 
    0.1955535, 0.1955531, 0.1955528, 0.195552, 0.1955525, 0.1955523, 
    0.1955529, 0.1955532, 0.195553, 0.1955541, 0.1955537, 0.1955559, 
    0.1955549, 0.1955576, 0.195557, 0.1955578, 0.1955574, 0.1955581, 
    0.1955574, 0.1955586, 0.1955589, 0.1955587, 0.1955594, 0.1955574, 
    0.1955581, 0.195553, 0.195553, 0.1955532, 0.1955526, 0.1955526, 
    0.1955521, 0.1955525, 0.1955527, 0.1955532, 0.1955535, 0.1955538, 
    0.1955544, 0.1955551, 0.1955562, 0.195557, 0.1955575, 0.1955572, 
    0.1955575, 0.1955572, 0.195557, 0.1955588, 0.1955578, 0.1955593, 
    0.1955592, 0.1955585, 0.1955592, 0.1955531, 0.1955529, 0.1955524, 
    0.1955528, 0.1955521, 0.1955525, 0.1955527, 0.1955536, 0.1955539, 
    0.1955541, 0.1955545, 0.195555, 0.195556, 0.1955569, 0.1955577, 
    0.1955576, 0.1955577, 0.1955578, 0.1955574, 0.1955579, 0.195558, 
    0.1955578, 0.1955592, 0.1955588, 0.1955592, 0.1955589, 0.195553, 
    0.1955532, 0.1955531, 0.1955533, 0.1955532, 0.195554, 0.1955543, 
    0.1955555, 0.195555, 0.1955559, 0.1955551, 0.1955552, 0.1955559, 
    0.1955551, 0.1955568, 0.1955556, 0.1955578, 0.1955566, 0.1955579, 
    0.1955577, 0.1955581, 0.1955584, 0.1955589, 0.1955597, 0.1955595, 
    0.1955603, 0.1955536, 0.195554, 0.1955539, 0.1955543, 0.1955546, 
    0.1955552, 0.1955562, 0.1955559, 0.1955566, 0.1955567, 0.1955556, 
    0.1955563, 0.1955542, 0.1955545, 0.1955543, 0.1955536, 0.1955559, 
    0.1955547, 0.195557, 0.1955563, 0.1955584, 0.1955573, 0.1955594, 
    0.1955604, 0.1955613, 0.1955623, 0.1955542, 0.1955539, 0.1955544, 
    0.195555, 0.1955556, 0.1955564, 0.1955564, 0.1955566, 0.195557, 
    0.1955573, 0.1955566, 0.1955574, 0.1955546, 0.195556, 0.1955538, 
    0.1955545, 0.1955549, 0.1955547, 0.1955558, 0.1955561, 0.1955571, 
    0.1955566, 0.1955601, 0.1955585, 0.1955632, 0.1955618, 0.1955538, 
    0.1955542, 0.1955553, 0.1955548, 0.1955564, 0.1955568, 0.1955572, 
    0.1955576, 0.1955577, 0.195558, 0.1955575, 0.1955579, 0.1955564, 
    0.1955571, 0.1955552, 0.1955556, 0.1955554, 0.1955552, 0.1955559, 
    0.1955566, 0.1955567, 0.1955569, 0.1955576, 0.1955564, 0.1955603, 
    0.1955578, 0.1955545, 0.1955552, 0.1955553, 0.195555, 0.1955568, 
    0.1955561, 0.195558, 0.1955574, 0.1955583, 0.1955579, 0.1955578, 
    0.1955573, 0.195557, 0.1955561, 0.1955555, 0.195555, 0.1955552, 
    0.1955557, 0.1955567, 0.1955577, 0.1955575, 0.1955582, 0.1955563, 
    0.1955571, 0.1955568, 0.1955576, 0.1955558, 0.1955573, 0.1955555, 
    0.1955556, 0.1955561, 0.1955571, 0.1955574, 0.1955576, 0.1955575, 
    0.1955567, 0.1955566, 0.1955561, 0.195556, 0.1955556, 0.1955553, 
    0.1955556, 0.1955559, 0.1955567, 0.1955575, 0.1955584, 0.1955587, 
    0.1955597, 0.1955588, 0.1955603, 0.195559, 0.1955613, 0.1955574, 
    0.195559, 0.1955561, 0.1955564, 0.195557, 0.1955583, 0.1955576, 
    0.1955584, 0.1955566, 0.1955557, 0.1955555, 0.1955551, 0.1955555, 
    0.1955555, 0.1955559, 0.1955557, 0.1955568, 0.1955562, 0.1955578, 
    0.1955584, 0.1955602, 0.1955613, 0.1955625, 0.1955631, 0.1955632, 
    0.1955633,
  0.1982741, 0.1982741, 0.1982741, 0.1982742, 0.1982742, 0.1982742, 
    0.1982741, 0.1982742, 0.1982741, 0.1982741, 0.1982743, 0.1982742, 
    0.1982745, 0.1982744, 0.1982747, 0.1982745, 0.1982747, 0.1982747, 
    0.1982748, 0.1982748, 0.198275, 0.1982748, 0.1982751, 0.1982749, 
    0.1982749, 0.1982748, 0.1982742, 0.1982743, 0.1982742, 0.1982742, 
    0.1982742, 0.1982742, 0.1982741, 0.198274, 0.1982741, 0.1982741, 
    0.1982742, 0.1982742, 0.1982743, 0.1982743, 0.1982744, 0.1982744, 
    0.1982746, 0.1982746, 0.1982748, 0.1982747, 0.1982748, 0.1982748, 
    0.1982748, 0.1982747, 0.1982747, 0.1982747, 0.1982744, 0.1982745, 
    0.1982743, 0.1982742, 0.1982741, 0.198274, 0.198274, 0.198274, 0.1982741, 
    0.1982742, 0.1982742, 0.1982743, 0.1982743, 0.1982744, 0.1982745, 
    0.1982746, 0.1982746, 0.1982747, 0.1982747, 0.1982748, 0.1982748, 
    0.1982748, 0.1982747, 0.1982748, 0.1982746, 0.1982746, 0.1982743, 
    0.1982742, 0.1982742, 0.1982741, 0.198274, 0.1982741, 0.1982741, 
    0.1982741, 0.1982742, 0.1982742, 0.1982743, 0.1982742, 0.1982745, 
    0.1982744, 0.1982747, 0.1982746, 0.1982747, 0.1982747, 0.1982748, 
    0.1982747, 0.1982748, 0.1982749, 0.1982748, 0.1982749, 0.1982747, 
    0.1982748, 0.1982742, 0.1982742, 0.1982742, 0.1982741, 0.1982741, 
    0.198274, 0.1982741, 0.1982741, 0.1982742, 0.1982742, 0.1982742, 
    0.1982743, 0.1982744, 0.1982745, 0.1982746, 0.1982747, 0.1982747, 
    0.1982747, 0.1982746, 0.1982746, 0.1982749, 0.1982747, 0.1982749, 
    0.1982749, 0.1982748, 0.1982749, 0.1982742, 0.1982741, 0.1982741, 
    0.1982741, 0.198274, 0.1982741, 0.1982741, 0.1982742, 0.1982743, 
    0.1982743, 0.1982743, 0.1982744, 0.1982745, 0.1982746, 0.1982747, 
    0.1982747, 0.1982747, 0.1982747, 0.1982747, 0.1982747, 0.1982748, 
    0.1982747, 0.1982749, 0.1982749, 0.1982749, 0.1982749, 0.1982742, 
    0.1982742, 0.1982742, 0.1982742, 0.1982742, 0.1982743, 0.1982743, 
    0.1982744, 0.1982744, 0.1982745, 0.1982744, 0.1982744, 0.1982745, 
    0.1982744, 0.1982746, 0.1982745, 0.1982747, 0.1982746, 0.1982747, 
    0.1982747, 0.1982748, 0.1982748, 0.1982749, 0.198275, 0.198275, 0.198275, 
    0.1982742, 0.1982743, 0.1982743, 0.1982743, 0.1982743, 0.1982744, 
    0.1982745, 0.1982745, 0.1982746, 0.1982746, 0.1982745, 0.1982745, 
    0.1982743, 0.1982743, 0.1982743, 0.1982742, 0.1982745, 0.1982743, 
    0.1982746, 0.1982745, 0.1982748, 0.1982747, 0.1982749, 0.1982751, 
    0.1982752, 0.1982753, 0.1982743, 0.1982743, 0.1982743, 0.1982744, 
    0.1982744, 0.1982746, 0.1982746, 0.1982746, 0.1982746, 0.1982747, 
    0.1982746, 0.1982747, 0.1982743, 0.1982745, 0.1982742, 0.1982743, 
    0.1982744, 0.1982743, 0.1982745, 0.1982745, 0.1982746, 0.1982746, 
    0.198275, 0.1982748, 0.1982754, 0.1982753, 0.1982742, 0.1982743, 
    0.1982744, 0.1982744, 0.1982746, 0.1982746, 0.1982747, 0.1982747, 
    0.1982747, 0.1982747, 0.1982747, 0.1982747, 0.1982746, 0.1982746, 
    0.1982744, 0.1982745, 0.1982744, 0.1982744, 0.1982745, 0.1982746, 
    0.1982746, 0.1982746, 0.1982747, 0.1982746, 0.198275, 0.1982747, 
    0.1982743, 0.1982744, 0.1982744, 0.1982744, 0.1982746, 0.1982745, 
    0.1982747, 0.1982747, 0.1982748, 0.1982747, 0.1982747, 0.1982747, 
    0.1982746, 0.1982745, 0.1982744, 0.1982744, 0.1982744, 0.1982745, 
    0.1982746, 0.1982747, 0.1982747, 0.1982748, 0.1982745, 0.1982746, 
    0.1982746, 0.1982747, 0.1982745, 0.1982747, 0.1982744, 0.1982745, 
    0.1982745, 0.1982746, 0.1982747, 0.1982747, 0.1982747, 0.1982746, 
    0.1982746, 0.1982745, 0.1982745, 0.1982745, 0.1982744, 0.1982744, 
    0.1982745, 0.1982746, 0.1982747, 0.1982748, 0.1982748, 0.198275, 
    0.1982749, 0.1982751, 0.1982749, 0.1982752, 0.1982747, 0.1982749, 
    0.1982745, 0.1982746, 0.1982746, 0.1982748, 0.1982747, 0.1982748, 
    0.1982746, 0.1982745, 0.1982744, 0.1982744, 0.1982744, 0.1982744, 
    0.1982745, 0.1982745, 0.1982746, 0.1982745, 0.1982747, 0.1982748, 
    0.198275, 0.1982752, 0.1982753, 0.1982754, 0.1982754, 0.1982755,
  0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985156, 0.1985156, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985156, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985156, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985158, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 
    0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985157, 0.1985158, 
    0.1985158, 0.1985158,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  8.606007, 8.606067, 8.606055, 8.606104, 8.606077, 8.606109, 8.606019, 
    8.606069, 8.606037, 8.606012, 8.606196, 8.606106, 8.606295, 8.606236, 
    8.606385, 8.606285, 8.606406, 8.606383, 8.606454, 8.606434, 8.606569, 
    8.606463, 8.606642, 8.606548, 8.606563, 8.606461, 8.606126, 8.606185, 
    8.606122, 8.606131, 8.606127, 8.606078, 8.606052, 8.606003, 8.606011, 
    8.606049, 8.606134, 8.606106, 8.606179, 8.606177, 8.606258, 8.606222, 
    8.606359, 8.60632, 8.606435, 8.606405, 8.606433, 8.606425, 8.606433, 
    8.606391, 8.606409, 8.606372, 8.606229, 8.606271, 8.606146, 8.606069, 
    8.606021, 8.605986, 8.605991, 8.606, 8.606049, 8.606095, 8.606131, 
    8.606154, 8.606177, 8.606245, 8.606283, 8.606366, 8.606353, 8.606377, 
    8.606402, 8.606444, 8.606438, 8.606455, 8.606378, 8.606429, 8.606344, 
    8.606367, 8.606179, 8.606113, 8.606082, 8.606058, 8.605994, 8.606038, 
    8.606021, 8.606063, 8.606089, 8.606075, 8.606155, 8.606124, 8.606285, 
    8.606215, 8.6064, 8.606356, 8.606411, 8.606382, 8.60643, 8.606387, 
    8.606462, 8.606495, 8.606467, 8.606552, 8.606384, 8.606433, 8.606075, 
    8.606077, 8.606087, 8.606043, 8.606041, 8.606002, 8.606037, 8.606051, 
    8.606091, 8.606112, 8.606133, 8.60618, 8.606232, 8.606305, 8.606359, 
    8.606394, 8.606372, 8.606392, 8.60637, 8.60636, 8.606481, 8.606409, 
    8.606542, 8.606533, 8.606456, 8.606534, 8.606079, 8.606067, 8.606025, 
    8.606058, 8.605998, 8.60603, 8.60605, 8.606124, 8.606141, 8.606155, 
    8.606186, 8.606224, 8.606291, 8.606349, 8.606404, 8.6064, 8.606401, 
    8.606414, 8.606383, 8.606419, 8.606424, 8.606409, 8.606532, 8.606483, 
    8.606533, 8.606503, 8.606071, 8.606091, 8.60608, 8.6061, 8.606086, 
    8.60615, 8.606169, 8.606259, 8.606223, 8.606282, 8.60623, 8.606238, 
    8.606282, 8.606233, 8.606345, 8.606267, 8.606414, 8.606334, 8.60642, 
    8.606404, 8.606429, 8.606451, 8.606499, 8.606586, 8.606567, 8.606635, 
    8.606121, 8.606147, 8.606145, 8.606173, 8.606193, 8.606237, 8.606308, 
    8.606281, 8.606331, 8.60634, 8.606266, 8.606311, 8.606165, 8.606187, 
    8.606174, 8.606123, 8.606286, 8.606202, 8.606359, 8.606313, 8.606448, 
    8.60638, 8.606557, 8.606642, 8.606722, 8.606807, 8.606162, 8.606144, 
    8.606176, 8.606219, 8.606261, 8.606316, 8.606322, 8.606332, 8.606359, 
    8.606381, 8.606335, 8.606387, 8.606191, 8.606295, 8.606136, 8.606183, 
    8.606216, 8.606203, 8.606278, 8.606297, 8.606368, 8.606331, 8.606621, 
    8.606455, 8.606873, 8.606766, 8.606138, 8.606162, 8.606245, 8.606206, 
    8.60632, 8.606348, 8.606371, 8.6064, 8.606404, 8.606421, 8.606393, 
    8.606421, 8.606316, 8.606362, 8.606236, 8.606266, 8.606253, 8.606237, 
    8.606285, 8.606335, 8.606338, 8.606353, 8.606396, 8.60632, 8.606636, 
    8.606411, 8.606188, 8.606233, 8.606241, 8.606223, 8.606345, 8.6063, 
    8.606421, 8.606388, 8.606442, 8.606416, 8.606411, 8.606377, 8.606356, 
    8.606302, 8.606259, 8.606226, 8.606234, 8.606271, 8.606339, 8.606403, 
    8.606389, 8.606438, 8.606312, 8.606363, 8.606343, 8.606397, 8.60628, 
    8.606376, 8.606256, 8.606267, 8.606299, 8.606366, 8.606382, 8.606399, 
    8.606389, 8.60634, 8.606333, 8.606299, 8.60629, 8.606264, 8.606243, 
    8.606262, 8.606282, 8.60634, 8.606393, 8.606452, 8.606466, 8.606586, 
    8.606492, 8.606637, 8.606513, 8.606722, 8.606383, 8.606513, 8.606301, 
    8.606322, 8.606357, 8.606441, 8.606397, 8.606449, 8.606333, 8.606271, 
    8.606257, 8.606228, 8.606257, 8.606256, 8.606284, 8.606275, 8.606342, 
    8.606306, 8.606411, 8.606449, 8.606627, 8.606724, 8.606821, 8.606862, 
    8.606874, 8.606879 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  3.991914e-15, 3.992308e-15, 3.992233e-15, 3.992547e-15, 3.992375e-15, 
    3.992579e-15, 3.991997e-15, 3.99232e-15, 3.992116e-15, 3.991954e-15, 
    3.993147e-15, 3.992561e-15, 3.993789e-15, 3.993409e-15, 3.994376e-15, 
    3.993725e-15, 3.994509e-15, 3.994365e-15, 3.994817e-15, 3.994688e-15, 
    3.99525e-15, 3.994877e-15, 3.995556e-15, 3.995165e-15, 3.995223e-15, 
    3.994863e-15, 3.992686e-15, 3.993071e-15, 3.992662e-15, 3.992717e-15, 
    3.992694e-15, 3.992376e-15, 3.992211e-15, 3.991889e-15, 3.991949e-15, 
    3.992188e-15, 3.992742e-15, 3.992559e-15, 3.993036e-15, 3.993026e-15, 
    3.993552e-15, 3.993314e-15, 3.994208e-15, 3.993956e-15, 3.994693e-15, 
    3.994507e-15, 3.994683e-15, 3.994631e-15, 3.994684e-15, 3.99441e-15, 
    3.994527e-15, 3.994288e-15, 3.993358e-15, 3.993628e-15, 3.992818e-15, 
    3.99232e-15, 3.99201e-15, 3.991784e-15, 3.991816e-15, 3.991875e-15, 
    3.99219e-15, 3.992492e-15, 3.992721e-15, 3.992873e-15, 3.993024e-15, 
    3.993461e-15, 3.99371e-15, 3.994255e-15, 3.994164e-15, 3.994324e-15, 
    3.994488e-15, 3.994754e-15, 3.994711e-15, 3.994827e-15, 3.994325e-15, 
    3.994656e-15, 3.99411e-15, 3.994258e-15, 3.993038e-15, 3.99261e-15, 
    3.992405e-15, 3.992246e-15, 3.99184e-15, 3.992119e-15, 3.992008e-15, 
    3.992277e-15, 3.992444e-15, 3.992363e-15, 3.992877e-15, 3.992676e-15, 
    3.993724e-15, 3.993272e-15, 3.994469e-15, 3.994183e-15, 3.994539e-15, 
    3.994358e-15, 3.994665e-15, 3.994389e-15, 3.994872e-15, 3.994973e-15, 
    3.994904e-15, 3.995183e-15, 3.994373e-15, 3.994681e-15, 3.992359e-15, 
    3.992372e-15, 3.992437e-15, 3.992154e-15, 3.992137e-15, 3.991886e-15, 
    3.992112e-15, 3.992206e-15, 3.992456e-15, 3.992599e-15, 3.992737e-15, 
    3.993041e-15, 3.993376e-15, 3.993853e-15, 3.994201e-15, 3.994434e-15, 
    3.994293e-15, 3.994417e-15, 3.994277e-15, 3.994213e-15, 3.994933e-15, 
    3.994526e-15, 3.995142e-15, 3.995109e-15, 3.994828e-15, 3.995113e-15, 
    3.992382e-15, 3.992306e-15, 3.992032e-15, 3.992246e-15, 3.991859e-15, 
    3.992072e-15, 3.992193e-15, 3.992674e-15, 3.992787e-15, 3.992882e-15, 
    3.993078e-15, 3.993326e-15, 3.993761e-15, 3.994144e-15, 3.994499e-15, 
    3.994474e-15, 3.994482e-15, 3.994559e-15, 3.994366e-15, 3.99459e-15, 
    3.994626e-15, 3.99453e-15, 3.995105e-15, 3.99494e-15, 3.995108e-15, 
    3.995002e-15, 3.992331e-15, 3.992461e-15, 3.992391e-15, 3.992522e-15, 
    3.992427e-15, 3.992841e-15, 3.992965e-15, 3.993556e-15, 3.99332e-15, 
    3.993703e-15, 3.993361e-15, 3.99342e-15, 3.993704e-15, 3.993381e-15, 
    3.994118e-15, 3.993608e-15, 3.994562e-15, 3.99404e-15, 3.994594e-15, 
    3.994497e-15, 3.994659e-15, 3.994802e-15, 3.994986e-15, 3.995319e-15, 
    3.995243e-15, 3.995527e-15, 3.992658e-15, 3.992824e-15, 3.992815e-15, 
    3.992993e-15, 3.993123e-15, 3.993413e-15, 3.993873e-15, 3.993701e-15, 
    3.994021e-15, 3.994084e-15, 3.9936e-15, 3.993892e-15, 3.99294e-15, 
    3.993088e-15, 3.993003e-15, 3.992668e-15, 3.993734e-15, 3.993183e-15, 
    3.994206e-15, 3.993908e-15, 3.994781e-15, 3.994341e-15, 3.9952e-15, 
    3.995556e-15, 3.995915e-15, 3.996309e-15, 3.992921e-15, 3.992807e-15, 
    3.993015e-15, 3.993294e-15, 3.993568e-15, 3.993925e-15, 3.993964e-15, 
    3.99403e-15, 3.994205e-15, 3.994351e-15, 3.994045e-15, 3.994388e-15, 
    3.993112e-15, 3.993784e-15, 3.992759e-15, 3.99306e-15, 3.99328e-15, 
    3.993189e-15, 3.993683e-15, 3.993798e-15, 3.994263e-15, 3.994025e-15, 
    3.995464e-15, 3.994825e-15, 3.996625e-15, 3.996117e-15, 3.992766e-15, 
    3.992923e-15, 3.993462e-15, 3.993206e-15, 3.993951e-15, 3.994133e-15, 
    3.994286e-15, 3.994472e-15, 3.994496e-15, 3.994608e-15, 3.994425e-15, 
    3.994602e-15, 3.993926e-15, 3.994228e-15, 3.993406e-15, 3.993603e-15, 
    3.993514e-15, 3.993413e-15, 3.993725e-15, 3.994049e-15, 3.994064e-15, 
    3.994167e-15, 3.994443e-15, 3.993955e-15, 3.995531e-15, 3.994542e-15, 
    3.993093e-15, 3.993385e-15, 3.993436e-15, 3.993321e-15, 3.994115e-15, 
    3.993826e-15, 3.994606e-15, 3.994396e-15, 3.994742e-15, 3.99457e-15, 
    3.994544e-15, 3.994324e-15, 3.994186e-15, 3.993837e-15, 3.993557e-15, 
    3.993339e-15, 3.99339e-15, 3.99363e-15, 3.994071e-15, 3.994495e-15, 
    3.994401e-15, 3.994716e-15, 3.993897e-15, 3.994236e-15, 3.994102e-15, 
    3.994452e-15, 3.993695e-15, 3.994315e-15, 3.993534e-15, 3.993604e-15, 
    3.99382e-15, 3.994253e-15, 3.994361e-15, 3.994462e-15, 3.994402e-15, 
    3.994083e-15, 3.994035e-15, 3.993817e-15, 3.993753e-15, 3.993589e-15, 
    3.99345e-15, 3.993575e-15, 3.993705e-15, 3.994087e-15, 3.994428e-15, 
    3.994803e-15, 3.994898e-15, 3.995317e-15, 3.994964e-15, 3.995535e-15, 
    3.995033e-15, 3.995912e-15, 3.994363e-15, 3.995034e-15, 3.993833e-15, 
    3.993964e-15, 3.994192e-15, 3.994736e-15, 3.994451e-15, 3.994788e-15, 
    3.994034e-15, 3.993634e-15, 3.993541e-15, 3.993351e-15, 3.993546e-15, 
    3.99353e-15, 3.993716e-15, 3.993657e-15, 3.9941e-15, 3.993862e-15, 
    3.994541e-15, 3.994787e-15, 3.995494e-15, 3.995925e-15, 3.996376e-15, 
    3.996572e-15, 3.996633e-15, 3.996658e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  9.819985, 9.86739, 9.858161, 9.896481, 9.87521, 9.900319, 9.829581, 
    9.869278, 9.843923, 9.824243, 9.971111, 9.89819, 10.0463, 10.00027, 
    10.11615, 10.03914, 10.13172, 10.11391, 10.16754, 10.15216, 10.22492, 
    10.17464, 10.2607, 10.21384, 10.22117, 10.17312, 9.912832, 9.962018, 
    9.909925, 9.916927, 9.913783, 9.875651, 9.856475, 9.816362, 9.823636, 
    9.853098, 9.920077, 9.897305, 9.954742, 9.953444, 10.01721, 9.988657, 
    10.09527, 10.06491, 10.1528, 10.13065, 10.15176, 10.14536, 10.15184, 
    10.11938, 10.13328, 10.10474, 9.994028, 10.02649, 9.928924, 9.870217, 
    9.831322, 9.803784, 9.807674, 9.815094, 9.853271, 9.889239, 9.916707, 
    9.935107, 9.953257, 10.00807, 10.03683, 10.10143, 10.08974, 10.10953, 
    10.12845, 10.16027, 10.15503, 10.16907, 10.10901, 10.1489, 10.08309, 
    10.10107, 9.958221, 9.903443, 9.880239, 9.859936, 9.810666, 9.844676, 
    9.831262, 9.863189, 9.883512, 9.873457, 9.935611, 9.91142, 10.03854, 
    9.984083, 10.12624, 10.09214, 10.13443, 10.11283, 10.14985, 10.11653, 
    10.17429, 10.19084, 10.17828, 10.21535, 10.11469, 10.15176, 9.873177, 
    9.874816, 9.882455, 9.848905, 9.846853, 9.816165, 9.843466, 9.855108, 
    9.884689, 9.902218, 9.918896, 9.955625, 9.996654, 10.05344, 10.09435, 
    10.12183, 10.10497, 10.11985, 10.10322, 10.09543, 10.18611, 10.13341, 
    10.21058, 10.20652, 10.1694, 10.20698, 9.875967, 9.866533, 9.83383, 
    9.859418, 9.812826, 9.838892, 9.853902, 9.911931, 9.924702, 9.936561, 
    9.960003, 9.990139, 10.04234, 10.08788, 10.12955, 10.12649, 10.12757, 
    10.1369, 10.11381, 10.14069, 10.14521, 10.1334, 10.20598, 10.18633, 
    10.20643, 10.19364, 9.869598, 9.885477, 9.876896, 9.893039, 9.881666, 
    9.932302, 9.947515, 10.01845, 9.989547, 10.03555, 9.994226, 10.00154, 
    10.03706, 9.996455, 10.08537, 10.02505, 10.13726, 10.07685, 10.14105, 
    10.12937, 10.14872, 10.16606, 10.19185, 10.23226, 10.22289, 10.25673, 
    9.909176, 9.929827, 9.928003, 9.949636, 9.965655, 10.00027, 10.05534, 
    10.03461, 10.07268, 10.08033, 10.0225, 10.05799, 9.943659, 9.962251, 
    9.951175, 9.910807, 10.03939, 9.973646, 10.09503, 10.0594, 10.16359, 
    10.1117, 10.21774, 10.2616, 10.30296, 10.35144, 9.941103, 9.927059, 
    9.952209, 9.98708, 10.01904, 10.06157, 10.06592, 10.07391, 10.09459, 
    10.11201, 10.07644, 10.11638, 9.966576, 10.04508, 9.921758, 9.959057, 
    9.98502, 9.97362, 10.03224, 10.04603, 10.10217, 10.07312, 10.25077, 
    10.16973, 10.38842, 10.32815, 9.922156, 9.941052, 10.00675, 9.975586, 
    10.06441, 10.08629, 10.1041, 10.12689, 10.12935, 10.14288, 10.12072, 
    10.142, 10.06166, 10.09751, 9.999304, 10.02316, 10.01218, 10.00015, 
    10.03731, 10.077, 10.07784, 10.09059, 10.12658, 10.06477, 10.26076, 
    10.13796, 9.961683, 9.998084, 10.00322, 9.989254, 10.0841, 10.04968, 
    10.14255, 10.11739, 10.15862, 10.13812, 10.13511, 10.10882, 10.09248, 
    10.05126, 10.01779, 9.991296, 9.997452, 10.02657, 10.07943, 10.12958, 
    10.11858, 10.15549, 10.05797, 10.0988, 10.08301, 10.1242, 10.03406, 
    10.11082, 10.0145, 10.02292, 10.049, 10.10157, 10.11322, 10.12567, 
    10.11798, 10.08077, 10.07468, 10.04836, 10.04111, 10.02109, 10.00453, 
    10.01966, 10.03556, 10.08078, 10.12165, 10.16631, 10.17725, 10.23362, 
    10.19094, 10.26143, 10.2015, 10.30536, 10.11526, 10.19973, 10.05018, 
    10.0658, 10.09411, 10.15918, 10.12401, 10.16515, 10.07444, 10.02758, 
    10.01546, 9.992907, 10.01598, 10.0141, 10.03621, 10.0291, 10.08228, 
    10.0537, 10.13504, 10.16482, 10.25319, 10.30515, 10.35819, 10.38166, 
    10.38881, 10.3918 ;

 WIND =
  8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  3.138606e-09, 3.097616e-09, 3.105489e-09, 3.073129e-09, 3.090987e-09, 
    3.069935e-09, 3.130199e-09, 3.09601e-09, 3.117737e-09, 3.134871e-09, 
    3.0125e-09, 3.071705e-09, 2.953781e-09, 2.989534e-09, 2.901578e-09, 
    2.959273e-09, 2.89026e-09, 2.903216e-09, 2.864647e-09, 2.875575e-09, 
    2.686875e-09, 2.859636e-09, 2.664886e-09, 2.693799e-09, 2.689212e-09, 
    2.860709e-09, 3.059584e-09, 3.019722e-09, 3.061981e-09, 3.056213e-09, 
    3.058801e-09, 3.090612e-09, 3.106929e-09, 3.141799e-09, 3.135403e-09, 
    3.109829e-09, 3.053627e-09, 3.072446e-09, 3.025547e-09, 3.026588e-09, 
    2.976245e-09, 2.998701e-09, 2.916935e-09, 2.939647e-09, 2.875117e-09, 
    2.891034e-09, 2.875859e-09, 2.880442e-09, 2.875799e-09, 2.899226e-09, 
    2.889134e-09, 2.909951e-09, 2.994463e-09, 2.969035e-09, 3.046398e-09, 
    3.095208e-09, 3.128679e-09, 3.152939e-09, 3.149482e-09, 3.142916e-09, 
    3.109681e-09, 3.07918e-09, 3.056397e-09, 3.041372e-09, 3.026738e-09, 
    2.983391e-09, 2.961049e-09, 2.912387e-09, 2.92104e-09, 2.906423e-09, 
    2.892629e-09, 2.869795e-09, 2.873526e-09, 2.863566e-09, 2.906813e-09, 
    2.877901e-09, 2.925994e-09, 2.912654e-09, 3.02275e-09, 3.067344e-09, 
    3.086734e-09, 3.103971e-09, 3.14683e-09, 3.117084e-09, 3.128731e-09, 
    3.101196e-09, 3.083986e-09, 3.092471e-09, 3.040964e-09, 3.060749e-09, 
    2.959737e-09, 3.002283e-09, 2.89423e-09, 2.91926e-09, 2.888305e-09, 
    2.904007e-09, 2.87722e-09, 2.901302e-09, 2.859883e-09, 2.708462e-09, 
    2.857075e-09, 2.692839e-09, 2.90265e-09, 2.875856e-09, 3.092708e-09, 
    3.09132e-09, 3.084876e-09, 3.113436e-09, 3.115205e-09, 3.141973e-09, 
    3.118133e-09, 3.108105e-09, 3.082998e-09, 3.068361e-09, 3.054599e-09, 
    3.024839e-09, 2.992384e-09, 2.948342e-09, 2.917622e-09, 2.897441e-09, 
    2.909779e-09, 2.89888e-09, 2.911069e-09, 2.916825e-09, 2.711564e-09, 
    2.889038e-09, 2.695842e-09, 2.698409e-09, 2.863329e-09, 2.698119e-09, 
    3.090347e-09, 3.098348e-09, 3.126493e-09, 3.104417e-09, 3.144921e-09, 
    3.122093e-09, 3.109138e-09, 3.060324e-09, 3.049845e-09, 3.040192e-09, 
    3.021343e-09, 2.997542e-09, 2.956821e-09, 2.922426e-09, 2.891832e-09, 
    2.894049e-09, 2.893268e-09, 2.886523e-09, 2.903292e-09, 2.883792e-09, 
    2.880546e-09, 2.889047e-09, 2.698754e-09, 2.711402e-09, 2.698464e-09, 
    2.706637e-09, 3.095743e-09, 3.082335e-09, 3.089563e-09, 3.076003e-09, 
    3.085538e-09, 3.043646e-09, 3.031342e-09, 2.975281e-09, 2.998004e-09, 
    2.962038e-09, 2.994307e-09, 2.988527e-09, 2.960866e-09, 2.992545e-09, 
    2.924292e-09, 2.97015e-09, 2.886262e-09, 2.930657e-09, 2.883531e-09, 
    2.891963e-09, 2.878037e-09, 2.865692e-09, 2.707796e-09, 2.682306e-09, 
    2.688124e-09, 2.667288e-09, 3.062601e-09, 3.045662e-09, 3.047151e-09, 
    3.029641e-09, 3.01684e-09, 2.989529e-09, 2.946897e-09, 2.962764e-09, 
    2.933792e-09, 2.928053e-09, 2.972133e-09, 2.944881e-09, 3.034452e-09, 
    3.019545e-09, 3.028405e-09, 3.061252e-09, 2.959081e-09, 3.010503e-09, 
    2.917119e-09, 2.943816e-09, 2.867444e-09, 2.904836e-09, 2.691346e-09, 
    2.664345e-09, 2.639608e-09, 2.611445e-09, 3.036516e-09, 3.047921e-09, 
    3.027577e-09, 2.999932e-09, 2.97482e-09, 2.94217e-09, 2.93888e-09, 
    2.932869e-09, 2.91744e-09, 2.904609e-09, 2.930968e-09, 2.901413e-09, 
    3.016099e-09, 2.954716e-09, 3.052252e-09, 3.022091e-09, 3.001548e-09, 
    3.010527e-09, 2.964592e-09, 2.953999e-09, 2.91184e-09, 2.933462e-09, 
    2.670937e-09, 2.863091e-09, 2.590493e-09, 2.624871e-09, 3.051927e-09, 
    3.036559e-09, 2.984434e-09, 3.008974e-09, 2.940024e-09, 2.923606e-09, 
    2.910422e-09, 2.893757e-09, 2.891976e-09, 2.88222e-09, 2.898245e-09, 
    2.882852e-09, 2.942101e-09, 2.915279e-09, 2.990295e-09, 2.971622e-09, 
    2.980181e-09, 2.98963e-09, 2.960687e-09, 2.930547e-09, 2.929922e-09, 
    2.92041e-09, 2.893971e-09, 2.939752e-09, 2.664873e-09, 2.885748e-09, 
    3.020003e-09, 2.991252e-09, 2.98721e-09, 2.998235e-09, 2.925242e-09, 
    2.951208e-09, 2.882459e-09, 2.900673e-09, 2.87097e-09, 2.88564e-09, 
    2.887813e-09, 2.906948e-09, 2.919008e-09, 2.950004e-09, 2.975796e-09, 
    2.996631e-09, 2.991758e-09, 2.968975e-09, 2.928729e-09, 2.89181e-09, 
    2.899803e-09, 2.873203e-09, 2.944899e-09, 2.91433e-09, 2.926054e-09, 
    2.895712e-09, 2.963186e-09, 2.905471e-09, 2.978365e-09, 2.971807e-09, 
    2.951729e-09, 2.912276e-09, 2.903727e-09, 2.894645e-09, 2.900244e-09, 
    2.927726e-09, 2.932291e-09, 2.952216e-09, 2.957767e-09, 2.973233e-09, 
    2.986174e-09, 2.974342e-09, 2.962031e-09, 2.927719e-09, 2.897572e-09, 
    2.865515e-09, 2.857799e-09, 2.681485e-09, 2.708429e-09, 2.664471e-09, 
    2.701673e-09, 2.638214e-09, 2.902222e-09, 2.702771e-09, 2.950826e-09, 
    2.938972e-09, 2.917798e-09, 2.870566e-09, 2.895853e-09, 2.866335e-09, 
    2.932471e-09, 2.968191e-09, 2.977612e-09, 2.995353e-09, 2.977209e-09, 
    2.978676e-09, 2.961531e-09, 2.967016e-09, 2.926595e-09, 2.948148e-09, 
    2.887865e-09, 2.866568e-09, 2.669451e-09, 2.638323e-09, 2.607579e-09, 
    2.594287e-09, 2.590274e-09, 2.588601e-09 ;

 W_SCALAR =
  0.6251353, 0.6267943, 0.6264719, 0.6278089, 0.6270673, 0.6279426, 
    0.6254717, 0.6268601, 0.6259739, 0.6252846, 0.6303998, 0.6278685, 
    0.6330233, 0.6314129, 0.6354543, 0.6327729, 0.6359942, 0.6353768, 
    0.6372336, 0.6367019, 0.6390741, 0.6374789, 0.6403017, 0.6386933, 
    0.6389451, 0.6374263, 0.6283781, 0.630085, 0.6282769, 0.6285205, 
    0.6284112, 0.6270827, 0.6264129, 0.6250083, 0.6252634, 0.6262949, 
    0.62863, 0.6278377, 0.6298333, 0.6297882, 0.6320065, 0.6310068, 
    0.6347294, 0.6336725, 0.6367241, 0.6359574, 0.6366882, 0.6364666, 
    0.636691, 0.6355664, 0.6360484, 0.6350582, 0.6311942, 0.6323311, 
    0.6289374, 0.6268929, 0.6255327, 0.6245668, 0.6247034, 0.6249638, 
    0.6263009, 0.6275567, 0.6285129, 0.6291522, 0.6297818, 0.631686, 
    0.6326924, 0.6349431, 0.6345371, 0.6352248, 0.6358811, 0.6369825, 
    0.6368012, 0.6372863, 0.6352065, 0.6365892, 0.6343058, 0.6349307, 
    0.6299535, 0.6280515, 0.6272427, 0.6265339, 0.6248084, 0.6260003, 
    0.6255305, 0.6266476, 0.627357, 0.6270062, 0.6291697, 0.628329, 0.632752, 
    0.6308487, 0.6358045, 0.6346204, 0.6360882, 0.6353394, 0.6366222, 
    0.6354678, 0.6374667, 0.6379016, 0.6376044, 0.6387454, 0.6354038, 
    0.6366882, 0.6269963, 0.6270536, 0.6273201, 0.6261482, 0.6260765, 
    0.6250014, 0.625958, 0.6263651, 0.6273981, 0.6280087, 0.628589, 
    0.6298638, 0.6312862, 0.6332723, 0.6346972, 0.6356515, 0.6350664, 
    0.6355829, 0.6350055, 0.6347347, 0.6377387, 0.6360529, 0.6385813, 
    0.6384416, 0.6372979, 0.6384573, 0.6270937, 0.6267644, 0.6256206, 
    0.6265158, 0.6248842, 0.6257978, 0.6263229, 0.6283467, 0.6287908, 
    0.6292027, 0.6300155, 0.631058, 0.6328849, 0.6344721, 0.6359192, 
    0.6358132, 0.6358505, 0.6361737, 0.6353732, 0.636305, 0.6364614, 
    0.6360526, 0.6384228, 0.6377462, 0.6384386, 0.637998, 0.6268715, 
    0.6274255, 0.6271262, 0.627689, 0.6272926, 0.6290547, 0.6295826, 
    0.6320496, 0.6310375, 0.6326477, 0.6312011, 0.6314576, 0.6327004, 
    0.6312793, 0.6343848, 0.6322804, 0.6361862, 0.6340882, 0.6363176, 
    0.635913, 0.6365828, 0.6371825, 0.6379364, 0.6393263, 0.6390046, 
    0.6401659, 0.628251, 0.6289688, 0.6289055, 0.6296563, 0.6302112, 
    0.6314132, 0.6333387, 0.632615, 0.6339433, 0.6342098, 0.6321916, 
    0.6334312, 0.6294489, 0.6300933, 0.6297096, 0.6283076, 0.6327819, 
    0.6304877, 0.6347207, 0.6334803, 0.637097, 0.6352998, 0.6388274, 
    0.6403326, 0.641747, 0.6433983, 0.6293603, 0.6288727, 0.6297455, 
    0.6309522, 0.6320706, 0.6335561, 0.6337079, 0.6339859, 0.6347058, 
    0.6353109, 0.634074, 0.6354625, 0.6302429, 0.6329808, 0.6286885, 
    0.6299827, 0.6308811, 0.6304869, 0.6325322, 0.6330138, 0.634969, 
    0.6339586, 0.6399614, 0.6373093, 0.6446536, 0.6426059, 0.6287023, 
    0.6293585, 0.6316399, 0.6305549, 0.6336551, 0.6344171, 0.6350361, 
    0.6358271, 0.6359124, 0.6363807, 0.6356131, 0.6363503, 0.6335592, 
    0.6348073, 0.6313792, 0.6322145, 0.6318303, 0.6314088, 0.6327093, 
    0.6340935, 0.6341228, 0.6345664, 0.6358159, 0.6336676, 0.6403037, 
    0.63621, 0.6300737, 0.6313363, 0.6315163, 0.6310275, 0.6343407, 
    0.6331412, 0.6363693, 0.6354976, 0.6369254, 0.6362162, 0.6361118, 
    0.6352001, 0.6346322, 0.6331963, 0.6320267, 0.6310984, 0.6313143, 
    0.6323338, 0.6341781, 0.6359202, 0.6355388, 0.636817, 0.6334305, 
    0.6348518, 0.6343027, 0.6357338, 0.6325958, 0.635269, 0.6319116, 
    0.6322063, 0.6331174, 0.6349483, 0.6353527, 0.6357846, 0.6355181, 
    0.6342248, 0.6340128, 0.6330952, 0.6328419, 0.6321421, 0.6315626, 
    0.6320921, 0.6326481, 0.6342253, 0.635645, 0.6371911, 0.637569, 
    0.6393728, 0.6379049, 0.6403264, 0.6382684, 0.6418286, 0.6354235, 
    0.6382074, 0.6331588, 0.6337036, 0.6346887, 0.6369447, 0.635727, 
    0.6371508, 0.6340044, 0.632369, 0.6319454, 0.6311548, 0.6319634, 
    0.6318977, 0.6326709, 0.6324225, 0.6342776, 0.6332815, 0.6361092, 
    0.6371396, 0.6400443, 0.6418217, 0.6436279, 0.6444244, 0.6446668, 
    0.6447681,
  0.546122, 0.5481663, 0.547769, 0.5494168, 0.5485029, 0.5495816, 0.5465365, 
    0.5482475, 0.5471554, 0.546306, 0.5526108, 0.5494903, 0.5558459, 
    0.5538599, 0.5588443, 0.5555371, 0.5595104, 0.5587488, 0.5610396, 
    0.5603836, 0.5633109, 0.5613422, 0.564826, 0.5628408, 0.5631516, 
    0.5612773, 0.5501185, 0.5522227, 0.5499938, 0.550294, 0.5501593, 
    0.5485218, 0.5476962, 0.5459654, 0.5462797, 0.5475509, 0.550429, 
    0.5494523, 0.5519123, 0.5518568, 0.554592, 0.5533592, 0.5579502, 
    0.5566465, 0.560411, 0.5594651, 0.5603666, 0.5600932, 0.5603701, 
    0.5589826, 0.5595772, 0.5583557, 0.5535902, 0.5549921, 0.550808, 
    0.5482879, 0.5466116, 0.5454214, 0.5455897, 0.5459106, 0.5475582, 
    0.5491059, 0.5502846, 0.5510727, 0.5518488, 0.5541967, 0.5554377, 
    0.5582138, 0.5577129, 0.5585612, 0.5593709, 0.5607297, 0.5605062, 
    0.5611046, 0.5585387, 0.5602445, 0.5574276, 0.5581985, 0.5520605, 
    0.5497158, 0.548719, 0.5478454, 0.5457191, 0.5471878, 0.546609, 
    0.5479856, 0.5488598, 0.5484275, 0.5510942, 0.5500579, 0.5555113, 
    0.5531643, 0.5592765, 0.5578157, 0.5596264, 0.5587026, 0.5602852, 
    0.558861, 0.5613272, 0.5618639, 0.5614972, 0.5629051, 0.558782, 
    0.5603667, 0.5484154, 0.5484859, 0.5488144, 0.5473701, 0.5472817, 
    0.5459569, 0.5471357, 0.5476375, 0.5489105, 0.5496632, 0.5503784, 
    0.55195, 0.5537037, 0.556153, 0.5579104, 0.5590876, 0.5583658, 0.5590031, 
    0.5582907, 0.5579567, 0.5616629, 0.5595828, 0.5627027, 0.5625302, 
    0.5611189, 0.5625496, 0.5485354, 0.5481296, 0.5467199, 0.5478232, 
    0.5458125, 0.5469384, 0.5475854, 0.5500798, 0.5506272, 0.5511349, 
    0.552137, 0.5534223, 0.5556751, 0.5576328, 0.559418, 0.5592872, 
    0.5593333, 0.5597319, 0.5587444, 0.559894, 0.5600869, 0.5595825, 
    0.5625071, 0.561672, 0.5625265, 0.5619829, 0.5482615, 0.5489443, 
    0.5485753, 0.5492691, 0.5487804, 0.5509526, 0.5516033, 0.5546451, 
    0.5533971, 0.5553826, 0.5535988, 0.5539151, 0.5554476, 0.5536952, 
    0.557525, 0.5549297, 0.5597474, 0.5571592, 0.5599095, 0.5594102, 
    0.5602366, 0.5609765, 0.5619068, 0.5636221, 0.563225, 0.5646584, 
    0.5499617, 0.5508466, 0.5507686, 0.5516941, 0.5523783, 0.5538603, 
    0.5562348, 0.5553423, 0.5569804, 0.5573092, 0.5548201, 0.5563489, 
    0.5514385, 0.5522329, 0.5517598, 0.5500316, 0.5555482, 0.5527192, 
    0.5579395, 0.5564095, 0.5608711, 0.5586538, 0.5630064, 0.5648642, 
    0.5666101, 0.5686489, 0.5513292, 0.5507281, 0.5518041, 0.5532919, 
    0.5546709, 0.5565029, 0.5566902, 0.5570331, 0.5579211, 0.5586674, 
    0.5571417, 0.5588545, 0.5524173, 0.5557935, 0.550501, 0.5520964, 
    0.5532042, 0.5527182, 0.5552402, 0.5558341, 0.5582457, 0.5569993, 
    0.564406, 0.561133, 0.5701991, 0.5676705, 0.5505182, 0.551327, 0.5541399, 
    0.552802, 0.5566251, 0.5575649, 0.5583284, 0.5593042, 0.5594094, 
    0.5599873, 0.5590403, 0.5599499, 0.5565068, 0.5580462, 0.5538184, 
    0.5548484, 0.5543746, 0.5538548, 0.5554585, 0.5571658, 0.557202, 
    0.5577492, 0.5592904, 0.5566405, 0.5648284, 0.5597767, 0.5522088, 
    0.5537655, 0.5539874, 0.5533847, 0.5574707, 0.5559913, 0.5599732, 
    0.5588979, 0.5606593, 0.5597843, 0.5596555, 0.5585308, 0.5578303, 
    0.5560592, 0.5546168, 0.5534721, 0.5537383, 0.5549955, 0.5572701, 
    0.5594191, 0.5589486, 0.5605255, 0.5563481, 0.5581011, 0.5574238, 
    0.5591892, 0.5553185, 0.5586159, 0.5544749, 0.5548382, 0.5559619, 
    0.5582201, 0.558719, 0.5592519, 0.558923, 0.5573277, 0.5570661, 
    0.5559345, 0.5556221, 0.5547591, 0.5540445, 0.5546975, 0.5553831, 
    0.5573283, 0.5590797, 0.5609871, 0.5614535, 0.5636794, 0.561868, 
    0.5648565, 0.5623165, 0.5667108, 0.5588064, 0.5622413, 0.5560129, 
    0.5566849, 0.5579, 0.5606831, 0.5591809, 0.5609375, 0.5570559, 0.555039, 
    0.5545165, 0.5535418, 0.5545388, 0.5544577, 0.5554113, 0.5551049, 
    0.5573929, 0.5561642, 0.5596523, 0.5609236, 0.5645083, 0.5667024, 
    0.5689324, 0.5699161, 0.5702153, 0.5703405,
  0.5139007, 0.5161509, 0.5157135, 0.5175276, 0.5165213, 0.5177091, 
    0.5143569, 0.5162403, 0.5150381, 0.5141032, 0.5210451, 0.5176085, 
    0.5246094, 0.5224211, 0.5279146, 0.5242691, 0.528649, 0.5278093, 
    0.5303354, 0.5296119, 0.5328408, 0.5306692, 0.5345126, 0.5323222, 
    0.5326651, 0.5305976, 0.5183002, 0.5206175, 0.5181628, 0.5184935, 
    0.5183451, 0.5165422, 0.5156334, 0.5137285, 0.5140744, 0.5154734, 
    0.5186421, 0.5175667, 0.5202757, 0.5202146, 0.5232277, 0.5218695, 
    0.5269288, 0.5254918, 0.5296421, 0.528599, 0.5295932, 0.5292917, 
    0.5295971, 0.5280671, 0.5287228, 0.5273759, 0.522124, 0.5236686, 
    0.5190594, 0.5162846, 0.5144396, 0.5131298, 0.513315, 0.5136681, 
    0.5154815, 0.5171853, 0.5184832, 0.5193509, 0.5202057, 0.5227922, 
    0.5241597, 0.5272194, 0.5266673, 0.5276024, 0.5284952, 0.5299937, 
    0.5297471, 0.5304071, 0.5275776, 0.5294585, 0.5263528, 0.5272026, 
    0.5204389, 0.5178568, 0.5167593, 0.5157976, 0.5134574, 0.5150738, 
    0.5144367, 0.5159519, 0.5169144, 0.5164384, 0.5193747, 0.5182335, 
    0.5242407, 0.5216548, 0.5283911, 0.5267806, 0.5287769, 0.5277584, 
    0.5295034, 0.5279329, 0.5306526, 0.5312446, 0.5308401, 0.5323932, 
    0.5278459, 0.5295932, 0.5164251, 0.5165027, 0.5168644, 0.5152744, 
    0.5151771, 0.513719, 0.5150164, 0.5155687, 0.5169701, 0.5177988, 
    0.5185864, 0.5203171, 0.522249, 0.5249479, 0.526885, 0.5281828, 
    0.5273871, 0.5280896, 0.5273043, 0.5269361, 0.5310228, 0.5287289, 
    0.5321699, 0.5319796, 0.5304228, 0.532001, 0.5165572, 0.5161104, 
    0.5145588, 0.5157731, 0.5135602, 0.5147992, 0.5155115, 0.5182576, 
    0.5188603, 0.5194194, 0.5205231, 0.521939, 0.5244212, 0.526579, 
    0.5285471, 0.5284029, 0.5284537, 0.5288932, 0.5278044, 0.529072, 
    0.5292847, 0.5287285, 0.5319541, 0.531033, 0.5319755, 0.5313758, 
    0.5162556, 0.5170074, 0.5166012, 0.517365, 0.516827, 0.5192186, 
    0.5199353, 0.5232862, 0.5219113, 0.5240989, 0.5221335, 0.5224819, 
    0.5241706, 0.5222397, 0.5264602, 0.5235998, 0.5289103, 0.5260569, 
    0.5290891, 0.5285386, 0.5294499, 0.5302659, 0.5312918, 0.5331842, 
    0.5327461, 0.5343277, 0.5181276, 0.519102, 0.519016, 0.5200353, 0.520789, 
    0.5224215, 0.5250381, 0.5240544, 0.5258599, 0.5262222, 0.5234791, 
    0.5251638, 0.5197538, 0.5206288, 0.5201077, 0.5182045, 0.5242813, 
    0.5211644, 0.5269171, 0.5252306, 0.5301495, 0.5277045, 0.5325049, 
    0.5345548, 0.5364818, 0.5387327, 0.5196335, 0.5189716, 0.5201565, 
    0.5217954, 0.5233147, 0.5253335, 0.5255399, 0.5259179, 0.5268968, 
    0.5277196, 0.5260376, 0.5279258, 0.5208319, 0.5245516, 0.5187214, 
    0.5204785, 0.5216987, 0.5211633, 0.5239419, 0.5245965, 0.5272546, 
    0.5258808, 0.5340492, 0.5304384, 0.5404447, 0.5376524, 0.5187403, 
    0.5196311, 0.5227296, 0.5212557, 0.5254682, 0.5265041, 0.5273458, 
    0.5284217, 0.5285377, 0.5291749, 0.5281307, 0.5291336, 0.5253378, 
    0.5270347, 0.5223754, 0.5235103, 0.5229882, 0.5224155, 0.5241826, 
    0.5260642, 0.5261041, 0.5267072, 0.5284064, 0.5254852, 0.5345153, 
    0.5289426, 0.5206022, 0.5223171, 0.5225616, 0.5218976, 0.5264003, 
    0.5247697, 0.5291593, 0.5279736, 0.529916, 0.528951, 0.528809, 0.5275689, 
    0.5267966, 0.5248445, 0.5232551, 0.5219939, 0.5222871, 0.5236723, 
    0.5261792, 0.5285484, 0.5280296, 0.5297685, 0.5251629, 0.5270953, 
    0.5263487, 0.5282949, 0.5240283, 0.5276627, 0.5230986, 0.5234991, 
    0.5247373, 0.5272264, 0.5277764, 0.528364, 0.5280014, 0.5262427, 
    0.5259544, 0.5247071, 0.5243628, 0.5234119, 0.5226244, 0.523344, 
    0.5240994, 0.5262434, 0.5281741, 0.5302775, 0.5307919, 0.5332475, 
    0.531249, 0.5345464, 0.5317438, 0.536593, 0.5278728, 0.5316609, 
    0.5247936, 0.5255342, 0.5268735, 0.5299422, 0.5282857, 0.5302228, 
    0.525943, 0.5237203, 0.5231445, 0.5220706, 0.5231691, 0.5230798, 
    0.5241305, 0.5237929, 0.5263145, 0.5249603, 0.5288056, 0.5302075, 
    0.5341621, 0.5365836, 0.5390458, 0.5401321, 0.5404627, 0.5406008,
  0.5071029, 0.5094935, 0.5090288, 0.5109567, 0.5098872, 0.5111496, 
    0.5075876, 0.5095885, 0.5083112, 0.507318, 0.5146972, 0.5110427, 
    0.5184905, 0.5161612, 0.5220108, 0.5181282, 0.5227934, 0.5218986, 
    0.5245908, 0.5238196, 0.5272627, 0.5249467, 0.5290464, 0.5267095, 
    0.5270752, 0.5248704, 0.5117781, 0.5142424, 0.5116321, 0.5119835, 
    0.5118257, 0.5099094, 0.5089437, 0.50692, 0.5072874, 0.5087736, 
    0.5121415, 0.5109982, 0.5138788, 0.5138137, 0.5170196, 0.5155743, 
    0.5209606, 0.51943, 0.5238518, 0.5227401, 0.5237997, 0.5234783, 
    0.5238038, 0.5221732, 0.5228719, 0.5214369, 0.5158451, 0.517489, 
    0.5125853, 0.5096357, 0.5076753, 0.5062842, 0.5064809, 0.5068558, 
    0.5087823, 0.5105929, 0.5119725, 0.5128953, 0.5138044, 0.5165562, 
    0.5180117, 0.5212702, 0.520682, 0.5216782, 0.5226294, 0.5242265, 
    0.5239637, 0.5246673, 0.5216517, 0.5236561, 0.520347, 0.5212523, 
    0.5140524, 0.5113066, 0.5101401, 0.5091181, 0.5066321, 0.5083491, 
    0.5076723, 0.5092821, 0.5103049, 0.5097991, 0.5129206, 0.5117072, 
    0.5180979, 0.5153458, 0.5225185, 0.5208027, 0.5229297, 0.5218444, 
    0.5237039, 0.5220304, 0.5249291, 0.5255602, 0.525129, 0.5267852, 
    0.5219376, 0.5237997, 0.5097849, 0.5098674, 0.5102518, 0.5085623, 
    0.5084589, 0.50691, 0.5082881, 0.508875, 0.5103642, 0.5112451, 0.5120823, 
    0.5139229, 0.5159781, 0.5188509, 0.520914, 0.5222966, 0.5214487, 
    0.5221973, 0.5213605, 0.5209683, 0.5253238, 0.5228785, 0.526547, 
    0.526344, 0.5246841, 0.5263669, 0.5099254, 0.5094505, 0.507802, 
    0.5090922, 0.5067413, 0.5080574, 0.508814, 0.5117327, 0.5123736, 
    0.5129681, 0.514142, 0.5156483, 0.5182902, 0.5205879, 0.5226848, 
    0.5225312, 0.5225852, 0.5230536, 0.5218934, 0.5232441, 0.5234709, 
    0.5228781, 0.5263168, 0.5253346, 0.5263397, 0.5257002, 0.5096048, 
    0.5104038, 0.5099721, 0.5107839, 0.510212, 0.5127546, 0.5135168, 
    0.5170819, 0.5156187, 0.517947, 0.5158552, 0.5162259, 0.5180233, 
    0.5159682, 0.5204614, 0.5174158, 0.5230719, 0.5200319, 0.5232623, 
    0.5226757, 0.5236469, 0.5245167, 0.5256106, 0.527629, 0.5271617, 
    0.5288491, 0.5115945, 0.5126305, 0.5125392, 0.5136232, 0.5144247, 
    0.5161617, 0.5189469, 0.5178996, 0.5198221, 0.520208, 0.5172873, 
    0.5190808, 0.5133237, 0.5142543, 0.5137001, 0.5116764, 0.5181412, 
    0.5148242, 0.5209481, 0.5191519, 0.5243927, 0.521787, 0.5269044, 
    0.5290914, 0.5311483, 0.5335522, 0.5131958, 0.5124919, 0.513752, 
    0.5154954, 0.5171123, 0.5192615, 0.5194813, 0.5198839, 0.5209265, 
    0.521803, 0.5200114, 0.5220227, 0.5144705, 0.518429, 0.5122259, 
    0.5140945, 0.5153926, 0.514823, 0.5177799, 0.5184767, 0.5213076, 
    0.5198442, 0.5285518, 0.5247006, 0.5353815, 0.5323984, 0.512246, 
    0.5131932, 0.5164895, 0.5149213, 0.5194049, 0.5205082, 0.5214048, 
    0.5225511, 0.5226747, 0.5233538, 0.5222411, 0.5233098, 0.5192661, 
    0.5210734, 0.5161126, 0.5173204, 0.5167648, 0.5161553, 0.5180361, 
    0.5200396, 0.5200821, 0.5207245, 0.5225348, 0.519423, 0.5290493, 
    0.5231063, 0.5142261, 0.5160505, 0.5163108, 0.5156042, 0.5203976, 
    0.5186611, 0.5233372, 0.5220737, 0.5241438, 0.5231152, 0.5229639, 
    0.5216425, 0.5208198, 0.5187408, 0.5170488, 0.5157066, 0.5160187, 
    0.5174929, 0.5201621, 0.5226861, 0.5221333, 0.5239865, 0.5190799, 
    0.5211378, 0.5203426, 0.5224159, 0.5178719, 0.5217424, 0.5168823, 
    0.5173085, 0.5186266, 0.5212776, 0.5218636, 0.5224897, 0.5221033, 
    0.5202298, 0.5199227, 0.5185946, 0.5182279, 0.5172157, 0.5163777, 
    0.5171434, 0.5179476, 0.5202305, 0.5222873, 0.5245291, 0.5250775, 
    0.5276965, 0.525565, 0.5290824, 0.5260926, 0.531267, 0.5219662, 
    0.5260041, 0.5186865, 0.5194752, 0.5209016, 0.5241717, 0.5224062, 
    0.5244708, 0.5199106, 0.5175439, 0.5169312, 0.5157883, 0.5169573, 
    0.5168622, 0.5179807, 0.5176213, 0.5203062, 0.5188641, 0.5229602, 
    0.5244544, 0.5286723, 0.531257, 0.5338867, 0.5350474, 0.5354007, 0.5355483,
  0.5311316, 0.5336009, 0.5331207, 0.5351133, 0.5340078, 0.5353128, 
    0.5316319, 0.5336991, 0.5323793, 0.5313537, 0.5389836, 0.5352023, 
    0.5429142, 0.5404999, 0.5465672, 0.5425386, 0.54738, 0.5464507, 
    0.5492477, 0.5484462, 0.5520267, 0.5496178, 0.5538836, 0.5514511, 
    0.5518317, 0.5495384, 0.5359627, 0.5385127, 0.5358117, 0.5361752, 
    0.5360121, 0.5340307, 0.5330327, 0.5309427, 0.5313221, 0.532857, 
    0.5363387, 0.5351563, 0.5381364, 0.538069, 0.5413894, 0.539892, 
    0.5454769, 0.5438886, 0.5484797, 0.5473246, 0.5484254, 0.5480916, 
    0.5484298, 0.5467359, 0.5474616, 0.5459713, 0.5401724, 0.5418758, 
    0.5367977, 0.5337478, 0.5317227, 0.5302864, 0.5304894, 0.5308765, 
    0.532866, 0.5347372, 0.5361639, 0.5371185, 0.5380594, 0.5409091, 
    0.5424178, 0.5457982, 0.5451877, 0.5462219, 0.5472097, 0.5488691, 
    0.5485959, 0.5493273, 0.5461944, 0.5482763, 0.54484, 0.5457796, 0.538316, 
    0.5354752, 0.5342691, 0.533213, 0.5306455, 0.5324185, 0.5317195, 
    0.5333824, 0.5344395, 0.5339166, 0.5371446, 0.5358894, 0.5425072, 
    0.5396553, 0.5470945, 0.545313, 0.5475215, 0.5463943, 0.548326, 
    0.5465875, 0.5495994, 0.5502557, 0.5498072, 0.5515298, 0.5464912, 
    0.5484256, 0.533902, 0.5339873, 0.5343845, 0.5326387, 0.5325319, 
    0.5309324, 0.5323555, 0.5329617, 0.5345007, 0.5354115, 0.5362774, 
    0.538182, 0.5403102, 0.5432879, 0.5454285, 0.546864, 0.5459836, 
    0.5467609, 0.5458921, 0.5454848, 0.5500098, 0.5474684, 0.551282, 
    0.5510709, 0.5493447, 0.5510947, 0.5340472, 0.5335565, 0.5318534, 
    0.5331861, 0.5307582, 0.5321172, 0.5328988, 0.5359158, 0.5365788, 
    0.5371939, 0.5384088, 0.5399686, 0.5427065, 0.5450901, 0.5472671, 
    0.5471076, 0.5471638, 0.5476503, 0.5464453, 0.5478482, 0.5480838, 
    0.547468, 0.5510426, 0.550021, 0.5510664, 0.5504012, 0.5337159, 
    0.5345417, 0.5340955, 0.5349346, 0.5343435, 0.5369729, 0.5377616, 
    0.5414539, 0.5399379, 0.5423506, 0.5401829, 0.540567, 0.5424298, 0.5403, 
    0.5449588, 0.5418, 0.5476693, 0.544513, 0.5478672, 0.5472577, 0.5482667, 
    0.5491707, 0.5503081, 0.5524079, 0.5519215, 0.5536782, 0.5357729, 
    0.5368446, 0.53675, 0.5378717, 0.5387015, 0.5405004, 0.5433876, 
    0.5423016, 0.5442954, 0.5446958, 0.5416667, 0.5435264, 0.5375618, 
    0.538525, 0.5379514, 0.5358575, 0.5425521, 0.5391151, 0.5454639, 
    0.5436001, 0.5490418, 0.5463348, 0.5516539, 0.5539305, 0.5560735, 
    0.5585806, 0.5374294, 0.5367011, 0.5380051, 0.5398102, 0.5414854, 
    0.5437139, 0.5439418, 0.5443595, 0.5454414, 0.5463514, 0.5444918, 
    0.5465796, 0.5387488, 0.5428504, 0.5364259, 0.5383596, 0.5397037, 
    0.5391139, 0.5421774, 0.5428999, 0.5458371, 0.5443184, 0.5533686, 
    0.5493619, 0.56049, 0.5573769, 0.5364467, 0.5374268, 0.54084, 0.5392156, 
    0.5438626, 0.5450073, 0.545938, 0.5471284, 0.5472568, 0.5479622, 
    0.5468063, 0.5479165, 0.5437186, 0.545594, 0.5404496, 0.5417011, 
    0.5411252, 0.5404938, 0.542443, 0.5445211, 0.5445652, 0.5452318, 
    0.5471114, 0.5438814, 0.5538865, 0.547705, 0.5384958, 0.5403852, 
    0.5406549, 0.5399229, 0.5448925, 0.5430912, 0.547945, 0.5466325, 
    0.5487831, 0.5477143, 0.5475571, 0.5461848, 0.5453308, 0.5431738, 
    0.5414196, 0.540029, 0.5403523, 0.54188, 0.5446482, 0.5472685, 0.5466944, 
    0.5486196, 0.5435255, 0.5456609, 0.5448354, 0.546988, 0.5422728, 
    0.5462885, 0.5412471, 0.5416888, 0.5430554, 0.5458059, 0.5464143, 
    0.5470645, 0.5466632, 0.5447184, 0.5443997, 0.5430221, 0.542642, 
    0.5415926, 0.5407242, 0.5415177, 0.5423512, 0.5447191, 0.5468544, 
    0.5491836, 0.5497537, 0.5524781, 0.5502606, 0.5539211, 0.5508093, 
    0.5561973, 0.5465209, 0.5507173, 0.5431175, 0.5439355, 0.5454156, 
    0.5488122, 0.5469778, 0.549123, 0.5443872, 0.5419328, 0.5412977, 
    0.5401136, 0.5413248, 0.5412263, 0.5423856, 0.542013, 0.5447977, 
    0.5433016, 0.5475532, 0.5491059, 0.5534941, 0.5561869, 0.5589296, 
    0.5601412, 0.56051, 0.5606642,
  0.5352567, 0.5381001, 0.5375467, 0.539844, 0.538569, 0.5400741, 0.5358325, 
    0.5382132, 0.5366928, 0.5355123, 0.5443151, 0.5399465, 0.5488689, 
    0.5460703, 0.5531131, 0.5484331, 0.554059, 0.5529775, 0.556235, 
    0.5553008, 0.5594782, 0.5566664, 0.5616494, 0.5588059, 0.5592504, 
    0.5565737, 0.5408241, 0.5437704, 0.5406498, 0.5410694, 0.5408811, 
    0.5385954, 0.5374454, 0.5350395, 0.5354759, 0.537243, 0.5412582, 
    0.5398935, 0.5433353, 0.5432574, 0.5471008, 0.5453663, 0.5518451, 0.55, 
    0.5553398, 0.5539945, 0.5552766, 0.5548877, 0.5552816, 0.5533093, 
    0.554154, 0.5524199, 0.545691, 0.5476646, 0.5417883, 0.5382693, 
    0.5359369, 0.5342847, 0.5345182, 0.5349634, 0.5372533, 0.5394101, 
    0.5410564, 0.5421589, 0.5432462, 0.5465443, 0.548293, 0.5522187, 
    0.551509, 0.5527113, 0.5538608, 0.5557936, 0.5554752, 0.5563276, 
    0.5526794, 0.5551028, 0.551105, 0.552197, 0.543543, 0.5402614, 0.5388703, 
    0.5376531, 0.5346977, 0.5367379, 0.5359333, 0.5378482, 0.5390668, 
    0.5384639, 0.5421891, 0.5407395, 0.5483968, 0.5450924, 0.5537266, 
    0.5516546, 0.5542238, 0.552912, 0.5551607, 0.5531367, 0.5566449, 
    0.5574104, 0.5568873, 0.5588979, 0.5530246, 0.5552766, 0.5384471, 
    0.5385454, 0.5390034, 0.5369915, 0.5368685, 0.5350276, 0.5366654, 
    0.5373636, 0.5391374, 0.540188, 0.5411875, 0.543388, 0.5458506, 
    0.5493026, 0.5517888, 0.5534584, 0.5524343, 0.5533384, 0.5523278, 
    0.5518543, 0.5571236, 0.5541619, 0.5586085, 0.5583619, 0.5563479, 
    0.5583897, 0.5386144, 0.5380488, 0.5360874, 0.5376221, 0.5348273, 
    0.536391, 0.5372912, 0.54077, 0.5415354, 0.5422459, 0.5436503, 0.545455, 
    0.5486279, 0.5513955, 0.5539277, 0.5537419, 0.5538073, 0.5543738, 
    0.5529712, 0.5546042, 0.5548786, 0.5541614, 0.5583289, 0.5571367, 
    0.5583566, 0.5575802, 0.5382326, 0.5391846, 0.5386701, 0.5396377, 
    0.538956, 0.5419907, 0.5429021, 0.5471756, 0.5454196, 0.5482152, 
    0.5457032, 0.5461479, 0.5483069, 0.5458387, 0.5512429, 0.5475767, 
    0.5543958, 0.550725, 0.5546262, 0.5539167, 0.5550916, 0.5561451, 
    0.5574716, 0.5599237, 0.5593554, 0.561409, 0.540605, 0.5418425, 
    0.5417333, 0.5430293, 0.5439888, 0.5460709, 0.5494182, 0.5481583, 
    0.5504722, 0.5509374, 0.5474222, 0.5495794, 0.5426711, 0.5437847, 
    0.5431215, 0.5407027, 0.5484488, 0.5444672, 0.5518299, 0.549665, 
    0.5559949, 0.5528427, 0.5590427, 0.5617042, 0.5642141, 0.5671557, 
    0.5425181, 0.5416767, 0.5431835, 0.5452718, 0.5472121, 0.5497969, 
    0.5500616, 0.5505467, 0.5518039, 0.552862, 0.5507003, 0.5531275, 
    0.5440435, 0.5487949, 0.5413589, 0.5435934, 0.5451484, 0.5444658, 
    0.5480143, 0.5488523, 0.5522639, 0.5504989, 0.5610469, 0.556368, 
    0.5694002, 0.5657426, 0.5413829, 0.5425151, 0.5464643, 0.5445836, 
    0.5499696, 0.5512993, 0.5523812, 0.5537661, 0.5539156, 0.5547369, 
    0.5533913, 0.5546837, 0.5498025, 0.5519812, 0.546012, 0.5474621, 
    0.5467947, 0.5460632, 0.5483224, 0.5507344, 0.5507857, 0.5515602, 
    0.5537463, 0.5499915, 0.5616528, 0.5544374, 0.5437509, 0.5459375, 
    0.5462497, 0.5454021, 0.5511659, 0.5490742, 0.5547169, 0.553189, 
    0.5556933, 0.5544482, 0.5542652, 0.5526682, 0.5516752, 0.5491701, 
    0.5471358, 0.545525, 0.5458993, 0.5476694, 0.550882, 0.5539292, 0.553261, 
    0.5555028, 0.5495782, 0.552059, 0.5510997, 0.5536027, 0.5481249, 
    0.5527889, 0.5469359, 0.5474478, 0.5490327, 0.5522276, 0.5529352, 
    0.5536917, 0.5532248, 0.5509636, 0.5505934, 0.5489941, 0.5485531, 
    0.5473363, 0.54633, 0.5472495, 0.5482159, 0.5509644, 0.5534472, 
    0.5561602, 0.5568249, 0.5600058, 0.5574162, 0.5616933, 0.5580566, 
    0.5643591, 0.5530592, 0.5579491, 0.5491048, 0.5500543, 0.5517739, 
    0.5557271, 0.5535909, 0.5560895, 0.550579, 0.5477307, 0.5469945, 
    0.5456229, 0.5470259, 0.5469117, 0.5482557, 0.5478237, 0.5510558, 
    0.5493185, 0.5542607, 0.5560697, 0.5611937, 0.564347, 0.5675656, 
    0.5689899, 0.5694237, 0.5696052,
  0.5840973, 0.5875084, 0.5868435, 0.5896071, 0.5880722, 0.5898844, 0.584787, 
    0.5876443, 0.5858185, 0.5844033, 0.5950112, 0.5897306, 0.6005507, 
    0.597142, 0.6057469, 0.600019, 0.6069095, 0.6055803, 0.6095902, 
    0.6084383, 0.6136027, 0.6101228, 0.6163003, 0.6127692, 0.6133202, 
    0.6100085, 0.5907888, 0.594351, 0.5905786, 0.5910849, 0.5908576, 
    0.588104, 0.5867218, 0.5838373, 0.5843598, 0.5864788, 0.5913127, 
    0.5896668, 0.5938239, 0.5937297, 0.5983955, 0.5962867, 0.6041909, 
    0.6019322, 0.6084863, 0.6068302, 0.6084084, 0.6079293, 0.6084146, 
    0.605988, 0.6070263, 0.6048959, 0.5966811, 0.5990822, 0.591953, 
    0.5877119, 0.5849121, 0.5829342, 0.5832134, 0.5837461, 0.5864912, 
    0.5890844, 0.5910691, 0.5924008, 0.5937161, 0.5977183, 0.599848, 
    0.6046491, 0.603779, 0.6052536, 0.6066657, 0.6090457, 0.6086532, 
    0.6097046, 0.6052144, 0.6081943, 0.6032842, 0.6046225, 0.5940755, 
    0.5901102, 0.5884346, 0.5869713, 0.5834281, 0.5858726, 0.5849077, 
    0.5872058, 0.5886711, 0.5879459, 0.5924373, 0.5906867, 0.5999746, 
    0.5959541, 0.6065008, 0.6039575, 0.6071122, 0.6054999, 0.6082657, 
    0.6057759, 0.6100964, 0.6110422, 0.6103957, 0.6128832, 0.6056382, 
    0.6084085, 0.5879256, 0.5880438, 0.5885949, 0.5861769, 0.5860293, 
    0.583823, 0.5857856, 0.5866236, 0.5887561, 0.5900217, 0.5912274, 
    0.5938878, 0.596875, 0.6010801, 0.604122, 0.6061711, 0.6049135, 
    0.6060237, 0.6047829, 0.6042023, 0.6106877, 0.6070361, 0.6125247, 
    0.6122194, 0.6097297, 0.6122538, 0.5881268, 0.5874467, 0.5850925, 
    0.5869341, 0.5835832, 0.5854565, 0.5865366, 0.5907236, 0.5916475, 
    0.5925061, 0.5942054, 0.5963944, 0.6002566, 0.60364, 0.6067479, 
    0.6065195, 0.6065999, 0.6072967, 0.6055726, 0.6075803, 0.6079181, 
    0.6070355, 0.6121785, 0.6107038, 0.6122129, 0.6112521, 0.5876677, 
    0.5888129, 0.5881938, 0.5893586, 0.5885379, 0.5921975, 0.5932996, 
    0.5984865, 0.5963513, 0.5997532, 0.5966958, 0.5972363, 0.5998651, 
    0.5968605, 0.6034531, 0.598975, 0.6073238, 0.6028191, 0.6076075, 
    0.6067345, 0.6081806, 0.6094794, 0.6111178, 0.6141555, 0.6134504, 
    0.6160011, 0.5905246, 0.5920184, 0.5918865, 0.5934536, 0.5946156, 
    0.5971426, 0.6012213, 0.5996838, 0.6025097, 0.603079, 0.5987869, 
    0.6014182, 0.5930202, 0.5943683, 0.5935651, 0.5906424, 0.6000381, 
    0.5951956, 0.6041725, 0.6015228, 0.609294, 0.6054149, 0.6130627, 
    0.6163685, 0.6194988, 0.6231837, 0.5928351, 0.5918182, 0.5936402, 
    0.5961719, 0.5985309, 0.6016841, 0.6020076, 0.6026009, 0.6041405, 
    0.6054386, 0.6027889, 0.6057645, 0.5946819, 0.6004604, 0.5914344, 
    0.5941365, 0.5960222, 0.5951939, 0.5995083, 0.6005304, 0.6047046, 
    0.6025425, 0.6155508, 0.6097545, 0.6260076, 0.6214114, 0.5914633, 
    0.5928315, 0.597621, 0.5953367, 0.6018951, 0.6035222, 0.6048485, 
    0.6065493, 0.606733, 0.6077437, 0.6060886, 0.6076782, 0.6016908, 
    0.6043578, 0.5970711, 0.5988355, 0.5980229, 0.5971333, 0.5998839, 
    0.6028305, 0.6028933, 0.6038418, 0.606525, 0.6019219, 0.6163046, 
    0.607375, 0.5943274, 0.5969806, 0.5973601, 0.5963302, 0.6033589, 
    0.6008013, 0.607719, 0.6058401, 0.6089221, 0.6073884, 0.6071631, 
    0.6052006, 0.6039827, 0.6009184, 0.5984381, 0.5964794, 0.5969341, 
    0.599088, 0.6030113, 0.6067499, 0.6059287, 0.6086873, 0.6014168, 
    0.6044532, 0.6032777, 0.6063484, 0.5996431, 0.6053487, 0.5981948, 
    0.598818, 0.6007506, 0.6046601, 0.6055284, 0.6064579, 0.6058841, 
    0.6031111, 0.6026581, 0.6007035, 0.6001653, 0.5986822, 0.5974577, 
    0.5985765, 0.599754, 0.6031122, 0.6061573, 0.609498, 0.6103187, 
    0.6142573, 0.6110493, 0.6163548, 0.6118414, 0.61968, 0.6056807, 
    0.6117085, 0.6008386, 0.6019986, 0.6041037, 0.6089638, 0.6063339, 
    0.6094108, 0.6026403, 0.5991626, 0.5982661, 0.5965983, 0.5983043, 
    0.5981653, 0.5998026, 0.5992759, 0.603224, 0.6010996, 0.6071576, 
    0.6093863, 0.6157333, 0.6196648, 0.6236987, 0.6254905, 0.6260372, 
    0.6262659,
  0.6622251, 0.667787, 0.6666976, 0.6712429, 0.6687129, 0.6717015, 0.6633443, 
    0.6680101, 0.6650231, 0.6627214, 0.6802661, 0.6714472, 0.6897115, 
    0.6838751, 0.6987642, 0.6887959, 0.7008165, 0.6984711, 0.7055876, 
    0.7035306, 0.7128337, 0.7065421, 0.7177787, 0.711318, 0.7123192, 
    0.706337, 0.6732006, 0.679154, 0.6728517, 0.6736924, 0.6733148, 
    0.6687651, 0.6664985, 0.6618038, 0.6626506, 0.6661011, 0.6740712, 
    0.6713416, 0.678268, 0.6781098, 0.6860123, 0.682423, 0.6960332, 
    0.6920996, 0.7036162, 0.7006762, 0.7034775, 0.7026251, 0.7034886, 
    0.6991889, 0.7010233, 0.6972684, 0.683092, 0.6871875, 0.6751375, 
    0.6681209, 0.6635476, 0.6603438, 0.6607947, 0.6616562, 0.6661214, 
    0.6703798, 0.6736662, 0.6758848, 0.6780871, 0.6848564, 0.688502, 
    0.6968355, 0.6953132, 0.6978964, 0.7003853, 0.7046142, 0.7039137, 
    0.7057924, 0.6978275, 0.7030964, 0.6944497, 0.696789, 0.6786907, 
    0.6720755, 0.669309, 0.6669067, 0.6611419, 0.6651114, 0.6635405, 
    0.6672908, 0.6696985, 0.6685052, 0.6759457, 0.6730312, 0.6887195, 
    0.6818596, 0.7000939, 0.6956249, 0.7011755, 0.6983296, 0.7032234, 
    0.6988153, 0.7064946, 0.7081949, 0.707032, 0.7115248, 0.6985729, 
    0.7034777, 0.6684719, 0.6686662, 0.6695728, 0.6656079, 0.665367, 
    0.6617807, 0.6649695, 0.6663378, 0.6698384, 0.6719288, 0.6739292, 
    0.6783753, 0.6834213, 0.6906251, 0.6959125, 0.6995119, 0.6972993, 
    0.6992519, 0.6970701, 0.6960531, 0.7075568, 0.7010406, 0.7108742, 
    0.710321, 0.7058373, 0.7103833, 0.6688027, 0.6676859, 0.6638409, 
    0.6668458, 0.6613927, 0.6644333, 0.6661956, 0.6730922, 0.6746284, 
    0.6760606, 0.6789091, 0.6826056, 0.6892048, 0.6950704, 0.7005307, 
    0.7001271, 0.7002691, 0.7015024, 0.6984575, 0.7020053, 0.7026053, 
    0.7010396, 0.710247, 0.7075858, 0.7103093, 0.7085733, 0.6680484, 
    0.6699321, 0.6689128, 0.6708325, 0.6694789, 0.6755454, 0.6773884, 
    0.6861679, 0.6825325, 0.688339, 0.683117, 0.6840357, 0.6885313, 
    0.6833967, 0.6947443, 0.6870038, 0.7015504, 0.6936398, 0.7020535, 
    0.7005069, 0.703072, 0.7053893, 0.7083312, 0.713842, 0.7125562, 
    0.7172273, 0.672762, 0.6752465, 0.6750265, 0.6776466, 0.6795995, 
    0.6838763, 0.6908692, 0.6882197, 0.6931019, 0.6940922, 0.6866817, 
    0.6912096, 0.6769205, 0.6791831, 0.6778336, 0.6729575, 0.6888287, 
    0.6805773, 0.6960008, 0.6913906, 0.7050577, 0.69818, 0.711851, 0.7179045, 
    0.7237219, 0.7306815, 0.6766108, 0.6749127, 0.6779597, 0.6822283, 
    0.6862438, 0.6916698, 0.6922304, 0.6932604, 0.6959449, 0.6982217, 
    0.6935872, 0.6987953, 0.6797111, 0.6895558, 0.6742736, 0.6787933, 
    0.6819748, 0.6805745, 0.6879184, 0.6896765, 0.6969327, 0.6931587, 
    0.7163987, 0.7058818, 0.7360995, 0.7273188, 0.6743218, 0.6766047, 
    0.6846905, 0.6808156, 0.6920354, 0.6948648, 0.6971852, 0.7001796, 
    0.7005044, 0.7022954, 0.6993665, 0.702179, 0.6916814, 0.6963252, 
    0.6837546, 0.6867648, 0.685376, 0.6838604, 0.6885635, 0.6936597, 
    0.6937689, 0.6954229, 0.7001367, 0.6920817, 0.7177866, 0.7016411, 
    0.6791143, 0.6836007, 0.6842463, 0.6824966, 0.6945799, 0.6901437, 
    0.7022516, 0.6989285, 0.7043934, 0.7016648, 0.7012656, 0.6978035, 
    0.6956691, 0.6903458, 0.686085, 0.6827497, 0.6835218, 0.6871974, 
    0.6939742, 0.7005342, 0.6990844, 0.7039744, 0.6912072, 0.6964923, 
    0.6944383, 0.6998248, 0.6881498, 0.6980637, 0.6856694, 0.686735, 
    0.6900563, 0.6968548, 0.6983797, 0.7000182, 0.6990059, 0.6941482, 
    0.6933598, 0.689975, 0.6890477, 0.6865026, 0.6844125, 0.6863217, 
    0.6883404, 0.6941499, 0.6994876, 0.7054225, 0.7068936, 0.7140281, 
    0.7082077, 0.7178792, 0.7096372, 0.7240614, 0.6986477, 0.709397, 
    0.6902081, 0.6922147, 0.6958807, 0.7044679, 0.6997992, 0.7052665, 
    0.6933289, 0.6873254, 0.6857913, 0.6829515, 0.6858565, 0.6856191, 
    0.6884239, 0.6875196, 0.6943448, 0.6906586, 0.7012557, 0.7052227, 
    0.7167343, 0.7240329, 0.731664, 0.7351019, 0.7361569, 0.7365991,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.540215e-11, 3.555962e-11, 3.552893e-11, 3.5656e-11, 3.558547e-11, 
    3.566862e-11, 3.54339e-11, 3.556559e-11, 3.548146e-11, 3.541603e-11, 
    3.59025e-11, 3.566137e-11, 3.615359e-11, 3.59994e-11, 3.638688e-11, 
    3.612946e-11, 3.64388e-11, 3.637941e-11, 3.655819e-11, 3.650689e-11, 
    3.673565e-11, 3.658175e-11, 3.685438e-11, 3.669885e-11, 3.67231e-11, 
    3.657647e-11, 3.57102e-11, 3.587273e-11, 3.570048e-11, 3.572366e-11, 
    3.571322e-11, 3.558675e-11, 3.552302e-11, 3.538981e-11, 3.541394e-11, 
    3.551177e-11, 3.57338e-11, 3.565835e-11, 3.584848e-11, 3.584419e-11, 
    3.605606e-11, 3.596046e-11, 3.631713e-11, 3.621561e-11, 3.650899e-11, 
    3.643509e-11, 3.650543e-11, 3.648404e-11, 3.65056e-11, 3.639733e-11, 
    3.644362e-11, 3.63484e-11, 3.597881e-11, 3.608751e-11, 3.576331e-11, 
    3.556857e-11, 3.54395e-11, 3.534797e-11, 3.536083e-11, 3.538549e-11, 
    3.551226e-11, 3.563159e-11, 3.572261e-11, 3.578346e-11, 3.584346e-11, 
    3.602523e-11, 3.612159e-11, 3.633753e-11, 3.629856e-11, 3.636454e-11, 
    3.64277e-11, 3.65337e-11, 3.651623e-11, 3.65629e-11, 3.636262e-11, 
    3.649566e-11, 3.627603e-11, 3.633605e-11, 3.585998e-11, 3.567887e-11, 
    3.56018e-11, 3.553447e-11, 3.537074e-11, 3.548375e-11, 3.543914e-11, 
    3.554516e-11, 3.561255e-11, 3.557916e-11, 3.578508e-11, 3.570491e-11, 
    3.612725e-11, 3.594518e-11, 3.642038e-11, 3.630648e-11, 3.644757e-11, 
    3.637555e-11, 3.649889e-11, 3.638782e-11, 3.658023e-11, 3.662219e-11, 
    3.659342e-11, 3.670362e-11, 3.638142e-11, 3.650502e-11, 3.557844e-11, 
    3.558388e-11, 3.560918e-11, 3.549773e-11, 3.549091e-11, 3.538891e-11, 
    3.547958e-11, 3.551822e-11, 3.561637e-11, 3.567439e-11, 3.572959e-11, 
    3.585114e-11, 3.598691e-11, 3.617702e-11, 3.631381e-11, 3.64055e-11, 
    3.634923e-11, 3.639884e-11, 3.634329e-11, 3.631722e-11, 3.660636e-11, 
    3.644389e-11, 3.668766e-11, 3.667417e-11, 3.65637e-11, 3.667558e-11, 
    3.558763e-11, 3.555628e-11, 3.544764e-11, 3.553259e-11, 3.537774e-11, 
    3.546435e-11, 3.551411e-11, 3.570649e-11, 3.574881e-11, 3.578805e-11, 
    3.586555e-11, 3.596506e-11, 3.613985e-11, 3.629207e-11, 3.643123e-11, 
    3.642097e-11, 3.642454e-11, 3.645556e-11, 3.637854e-11, 3.646814e-11, 
    3.648312e-11, 3.644379e-11, 3.667225e-11, 3.660695e-11, 3.667373e-11, 
    3.663115e-11, 3.556641e-11, 3.561901e-11, 3.55905e-11, 3.564402e-11, 
    3.560622e-11, 3.577394e-11, 3.58242e-11, 3.605987e-11, 3.596308e-11, 
    3.611713e-11, 3.597866e-11, 3.600318e-11, 3.612195e-11, 3.598605e-11, 
    3.628351e-11, 3.608163e-11, 3.645673e-11, 3.625484e-11, 3.64693e-11, 
    3.643031e-11, 3.649474e-11, 3.655251e-11, 3.662519e-11, 3.67594e-11, 
    3.672824e-11, 3.684058e-11, 3.569751e-11, 3.576579e-11, 3.575979e-11, 
    3.583131e-11, 3.588421e-11, 3.599908e-11, 3.61834e-11, 3.6114e-11, 
    3.624131e-11, 3.626689e-11, 3.607334e-11, 3.619207e-11, 3.581118e-11, 
    3.587254e-11, 3.583598e-11, 3.570229e-11, 3.61296e-11, 3.591006e-11, 
    3.631559e-11, 3.619647e-11, 3.654416e-11, 3.63711e-11, 3.67111e-11, 
    3.685657e-11, 3.699372e-11, 3.715392e-11, 3.58031e-11, 3.575659e-11, 
    3.583976e-11, 3.595491e-11, 3.606185e-11, 3.620419e-11, 3.621873e-11, 
    3.624534e-11, 3.631444e-11, 3.637259e-11, 3.625364e-11, 3.638706e-11, 
    3.588668e-11, 3.614867e-11, 3.573849e-11, 3.586183e-11, 3.59476e-11, 
    3.590998e-11, 3.610558e-11, 3.615165e-11, 3.63392e-11, 3.624223e-11, 
    3.682051e-11, 3.656438e-11, 3.727608e-11, 3.707687e-11, 3.574031e-11, 
    3.580279e-11, 3.602058e-11, 3.591691e-11, 3.621361e-11, 3.628673e-11, 
    3.634614e-11, 3.642218e-11, 3.643033e-11, 3.647541e-11, 3.640148e-11, 
    3.647243e-11, 3.620407e-11, 3.632392e-11, 3.599529e-11, 3.607512e-11, 
    3.603835e-11, 3.599797e-11, 3.61224e-11, 3.625507e-11, 3.625791e-11, 
    3.63004e-11, 3.642025e-11, 3.621409e-11, 3.685333e-11, 3.645809e-11, 
    3.587098e-11, 3.599145e-11, 3.600869e-11, 3.596198e-11, 3.627929e-11, 
    3.616421e-11, 3.647432e-11, 3.639039e-11, 3.652779e-11, 3.645948e-11, 
    3.644934e-11, 3.636166e-11, 3.630698e-11, 3.616917e-11, 3.605705e-11, 
    3.59683e-11, 3.598886e-11, 3.608638e-11, 3.626309e-11, 3.643057e-11, 
    3.639381e-11, 3.651686e-11, 3.619127e-11, 3.632767e-11, 3.627483e-11, 
    3.641244e-11, 3.611198e-11, 3.636831e-11, 3.604646e-11, 3.607461e-11, 
    3.616182e-11, 3.633747e-11, 3.637637e-11, 3.641789e-11, 3.63922e-11, 
    3.626788e-11, 3.624749e-11, 3.615945e-11, 3.613509e-11, 3.606812e-11, 
    3.601258e-11, 3.606324e-11, 3.611636e-11, 3.626765e-11, 3.640402e-11, 
    3.655285e-11, 3.658931e-11, 3.676328e-11, 3.662152e-11, 3.685533e-11, 
    3.665633e-11, 3.700093e-11, 3.638316e-11, 3.665141e-11, 3.616582e-11, 
    3.6218e-11, 3.631247e-11, 3.652946e-11, 3.641227e-11, 3.654931e-11, 
    3.624668e-11, 3.608978e-11, 3.604925e-11, 3.597363e-11, 3.60509e-11, 
    3.604462e-11, 3.611861e-11, 3.609476e-11, 3.627256e-11, 3.617701e-11, 
    3.644856e-11, 3.654778e-11, 3.682833e-11, 3.700045e-11, 3.717597e-11, 
    3.725342e-11, 3.727701e-11, 3.728683e-11,
  1.802e-11, 1.815729e-11, 1.813058e-11, 1.824152e-11, 1.817996e-11, 
    1.825264e-11, 1.804781e-11, 1.816274e-11, 1.808935e-11, 1.803236e-11, 
    1.845753e-11, 1.824648e-11, 1.867786e-11, 1.854252e-11, 1.888324e-11, 
    1.865676e-11, 1.892903e-11, 1.887672e-11, 1.903441e-11, 1.898919e-11, 
    1.919136e-11, 1.90553e-11, 1.929651e-11, 1.915886e-11, 1.918036e-11, 
    1.905081e-11, 1.828891e-11, 1.84312e-11, 1.828048e-11, 1.830075e-11, 
    1.829166e-11, 1.818122e-11, 1.812564e-11, 1.800954e-11, 1.80306e-11, 
    1.81159e-11, 1.830986e-11, 1.824395e-11, 1.841029e-11, 1.840653e-11, 
    1.859237e-11, 1.850849e-11, 1.882191e-11, 1.873264e-11, 1.899107e-11, 
    1.892595e-11, 1.898801e-11, 1.896919e-11, 1.898825e-11, 1.889278e-11, 
    1.893366e-11, 1.884974e-11, 1.852418e-11, 1.861963e-11, 1.833549e-11, 
    1.816541e-11, 1.805284e-11, 1.797311e-11, 1.798437e-11, 1.800585e-11, 
    1.811639e-11, 1.822059e-11, 1.830014e-11, 1.835343e-11, 1.840599e-11, 
    1.856537e-11, 1.865e-11, 1.883997e-11, 1.880566e-11, 1.886382e-11, 
    1.891948e-11, 1.901303e-11, 1.899762e-11, 1.903888e-11, 1.88623e-11, 
    1.897958e-11, 1.878612e-11, 1.883895e-11, 1.842019e-11, 1.826173e-11, 
    1.819444e-11, 1.813571e-11, 1.799303e-11, 1.809151e-11, 1.805266e-11, 
    1.814515e-11, 1.8204e-11, 1.817489e-11, 1.835489e-11, 1.828483e-11, 
    1.865502e-11, 1.849522e-11, 1.891298e-11, 1.88127e-11, 1.893705e-11, 
    1.887356e-11, 1.898239e-11, 1.888444e-11, 1.905425e-11, 1.90913e-11, 
    1.906597e-11, 1.916334e-11, 1.887901e-11, 1.8988e-11, 1.817407e-11, 
    1.817882e-11, 1.820095e-11, 1.810375e-11, 1.809782e-11, 1.800896e-11, 
    1.808803e-11, 1.812173e-11, 1.820743e-11, 1.825817e-11, 1.830647e-11, 
    1.841283e-11, 1.853188e-11, 1.869886e-11, 1.881919e-11, 1.890001e-11, 
    1.885044e-11, 1.88942e-11, 1.884528e-11, 1.882238e-11, 1.907742e-11, 
    1.893404e-11, 1.914932e-11, 1.913739e-11, 1.903985e-11, 1.913874e-11, 
    1.818215e-11, 1.815484e-11, 1.806012e-11, 1.813423e-11, 1.79993e-11, 
    1.807477e-11, 1.811821e-11, 1.828627e-11, 1.832329e-11, 1.835762e-11, 
    1.842552e-11, 1.851278e-11, 1.866623e-11, 1.880014e-11, 1.892272e-11, 
    1.891373e-11, 1.89169e-11, 1.894431e-11, 1.887642e-11, 1.895546e-11, 
    1.896873e-11, 1.893403e-11, 1.91358e-11, 1.907808e-11, 1.913714e-11, 
    1.909956e-11, 1.816372e-11, 1.82097e-11, 1.818485e-11, 1.823158e-11, 
    1.819864e-11, 1.834525e-11, 1.83893e-11, 1.859594e-11, 1.851105e-11, 
    1.864625e-11, 1.852478e-11, 1.854628e-11, 1.865063e-11, 1.853134e-11, 
    1.879273e-11, 1.861533e-11, 1.894537e-11, 1.876764e-11, 1.895653e-11, 
    1.892219e-11, 1.897907e-11, 1.903004e-11, 1.909429e-11, 1.921297e-11, 
    1.918547e-11, 1.92849e-11, 1.827833e-11, 1.83381e-11, 1.833286e-11, 
    1.83955e-11, 1.844187e-11, 1.854257e-11, 1.870448e-11, 1.864353e-11, 
    1.875549e-11, 1.877799e-11, 1.860793e-11, 1.871226e-11, 1.837817e-11, 
    1.843197e-11, 1.839994e-11, 1.828303e-11, 1.865755e-11, 1.846497e-11, 
    1.882118e-11, 1.871642e-11, 1.902277e-11, 1.887017e-11, 1.917033e-11, 
    1.929912e-11, 1.942071e-11, 1.956305e-11, 1.837078e-11, 1.833013e-11, 
    1.840296e-11, 1.850388e-11, 1.859775e-11, 1.87228e-11, 1.873562e-11, 
    1.875909e-11, 1.881994e-11, 1.887114e-11, 1.876649e-11, 1.888399e-11, 
    1.844442e-11, 1.867431e-11, 1.831475e-11, 1.842271e-11, 1.849793e-11, 
    1.846494e-11, 1.863658e-11, 1.867711e-11, 1.884216e-11, 1.875679e-11, 
    1.926729e-11, 1.904079e-11, 1.967175e-11, 1.949466e-11, 1.831593e-11, 
    1.837065e-11, 1.856156e-11, 1.847063e-11, 1.873117e-11, 1.87955e-11, 
    1.884788e-11, 1.891488e-11, 1.892213e-11, 1.896188e-11, 1.889676e-11, 
    1.895931e-11, 1.872307e-11, 1.882851e-11, 1.853973e-11, 1.860985e-11, 
    1.857758e-11, 1.85422e-11, 1.865148e-11, 1.876813e-11, 1.877066e-11, 
    1.880812e-11, 1.891377e-11, 1.873223e-11, 1.929653e-11, 1.894724e-11, 
    1.843039e-11, 1.853606e-11, 1.855121e-11, 1.851023e-11, 1.878905e-11, 
    1.868784e-11, 1.896091e-11, 1.888697e-11, 1.900819e-11, 1.894792e-11, 
    1.893905e-11, 1.886176e-11, 1.88137e-11, 1.869247e-11, 1.859406e-11, 
    1.851618e-11, 1.853428e-11, 1.861987e-11, 1.877528e-11, 1.892277e-11, 
    1.889043e-11, 1.899897e-11, 1.871223e-11, 1.883225e-11, 1.878582e-11, 
    1.890698e-11, 1.864191e-11, 1.886745e-11, 1.858441e-11, 1.860917e-11, 
    1.868583e-11, 1.884038e-11, 1.887468e-11, 1.891128e-11, 1.88887e-11, 
    1.877924e-11, 1.876134e-11, 1.868397e-11, 1.866262e-11, 1.860378e-11, 
    1.855511e-11, 1.859957e-11, 1.86463e-11, 1.87793e-11, 1.889944e-11, 
    1.903077e-11, 1.906297e-11, 1.921687e-11, 1.909153e-11, 1.929848e-11, 
    1.912242e-11, 1.94276e-11, 1.88806e-11, 1.911731e-11, 1.868933e-11, 
    1.873527e-11, 1.881843e-11, 1.900976e-11, 1.890641e-11, 1.902731e-11, 
    1.876064e-11, 1.862281e-11, 1.858724e-11, 1.85209e-11, 1.858876e-11, 
    1.858324e-11, 1.864826e-11, 1.862736e-11, 1.878372e-11, 1.869967e-11, 
    1.893882e-11, 1.902637e-11, 1.927446e-11, 1.942709e-11, 1.958297e-11, 
    1.965191e-11, 1.967291e-11, 1.968169e-11,
  1.693475e-11, 1.708502e-11, 1.705576e-11, 1.717728e-11, 1.710984e-11, 
    1.718947e-11, 1.696518e-11, 1.709099e-11, 1.701063e-11, 1.694827e-11, 
    1.741415e-11, 1.718272e-11, 1.765603e-11, 1.750738e-11, 1.788183e-11, 
    1.763285e-11, 1.793221e-11, 1.787464e-11, 1.80482e-11, 1.799841e-11, 
    1.822114e-11, 1.80712e-11, 1.833708e-11, 1.81853e-11, 1.8209e-11, 
    1.806626e-11, 1.72292e-11, 1.738526e-11, 1.721997e-11, 1.724218e-11, 
    1.723222e-11, 1.711122e-11, 1.705038e-11, 1.69233e-11, 1.694634e-11, 
    1.70397e-11, 1.725217e-11, 1.717993e-11, 1.736229e-11, 1.735816e-11, 
    1.756211e-11, 1.747003e-11, 1.781436e-11, 1.771621e-11, 1.800048e-11, 
    1.792881e-11, 1.799711e-11, 1.797639e-11, 1.799738e-11, 1.789231e-11, 
    1.79373e-11, 1.784496e-11, 1.748725e-11, 1.759205e-11, 1.728027e-11, 
    1.709393e-11, 1.697068e-11, 1.688345e-11, 1.689577e-11, 1.691926e-11, 
    1.704024e-11, 1.715434e-11, 1.724151e-11, 1.729992e-11, 1.735757e-11, 
    1.753249e-11, 1.762542e-11, 1.783423e-11, 1.779648e-11, 1.786045e-11, 
    1.792168e-11, 1.802466e-11, 1.80077e-11, 1.805312e-11, 1.785878e-11, 
    1.798784e-11, 1.777499e-11, 1.78331e-11, 1.737319e-11, 1.719941e-11, 
    1.712572e-11, 1.706139e-11, 1.690524e-11, 1.7013e-11, 1.697049e-11, 
    1.707172e-11, 1.713617e-11, 1.710429e-11, 1.730152e-11, 1.722473e-11, 
    1.763093e-11, 1.745547e-11, 1.791454e-11, 1.780423e-11, 1.794102e-11, 
    1.787117e-11, 1.799093e-11, 1.788313e-11, 1.807005e-11, 1.811087e-11, 
    1.808296e-11, 1.819023e-11, 1.787716e-11, 1.799711e-11, 1.710339e-11, 
    1.710859e-11, 1.713282e-11, 1.70264e-11, 1.70199e-11, 1.692267e-11, 
    1.700918e-11, 1.704608e-11, 1.713992e-11, 1.719552e-11, 1.724845e-11, 
    1.736507e-11, 1.749571e-11, 1.76791e-11, 1.781137e-11, 1.790026e-11, 
    1.784574e-11, 1.789387e-11, 1.784006e-11, 1.781487e-11, 1.809557e-11, 
    1.793771e-11, 1.817479e-11, 1.816164e-11, 1.805421e-11, 1.816312e-11, 
    1.711224e-11, 1.708233e-11, 1.697864e-11, 1.705976e-11, 1.691209e-11, 
    1.699467e-11, 1.704224e-11, 1.722631e-11, 1.726689e-11, 1.730453e-11, 
    1.737898e-11, 1.747473e-11, 1.764324e-11, 1.779043e-11, 1.792525e-11, 
    1.791536e-11, 1.791884e-11, 1.794901e-11, 1.787431e-11, 1.796129e-11, 
    1.797589e-11, 1.79377e-11, 1.815988e-11, 1.809629e-11, 1.816136e-11, 
    1.811995e-11, 1.709205e-11, 1.714241e-11, 1.711519e-11, 1.716639e-11, 
    1.713031e-11, 1.729097e-11, 1.733927e-11, 1.756605e-11, 1.747284e-11, 
    1.76213e-11, 1.74879e-11, 1.751151e-11, 1.762613e-11, 1.749511e-11, 
    1.778228e-11, 1.758734e-11, 1.795018e-11, 1.775471e-11, 1.796246e-11, 
    1.792467e-11, 1.798727e-11, 1.80434e-11, 1.811415e-11, 1.824496e-11, 
    1.821463e-11, 1.832426e-11, 1.72176e-11, 1.728313e-11, 1.727737e-11, 
    1.734606e-11, 1.739693e-11, 1.750743e-11, 1.768526e-11, 1.76183e-11, 
    1.774133e-11, 1.776606e-11, 1.75792e-11, 1.769382e-11, 1.732706e-11, 
    1.738608e-11, 1.735093e-11, 1.722276e-11, 1.763371e-11, 1.742228e-11, 
    1.781355e-11, 1.769839e-11, 1.803539e-11, 1.786744e-11, 1.819795e-11, 
    1.833998e-11, 1.847412e-11, 1.863135e-11, 1.731895e-11, 1.727438e-11, 
    1.735424e-11, 1.746497e-11, 1.756802e-11, 1.77054e-11, 1.771949e-11, 
    1.774528e-11, 1.781218e-11, 1.786851e-11, 1.775343e-11, 1.788264e-11, 
    1.739976e-11, 1.765212e-11, 1.725753e-11, 1.737593e-11, 1.745844e-11, 
    1.742224e-11, 1.761066e-11, 1.765519e-11, 1.783664e-11, 1.774275e-11, 
    1.830487e-11, 1.805525e-11, 1.875147e-11, 1.855579e-11, 1.725881e-11, 
    1.731881e-11, 1.752829e-11, 1.742849e-11, 1.771459e-11, 1.778532e-11, 
    1.784291e-11, 1.791663e-11, 1.79246e-11, 1.796835e-11, 1.789669e-11, 
    1.796552e-11, 1.770569e-11, 1.782161e-11, 1.750431e-11, 1.75813e-11, 
    1.754587e-11, 1.750703e-11, 1.762702e-11, 1.775523e-11, 1.7758e-11, 
    1.779919e-11, 1.791546e-11, 1.771576e-11, 1.833715e-11, 1.795229e-11, 
    1.738433e-11, 1.750031e-11, 1.751692e-11, 1.747193e-11, 1.777822e-11, 
    1.766698e-11, 1.796729e-11, 1.788592e-11, 1.801933e-11, 1.795298e-11, 
    1.794323e-11, 1.785819e-11, 1.780532e-11, 1.767207e-11, 1.756397e-11, 
    1.747846e-11, 1.749833e-11, 1.759231e-11, 1.77631e-11, 1.792532e-11, 
    1.788973e-11, 1.800918e-11, 1.769378e-11, 1.782573e-11, 1.777468e-11, 
    1.790794e-11, 1.761652e-11, 1.786449e-11, 1.755337e-11, 1.758056e-11, 
    1.766477e-11, 1.783469e-11, 1.78724e-11, 1.791267e-11, 1.788782e-11, 
    1.776744e-11, 1.774776e-11, 1.766273e-11, 1.763927e-11, 1.757464e-11, 
    1.752119e-11, 1.757002e-11, 1.762135e-11, 1.77675e-11, 1.789965e-11, 
    1.804419e-11, 1.807965e-11, 1.824927e-11, 1.811113e-11, 1.83393e-11, 
    1.81452e-11, 1.848177e-11, 1.787894e-11, 1.813954e-11, 1.766861e-11, 
    1.77191e-11, 1.781055e-11, 1.802108e-11, 1.790731e-11, 1.80404e-11, 
    1.774699e-11, 1.759555e-11, 1.755648e-11, 1.748365e-11, 1.755815e-11, 
    1.755208e-11, 1.762349e-11, 1.760053e-11, 1.777236e-11, 1.767997e-11, 
    1.794298e-11, 1.803936e-11, 1.831275e-11, 1.848118e-11, 1.865333e-11, 
    1.872953e-11, 1.875275e-11, 1.876246e-11,
  1.733278e-11, 1.749766e-11, 1.746555e-11, 1.759896e-11, 1.75249e-11, 
    1.761234e-11, 1.736615e-11, 1.750422e-11, 1.741602e-11, 1.73476e-11, 
    1.785927e-11, 1.760493e-11, 1.812536e-11, 1.796177e-11, 1.837409e-11, 
    1.809986e-11, 1.842963e-11, 1.836616e-11, 1.855753e-11, 1.850261e-11, 
    1.874842e-11, 1.85829e-11, 1.887646e-11, 1.870883e-11, 1.8735e-11, 
    1.857745e-11, 1.765598e-11, 1.78275e-11, 1.764584e-11, 1.767024e-11, 
    1.765929e-11, 1.752642e-11, 1.745965e-11, 1.732022e-11, 1.734549e-11, 
    1.744792e-11, 1.768122e-11, 1.760186e-11, 1.780221e-11, 1.779767e-11, 
    1.802198e-11, 1.792068e-11, 1.829973e-11, 1.819161e-11, 1.85049e-11, 
    1.842586e-11, 1.850118e-11, 1.847833e-11, 1.850148e-11, 1.838563e-11, 
    1.843522e-11, 1.833345e-11, 1.793963e-11, 1.805494e-11, 1.771209e-11, 
    1.750746e-11, 1.73722e-11, 1.727652e-11, 1.729003e-11, 1.73158e-11, 
    1.744852e-11, 1.757376e-11, 1.76695e-11, 1.773368e-11, 1.779702e-11, 
    1.798942e-11, 1.809167e-11, 1.832162e-11, 1.828003e-11, 1.835053e-11, 
    1.841801e-11, 1.853157e-11, 1.851285e-11, 1.856297e-11, 1.834867e-11, 
    1.849096e-11, 1.825635e-11, 1.832037e-11, 1.781424e-11, 1.762326e-11, 
    1.754236e-11, 1.747172e-11, 1.730042e-11, 1.741863e-11, 1.737198e-11, 
    1.748306e-11, 1.755381e-11, 1.75188e-11, 1.773543e-11, 1.765106e-11, 
    1.809774e-11, 1.790468e-11, 1.841013e-11, 1.828856e-11, 1.843933e-11, 
    1.836232e-11, 1.849436e-11, 1.837551e-11, 1.858163e-11, 1.862667e-11, 
    1.859589e-11, 1.871426e-11, 1.836893e-11, 1.850118e-11, 1.751782e-11, 
    1.752353e-11, 1.755013e-11, 1.743333e-11, 1.74262e-11, 1.731953e-11, 
    1.741443e-11, 1.745492e-11, 1.755792e-11, 1.761898e-11, 1.767712e-11, 
    1.780528e-11, 1.794893e-11, 1.815076e-11, 1.829643e-11, 1.839439e-11, 
    1.833429e-11, 1.838735e-11, 1.832804e-11, 1.830028e-11, 1.86098e-11, 
    1.843568e-11, 1.869722e-11, 1.86827e-11, 1.856416e-11, 1.868434e-11, 
    1.752754e-11, 1.74947e-11, 1.738092e-11, 1.746993e-11, 1.730793e-11, 
    1.739852e-11, 1.745071e-11, 1.765281e-11, 1.769738e-11, 1.773874e-11, 
    1.782057e-11, 1.792586e-11, 1.811128e-11, 1.827336e-11, 1.842194e-11, 
    1.841103e-11, 1.841487e-11, 1.844814e-11, 1.836579e-11, 1.846167e-11, 
    1.847778e-11, 1.843567e-11, 1.868076e-11, 1.861058e-11, 1.868239e-11, 
    1.863669e-11, 1.750537e-11, 1.756066e-11, 1.753077e-11, 1.758699e-11, 
    1.754738e-11, 1.772385e-11, 1.777693e-11, 1.802633e-11, 1.792378e-11, 
    1.808713e-11, 1.794034e-11, 1.796631e-11, 1.809246e-11, 1.794826e-11, 
    1.82644e-11, 1.804977e-11, 1.844943e-11, 1.823403e-11, 1.846297e-11, 
    1.84213e-11, 1.849032e-11, 1.855223e-11, 1.863029e-11, 1.87747e-11, 
    1.874121e-11, 1.886229e-11, 1.764324e-11, 1.771523e-11, 1.770889e-11, 
    1.778438e-11, 1.78403e-11, 1.796182e-11, 1.815754e-11, 1.808382e-11, 
    1.821927e-11, 1.824652e-11, 1.804078e-11, 1.816696e-11, 1.77635e-11, 
    1.782838e-11, 1.778974e-11, 1.764891e-11, 1.810079e-11, 1.786819e-11, 
    1.829884e-11, 1.817199e-11, 1.85434e-11, 1.835823e-11, 1.872279e-11, 
    1.887967e-11, 1.902791e-11, 1.920184e-11, 1.775459e-11, 1.77056e-11, 
    1.779337e-11, 1.791513e-11, 1.802849e-11, 1.817971e-11, 1.819522e-11, 
    1.822363e-11, 1.829732e-11, 1.835939e-11, 1.823261e-11, 1.837497e-11, 
    1.784344e-11, 1.812105e-11, 1.768709e-11, 1.781723e-11, 1.790795e-11, 
    1.786813e-11, 1.80754e-11, 1.812442e-11, 1.832428e-11, 1.822084e-11, 
    1.884089e-11, 1.856532e-11, 1.93348e-11, 1.911825e-11, 1.76885e-11, 
    1.775442e-11, 1.798478e-11, 1.7875e-11, 1.818983e-11, 1.826773e-11, 
    1.833118e-11, 1.841244e-11, 1.842123e-11, 1.846947e-11, 1.839045e-11, 
    1.846634e-11, 1.818003e-11, 1.830771e-11, 1.795838e-11, 1.80431e-11, 
    1.800411e-11, 1.796137e-11, 1.809342e-11, 1.82346e-11, 1.823763e-11, 
    1.828302e-11, 1.84112e-11, 1.819111e-11, 1.887658e-11, 1.84518e-11, 
    1.782644e-11, 1.7954e-11, 1.797226e-11, 1.792277e-11, 1.825991e-11, 
    1.81374e-11, 1.846829e-11, 1.837858e-11, 1.852568e-11, 1.845251e-11, 
    1.844176e-11, 1.834802e-11, 1.828977e-11, 1.814301e-11, 1.802402e-11, 
    1.792995e-11, 1.79518e-11, 1.805522e-11, 1.824326e-11, 1.842202e-11, 
    1.838279e-11, 1.851448e-11, 1.816691e-11, 1.831226e-11, 1.825602e-11, 
    1.840286e-11, 1.808186e-11, 1.835501e-11, 1.801236e-11, 1.804228e-11, 
    1.813498e-11, 1.832214e-11, 1.836368e-11, 1.840808e-11, 1.838068e-11, 
    1.824805e-11, 1.822636e-11, 1.813272e-11, 1.81069e-11, 1.803576e-11, 
    1.797696e-11, 1.803068e-11, 1.808718e-11, 1.82481e-11, 1.839372e-11, 
    1.855312e-11, 1.859223e-11, 1.877949e-11, 1.862698e-11, 1.887896e-11, 
    1.866462e-11, 1.903641e-11, 1.837091e-11, 1.865834e-11, 1.81392e-11, 
    1.819479e-11, 1.829554e-11, 1.852763e-11, 1.840216e-11, 1.854894e-11, 
    1.822552e-11, 1.805879e-11, 1.801578e-11, 1.793566e-11, 1.801762e-11, 
    1.801094e-11, 1.808952e-11, 1.806425e-11, 1.825346e-11, 1.815171e-11, 
    1.844149e-11, 1.854778e-11, 1.884958e-11, 1.903573e-11, 1.922615e-11, 
    1.93105e-11, 1.93362e-11, 1.934696e-11,
  1.885987e-11, 1.9036e-11, 1.900169e-11, 1.914429e-11, 1.906511e-11, 
    1.91586e-11, 1.88955e-11, 1.904302e-11, 1.894877e-11, 1.887569e-11, 
    1.94228e-11, 1.915067e-11, 1.97078e-11, 1.953252e-11, 1.997456e-11, 
    1.968047e-11, 2.003417e-11, 1.996604e-11, 2.017149e-11, 2.011251e-11, 
    2.037665e-11, 2.019875e-11, 2.051436e-11, 2.033409e-11, 2.036223e-11, 
    2.01929e-11, 1.920525e-11, 1.93888e-11, 1.919441e-11, 1.922051e-11, 
    1.920879e-11, 1.906674e-11, 1.899539e-11, 1.884645e-11, 1.887344e-11, 
    1.898286e-11, 1.923225e-11, 1.914738e-11, 1.936169e-11, 1.935683e-11, 
    1.959701e-11, 1.948851e-11, 1.989476e-11, 1.97788e-11, 2.011497e-11, 
    2.003012e-11, 2.011098e-11, 2.008644e-11, 2.01113e-11, 1.998694e-11, 
    2.004017e-11, 1.993094e-11, 1.95088e-11, 1.963232e-11, 1.926526e-11, 
    1.904649e-11, 1.890196e-11, 1.879979e-11, 1.881421e-11, 1.884173e-11, 
    1.89835e-11, 1.911734e-11, 1.921971e-11, 1.928836e-11, 1.935614e-11, 
    1.956215e-11, 1.967169e-11, 1.991826e-11, 1.987363e-11, 1.994927e-11, 
    2.002169e-11, 2.014361e-11, 2.012352e-11, 2.017734e-11, 1.994727e-11, 
    2.010001e-11, 1.984823e-11, 1.991691e-11, 1.937461e-11, 1.917026e-11, 
    1.908379e-11, 1.900828e-11, 1.882531e-11, 1.895156e-11, 1.890173e-11, 
    1.902039e-11, 1.909602e-11, 1.905859e-11, 1.929023e-11, 1.919999e-11, 
    1.96782e-11, 1.947138e-11, 2.001323e-11, 1.988278e-11, 2.004457e-11, 
    1.996192e-11, 2.010366e-11, 1.997607e-11, 2.019739e-11, 2.024578e-11, 
    2.021271e-11, 2.033992e-11, 1.996901e-11, 2.011098e-11, 1.905754e-11, 
    1.906364e-11, 1.909208e-11, 1.896727e-11, 1.895965e-11, 1.884571e-11, 
    1.894707e-11, 1.899033e-11, 1.91004e-11, 1.916569e-11, 1.922786e-11, 
    1.936497e-11, 1.951878e-11, 1.973502e-11, 1.989122e-11, 1.999633e-11, 
    1.993184e-11, 1.998877e-11, 1.992514e-11, 1.989535e-11, 2.022765e-11, 
    2.004066e-11, 2.032159e-11, 2.030599e-11, 2.017862e-11, 2.030774e-11, 
    1.906793e-11, 1.903283e-11, 1.891128e-11, 1.900637e-11, 1.883332e-11, 
    1.893007e-11, 1.898584e-11, 1.920187e-11, 1.924953e-11, 1.929377e-11, 
    1.938134e-11, 1.949405e-11, 1.96927e-11, 1.986648e-11, 2.00259e-11, 
    2.00142e-11, 2.001832e-11, 2.005403e-11, 1.996565e-11, 2.006856e-11, 
    2.008586e-11, 2.004064e-11, 2.03039e-11, 2.022848e-11, 2.030565e-11, 
    2.025653e-11, 1.904424e-11, 1.910333e-11, 1.907139e-11, 1.913148e-11, 
    1.908913e-11, 1.927786e-11, 1.933466e-11, 1.960168e-11, 1.949183e-11, 
    1.966682e-11, 1.950957e-11, 1.953738e-11, 1.967256e-11, 1.951804e-11, 
    1.985688e-11, 1.96268e-11, 2.005541e-11, 1.982432e-11, 2.006995e-11, 
    2.002521e-11, 2.009931e-11, 2.016581e-11, 2.024966e-11, 2.04049e-11, 
    2.036889e-11, 2.049911e-11, 1.919162e-11, 1.926863e-11, 1.926184e-11, 
    1.934261e-11, 1.940246e-11, 1.953256e-11, 1.974228e-11, 1.966327e-11, 
    1.980846e-11, 1.983769e-11, 1.961715e-11, 1.975239e-11, 1.932027e-11, 
    1.938972e-11, 1.934835e-11, 1.919769e-11, 1.968146e-11, 1.943232e-11, 
    1.989381e-11, 1.975777e-11, 2.015632e-11, 1.995754e-11, 2.034908e-11, 
    2.051783e-11, 2.067737e-11, 2.086476e-11, 1.931074e-11, 1.925832e-11, 
    1.935222e-11, 1.948258e-11, 1.960398e-11, 1.976605e-11, 1.978268e-11, 
    1.981314e-11, 1.989218e-11, 1.995877e-11, 1.982279e-11, 1.997549e-11, 
    1.940585e-11, 1.970317e-11, 1.923853e-11, 1.937778e-11, 1.947489e-11, 
    1.943225e-11, 1.965425e-11, 1.970678e-11, 1.992111e-11, 1.981014e-11, 
    2.047611e-11, 2.017988e-11, 2.100809e-11, 2.077468e-11, 1.924003e-11, 
    1.931055e-11, 1.955716e-11, 1.94396e-11, 1.97769e-11, 1.986044e-11, 
    1.992851e-11, 2.001571e-11, 2.002514e-11, 2.007693e-11, 1.999211e-11, 
    2.007357e-11, 1.97664e-11, 1.990333e-11, 1.952888e-11, 1.961964e-11, 
    1.957786e-11, 1.953209e-11, 1.967355e-11, 1.982492e-11, 1.982816e-11, 
    1.987684e-11, 2.001442e-11, 1.977827e-11, 2.051453e-11, 2.0058e-11, 
    1.938763e-11, 1.952421e-11, 1.954375e-11, 1.949075e-11, 1.985206e-11, 
    1.97207e-11, 2.007566e-11, 1.997937e-11, 2.013729e-11, 2.005872e-11, 
    2.004718e-11, 1.994657e-11, 1.988408e-11, 1.972671e-11, 1.95992e-11, 
    1.949843e-11, 1.952184e-11, 1.963263e-11, 1.98342e-11, 2.002599e-11, 
    1.998389e-11, 2.012526e-11, 1.975233e-11, 1.990822e-11, 1.984788e-11, 
    2.000542e-11, 1.966117e-11, 1.995412e-11, 1.95867e-11, 1.961875e-11, 
    1.97181e-11, 1.991882e-11, 1.996338e-11, 2.001103e-11, 1.998162e-11, 
    1.983934e-11, 1.981608e-11, 1.971568e-11, 1.968801e-11, 1.961177e-11, 
    1.954878e-11, 1.960633e-11, 1.966687e-11, 1.983939e-11, 1.999562e-11, 
    2.016676e-11, 2.020877e-11, 2.041008e-11, 2.024613e-11, 2.05171e-11, 
    2.028661e-11, 2.068656e-11, 1.997116e-11, 2.027984e-11, 1.972262e-11, 
    1.978222e-11, 1.989028e-11, 2.01394e-11, 2.000468e-11, 2.016229e-11, 
    1.981517e-11, 1.963646e-11, 1.959037e-11, 1.950455e-11, 1.959233e-11, 
    1.958518e-11, 1.966937e-11, 1.96423e-11, 1.984514e-11, 1.973603e-11, 
    2.004689e-11, 2.016104e-11, 2.048544e-11, 2.068581e-11, 2.089093e-11, 
    2.098188e-11, 2.10096e-11, 2.10212e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
