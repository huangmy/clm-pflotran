netcdf ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-01-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 338 ;
	column = 338 ;
	pft = 5746 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "timestep fractional area burned for crop" ;
		BAF_CROP:units = "proportion" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "timestep fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "timestep fractional area burned" ;
		FAREA_BURNED:units = "proportion" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned in this timestep" ;
		LFC2:units = "per timestep" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "timestep fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/timestep" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 02/10/14 15:54:32" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "bandre" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c130821.nc" ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-01-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 10102 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "02/10/14" ;

 time_written =
  "15:54:32" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  4.726044e-14, 4.73878e-14, 4.736306e-14, 4.746568e-14, 4.740878e-14, 
    4.747595e-14, 4.728629e-14, 4.739284e-14, 4.732484e-14, 4.727194e-14, 
    4.766455e-14, 4.747026e-14, 4.786618e-14, 4.774249e-14, 4.805298e-14, 
    4.784692e-14, 4.809449e-14, 4.804707e-14, 4.818983e-14, 4.814895e-14, 
    4.833127e-14, 4.820869e-14, 4.842573e-14, 4.830203e-14, 4.832137e-14, 
    4.820464e-14, 4.750942e-14, 4.764037e-14, 4.750165e-14, 4.752034e-14, 
    4.751196e-14, 4.740994e-14, 4.735847e-14, 4.725073e-14, 4.72703e-14, 
    4.734945e-14, 4.752874e-14, 4.746793e-14, 4.76212e-14, 4.761774e-14, 
    4.77881e-14, 4.771132e-14, 4.799731e-14, 4.791613e-14, 4.815066e-14, 
    4.809171e-14, 4.814788e-14, 4.813086e-14, 4.814811e-14, 4.806164e-14, 
    4.809869e-14, 4.802259e-14, 4.77257e-14, 4.781302e-14, 4.755236e-14, 
    4.73953e-14, 4.729096e-14, 4.721684e-14, 4.722731e-14, 4.724729e-14, 
    4.734991e-14, 4.744636e-14, 4.751979e-14, 4.756888e-14, 4.761724e-14, 
    4.776339e-14, 4.784075e-14, 4.801371e-14, 4.798254e-14, 4.803536e-14, 
    4.808584e-14, 4.817051e-14, 4.815658e-14, 4.819386e-14, 4.803399e-14, 
    4.814025e-14, 4.796478e-14, 4.80128e-14, 4.763025e-14, 4.748435e-14, 
    4.742217e-14, 4.736781e-14, 4.723537e-14, 4.732684e-14, 4.729079e-14, 
    4.737657e-14, 4.743102e-14, 4.74041e-14, 4.757022e-14, 4.750566e-14, 
    4.784534e-14, 4.769915e-14, 4.807996e-14, 4.798894e-14, 4.810177e-14, 
    4.804421e-14, 4.81428e-14, 4.805408e-14, 4.820774e-14, 4.824116e-14, 
    4.821832e-14, 4.830607e-14, 4.804915e-14, 4.814787e-14, 4.740334e-14, 
    4.740773e-14, 4.74282e-14, 4.733819e-14, 4.733269e-14, 4.725018e-14, 
    4.732361e-14, 4.735486e-14, 4.743419e-14, 4.748107e-14, 4.752562e-14, 
    4.762352e-14, 4.773274e-14, 4.788534e-14, 4.799484e-14, 4.80682e-14, 
    4.802323e-14, 4.806293e-14, 4.801855e-14, 4.799774e-14, 4.822863e-14, 
    4.809903e-14, 4.829345e-14, 4.828271e-14, 4.819474e-14, 4.828392e-14, 
    4.741081e-14, 4.738554e-14, 4.729771e-14, 4.736645e-14, 4.72412e-14, 
    4.731131e-14, 4.735159e-14, 4.750698e-14, 4.754113e-14, 4.757274e-14, 
    4.763518e-14, 4.771525e-14, 4.785557e-14, 4.797753e-14, 4.808878e-14, 
    4.808064e-14, 4.808351e-14, 4.810833e-14, 4.804681e-14, 4.811843e-14, 
    4.813044e-14, 4.809903e-14, 4.828127e-14, 4.822924e-14, 4.828248e-14, 
    4.824861e-14, 4.739376e-14, 4.743628e-14, 4.741331e-14, 4.745651e-14, 
    4.742606e-14, 4.756134e-14, 4.760187e-14, 4.779137e-14, 4.771367e-14, 
    4.783734e-14, 4.772625e-14, 4.774593e-14, 4.784132e-14, 4.773226e-14, 
    4.797078e-14, 4.780908e-14, 4.81093e-14, 4.794797e-14, 4.81194e-14, 
    4.80883e-14, 4.81398e-14, 4.818588e-14, 4.824386e-14, 4.835071e-14, 
    4.832598e-14, 4.841531e-14, 4.749967e-14, 4.755476e-14, 4.754994e-14, 
    4.760759e-14, 4.76502e-14, 4.774254e-14, 4.789046e-14, 4.783487e-14, 
    4.793694e-14, 4.795738e-14, 4.780235e-14, 4.789755e-14, 4.759164e-14, 
    4.76411e-14, 4.761167e-14, 4.7504e-14, 4.784765e-14, 4.76714e-14, 
    4.799665e-14, 4.790135e-14, 4.817931e-14, 4.804112e-14, 4.831236e-14, 
    4.842806e-14, 4.853695e-14, 4.866394e-14, 4.758485e-14, 4.754742e-14, 
    4.761445e-14, 4.770708e-14, 4.779303e-14, 4.790716e-14, 4.791885e-14, 
    4.794021e-14, 4.799552e-14, 4.804202e-14, 4.794694e-14, 4.805368e-14, 
    4.765251e-14, 4.786295e-14, 4.753325e-14, 4.763259e-14, 4.770163e-14, 
    4.767138e-14, 4.782852e-14, 4.786551e-14, 4.801571e-14, 4.793812e-14, 
    4.839949e-14, 4.819558e-14, 4.876061e-14, 4.860298e-14, 4.753434e-14, 
    4.758473e-14, 4.775992e-14, 4.76766e-14, 4.791479e-14, 4.797331e-14, 
    4.80209e-14, 4.808167e-14, 4.808825e-14, 4.812424e-14, 4.806525e-14, 
    4.812192e-14, 4.79074e-14, 4.800331e-14, 4.773994e-14, 4.780409e-14, 
    4.777459e-14, 4.774221e-14, 4.784212e-14, 4.79484e-14, 4.795071e-14, 
    4.798477e-14, 4.808063e-14, 4.791576e-14, 4.842571e-14, 4.811095e-14, 
    4.763966e-14, 4.773657e-14, 4.775045e-14, 4.771292e-14, 4.796744e-14, 
    4.787529e-14, 4.812337e-14, 4.805638e-14, 4.816614e-14, 4.81116e-14, 
    4.810358e-14, 4.803351e-14, 4.798985e-14, 4.787951e-14, 4.778965e-14, 
    4.771837e-14, 4.773495e-14, 4.781324e-14, 4.795491e-14, 4.808883e-14, 
    4.80595e-14, 4.81578e-14, 4.789753e-14, 4.80067e-14, 4.79645e-14, 
    4.807452e-14, 4.783338e-14, 4.803863e-14, 4.778084e-14, 4.780347e-14, 
    4.787346e-14, 4.801408e-14, 4.804523e-14, 4.807841e-14, 4.805795e-14, 
    4.795851e-14, 4.794226e-14, 4.787177e-14, 4.785228e-14, 4.779855e-14, 
    4.775402e-14, 4.779469e-14, 4.783738e-14, 4.795857e-14, 4.806768e-14, 
    4.818653e-14, 4.821562e-14, 4.835419e-14, 4.824134e-14, 4.842745e-14, 
    4.826916e-14, 4.854308e-14, 4.805057e-14, 4.826458e-14, 4.787666e-14, 
    4.791852e-14, 4.799414e-14, 4.816754e-14, 4.8074e-14, 4.81834e-14, 
    4.794162e-14, 4.781592e-14, 4.778343e-14, 4.77227e-14, 4.778481e-14, 
    4.777977e-14, 4.783918e-14, 4.782009e-14, 4.796259e-14, 4.788608e-14, 
    4.810336e-14, 4.818255e-14, 4.840594e-14, 4.854264e-14, 4.868169e-14, 
    4.8743e-14, 4.876165e-14, 4.876945e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -1.76574e-14, -1.768033e-14, -1.767586e-14, -1.769436e-14, -1.768408e-14, 
    -1.76962e-14, -1.766203e-14, -1.768127e-14, -1.766897e-14, -1.765943e-14, 
    -1.773024e-14, -1.769518e-14, -1.776626e-14, -1.774404e-14, 
    -1.779968e-14, -1.776284e-14, -1.780707e-14, -1.779855e-14, 
    -1.782402e-14, -1.781673e-14, -1.784937e-14, -1.782739e-14, 
    -1.786615e-14, -1.784409e-14, -1.784757e-14, -1.782667e-14, 
    -1.770218e-14, -1.772591e-14, -1.770079e-14, -1.770417e-14, 
    -1.770264e-14, -1.768431e-14, -1.767511e-14, -1.765561e-14, 
    -1.765914e-14, -1.767344e-14, -1.770569e-14, -1.769471e-14, 
    -1.772223e-14, -1.772161e-14, -1.77522e-14, -1.773843e-14, -1.778965e-14, 
    -1.77751e-14, -1.781703e-14, -1.780651e-14, -1.781655e-14, -1.78135e-14, 
    -1.781659e-14, -1.780115e-14, -1.780777e-14, -1.779416e-14, 
    -1.774102e-14, -1.775669e-14, -1.770992e-14, -1.768178e-14, 
    -1.766288e-14, -1.764951e-14, -1.76514e-14, -1.765502e-14, -1.767352e-14, 
    -1.769083e-14, -1.770402e-14, -1.771285e-14, -1.772153e-14, 
    -1.774791e-14, -1.77617e-14, -1.779263e-14, -1.7787e-14, -1.779649e-14, 
    -1.780546e-14, -1.782059e-14, -1.78181e-14, -1.782477e-14, -1.779619e-14, 
    -1.781522e-14, -1.77838e-14, -1.779241e-14, -1.772411e-14, -1.769766e-14, 
    -1.76866e-14, -1.767673e-14, -1.765286e-14, -1.766936e-14, -1.766286e-14, 
    -1.767827e-14, -1.768808e-14, -1.768322e-14, -1.771309e-14, 
    -1.770149e-14, -1.776252e-14, -1.773628e-14, -1.780442e-14, 
    -1.778815e-14, -1.780831e-14, -1.779801e-14, -1.781566e-14, 
    -1.779978e-14, -1.782723e-14, -1.783323e-14, -1.782914e-14, 
    -1.784477e-14, -1.77989e-14, -1.781657e-14, -1.768309e-14, -1.768388e-14, 
    -1.768756e-14, -1.767141e-14, -1.767041e-14, -1.765552e-14, 
    -1.766875e-14, -1.767439e-14, -1.768863e-14, -1.769708e-14, 
    -1.770509e-14, -1.772268e-14, -1.774232e-14, -1.776965e-14, -1.77892e-14, 
    -1.78023e-14, -1.779426e-14, -1.780136e-14, -1.779343e-14, -1.77897e-14, 
    -1.7831e-14, -1.780785e-14, -1.784252e-14, -1.78406e-14, -1.782494e-14, 
    -1.784081e-14, -1.768444e-14, -1.767988e-14, -1.766409e-14, 
    -1.767645e-14, -1.765389e-14, -1.766655e-14, -1.767384e-14, 
    -1.770178e-14, -1.770786e-14, -1.771356e-14, -1.772476e-14, 
    -1.773913e-14, -1.776431e-14, -1.778613e-14, -1.780598e-14, 
    -1.780452e-14, -1.780503e-14, -1.780949e-14, -1.779849e-14, 
    -1.781129e-14, -1.781346e-14, -1.780782e-14, -1.784034e-14, 
    -1.783106e-14, -1.784056e-14, -1.783451e-14, -1.768135e-14, 
    -1.768902e-14, -1.768488e-14, -1.769267e-14, -1.76872e-14, -1.771157e-14, 
    -1.771886e-14, -1.775285e-14, -1.773886e-14, -1.776106e-14, -1.77411e-14, 
    -1.774465e-14, -1.776187e-14, -1.774217e-14, -1.778497e-14, 
    -1.775606e-14, -1.780966e-14, -1.778094e-14, -1.781146e-14, 
    -1.780589e-14, -1.781509e-14, -1.782334e-14, -1.783367e-14, 
    -1.785277e-14, -1.784834e-14, -1.786425e-14, -1.770041e-14, 
    -1.771036e-14, -1.770944e-14, -1.77198e-14, -1.772747e-14, -1.774401e-14, 
    -1.777054e-14, -1.776056e-14, -1.777882e-14, -1.77825e-14, -1.775472e-14, 
    -1.777183e-14, -1.771697e-14, -1.77259e-14, -1.772055e-14, -1.770122e-14, 
    -1.776292e-14, -1.773133e-14, -1.778954e-14, -1.777247e-14, 
    -1.782217e-14, -1.779753e-14, -1.784591e-14, -1.786663e-14, 
    -1.788589e-14, -1.790857e-14, -1.771573e-14, -1.770899e-14, 
    -1.772102e-14, -1.773773e-14, -1.775308e-14, -1.777352e-14, 
    -1.777559e-14, -1.777942e-14, -1.778931e-14, -1.779762e-14, 
    -1.778068e-14, -1.77997e-14, -1.772805e-14, -1.776563e-14, -1.770647e-14, 
    -1.772438e-14, -1.773673e-14, -1.773127e-14, -1.775941e-14, 
    -1.776604e-14, -1.779297e-14, -1.777903e-14, -1.786156e-14, 
    -1.782514e-14, -1.792566e-14, -1.789771e-14, -1.770664e-14, 
    -1.771569e-14, -1.774718e-14, -1.77322e-14, -1.777486e-14, -1.778536e-14, 
    -1.779384e-14, -1.780474e-14, -1.780589e-14, -1.781234e-14, 
    -1.780177e-14, -1.78119e-14, -1.777357e-14, -1.779071e-14, -1.774353e-14, 
    -1.775506e-14, -1.774975e-14, -1.774394e-14, -1.776185e-14, 
    -1.778096e-14, -1.77813e-14, -1.778743e-14, -1.780481e-14, -1.777503e-14, 
    -1.786637e-14, -1.781019e-14, -1.772555e-14, -1.774303e-14, 
    -1.774544e-14, -1.773869e-14, -1.778431e-14, -1.776781e-14, 
    -1.781217e-14, -1.780019e-14, -1.781979e-14, -1.781006e-14, 
    -1.780863e-14, -1.77961e-14, -1.778831e-14, -1.776858e-14, -1.775248e-14, 
    -1.773966e-14, -1.774264e-14, -1.775672e-14, -1.778211e-14, 
    -1.780602e-14, -1.78008e-14, -1.781831e-14, -1.777178e-14, -1.779135e-14, 
    -1.778381e-14, -1.780344e-14, -1.776031e-14, -1.779726e-14, 
    -1.775086e-14, -1.775493e-14, -1.776748e-14, -1.779272e-14, -1.77982e-14, 
    -1.780416e-14, -1.780047e-14, -1.778274e-14, -1.77798e-14, -1.776716e-14, 
    -1.77637e-14, -1.775404e-14, -1.774606e-14, -1.775337e-14, -1.776105e-14, 
    -1.778272e-14, -1.780225e-14, -1.782347e-14, -1.782863e-14, 
    -1.785352e-14, -1.783335e-14, -1.78667e-14, -1.78385e-14, -1.788719e-14, 
    -1.779929e-14, -1.783753e-14, -1.776803e-14, -1.777553e-14, 
    -1.778914e-14, -1.782015e-14, -1.780335e-14, -1.782296e-14, 
    -1.777968e-14, -1.775723e-14, -1.775133e-14, -1.774046e-14, 
    -1.775158e-14, -1.775067e-14, -1.776132e-14, -1.775789e-14, 
    -1.778344e-14, -1.776972e-14, -1.780862e-14, -1.782279e-14, 
    -1.786261e-14, -1.788698e-14, -1.791162e-14, -1.792251e-14, 
    -1.792581e-14, -1.79272e-14 ;

 CH4_SURF_DIFF_UNSAT =
  1.390431e-11, 1.377575e-11, 1.380085e-11, 1.369636e-11, 1.375444e-11, 
    1.368585e-11, 1.387836e-11, 1.377062e-11, 1.383951e-11, 1.389279e-11, 
    1.349103e-11, 1.369168e-11, 1.320386e-11, 1.332195e-11, 1.302103e-11, 
    1.322238e-11, 1.297968e-11, 1.302692e-11, 1.288376e-11, 1.292507e-11, 
    1.273885e-11, 1.286462e-11, 1.264053e-11, 1.276907e-11, 1.27491e-11, 
    1.286873e-11, 1.365155e-11, 1.351619e-11, 1.365953e-11, 1.364033e-11, 
    1.364895e-11, 1.375324e-11, 1.380546e-11, 1.391408e-11, 1.389443e-11, 
    1.381462e-11, 1.363168e-11, 1.369409e-11, 1.353621e-11, 1.35398e-11, 
    1.327869e-11, 1.335134e-11, 1.307609e-11, 1.315555e-11, 1.292335e-11, 
    1.298249e-11, 1.292614e-11, 1.294327e-11, 1.292592e-11, 1.301245e-11, 
    1.297551e-11, 1.305117e-11, 1.33378e-11, 1.325491e-11, 1.360737e-11, 
    1.376808e-11, 1.387366e-11, 1.3948e-11, 1.393752e-11, 1.391751e-11, 
    1.381415e-11, 1.371614e-11, 1.364091e-11, 1.359034e-11, 1.354031e-11, 
    1.330211e-11, 1.322832e-11, 1.305991e-11, 1.309063e-11, 1.303851e-11, 
    1.298835e-11, 1.290331e-11, 1.291738e-11, 1.287966e-11, 1.303989e-11, 
    1.293381e-11, 1.310806e-11, 1.306084e-11, 1.352668e-11, 1.367728e-11, 
    1.374075e-11, 1.379603e-11, 1.392945e-11, 1.383748e-11, 1.387382e-11, 
    1.378717e-11, 1.373178e-11, 1.375921e-11, 1.358896e-11, 1.365542e-11, 
    1.322392e-11, 1.336276e-11, 1.299422e-11, 1.308433e-11, 1.297244e-11, 
    1.302977e-11, 1.293125e-11, 1.301998e-11, 1.286557e-11, 1.283151e-11, 
    1.285481e-11, 1.276493e-11, 1.302486e-11, 1.292614e-11, 1.375997e-11, 
    1.375551e-11, 1.373467e-11, 1.382601e-11, 1.383157e-11, 1.391462e-11, 
    1.384075e-11, 1.380915e-11, 1.372856e-11, 1.368064e-11, 1.363491e-11, 
    1.353378e-11, 1.333115e-11, 1.318537e-11, 1.307853e-11, 1.300594e-11, 
    1.305054e-11, 1.301118e-11, 1.305517e-11, 1.307569e-11, 1.28443e-11, 
    1.297516e-11, 1.277793e-11, 1.278898e-11, 1.287876e-11, 1.278773e-11, 
    1.375237e-11, 1.377807e-11, 1.386686e-11, 1.379743e-11, 1.392363e-11, 
    1.385315e-11, 1.381244e-11, 1.365404e-11, 1.361896e-11, 1.358635e-11, 
    1.352168e-11, 1.334765e-11, 1.321409e-11, 1.309554e-11, 1.298542e-11, 
    1.299355e-11, 1.299068e-11, 1.296586e-11, 1.302719e-11, 1.295574e-11, 
    1.294368e-11, 1.297518e-11, 1.279046e-11, 1.28437e-11, 1.278921e-11, 
    1.282393e-11, 1.376972e-11, 1.372642e-11, 1.374983e-11, 1.370576e-11, 
    1.373683e-11, 1.359808e-11, 1.355618e-11, 1.327556e-11, 1.334913e-11, 
    1.323161e-11, 1.333729e-11, 1.33187e-11, 1.322774e-11, 1.333163e-11, 
    1.310213e-11, 1.325864e-11, 1.296489e-11, 1.312445e-11, 1.295477e-11, 
    1.29859e-11, 1.293429e-11, 1.288775e-11, 1.282878e-11, 1.271875e-11, 
    1.274436e-11, 1.265146e-11, 1.366158e-11, 1.360488e-11, 1.360988e-11, 
    1.35503e-11, 1.350606e-11, 1.332192e-11, 1.318043e-11, 1.323401e-11, 
    1.313529e-11, 1.311528e-11, 1.326513e-11, 1.317355e-11, 1.35668e-11, 
    1.35155e-11, 1.354607e-11, 1.365711e-11, 1.322171e-11, 1.348397e-11, 
    1.307675e-11, 1.316988e-11, 1.28944e-11, 1.30328e-11, 1.275843e-11, 
    1.263805e-11, 1.252315e-11, 1.238698e-11, 1.357383e-11, 1.361248e-11, 
    1.35432e-11, 1.33553e-11, 1.3274e-11, 1.316424e-11, 1.31529e-11, 
    1.313209e-11, 1.307787e-11, 1.303194e-11, 1.31255e-11, 1.302038e-11, 
    1.350357e-11, 1.320699e-11, 1.362706e-11, 1.352433e-11, 1.336042e-11, 
    1.348402e-11, 1.324011e-11, 1.320454e-11, 1.305795e-11, 1.313414e-11, 
    1.266793e-11, 1.287788e-11, 1.228201e-11, 1.24526e-11, 1.362595e-11, 
    1.357397e-11, 1.330545e-11, 1.347858e-11, 1.315684e-11, 1.309968e-11, 
    1.305284e-11, 1.29925e-11, 1.298595e-11, 1.294991e-11, 1.300887e-11, 
    1.295225e-11, 1.3164e-11, 1.30702e-11, 1.332438e-11, 1.326346e-11, 
    1.329156e-11, 1.332224e-11, 1.322706e-11, 1.312403e-11, 1.312181e-11, 
    1.308842e-11, 1.299341e-11, 1.315591e-11, 1.264043e-11, 1.296312e-11, 
    1.351704e-11, 1.332752e-11, 1.331443e-11, 1.334985e-11, 1.310544e-11, 
    1.31951e-11, 1.295079e-11, 1.301769e-11, 1.290774e-11, 1.296259e-11, 
    1.297063e-11, 1.304037e-11, 1.308344e-11, 1.319101e-11, 1.327722e-11, 
    1.334473e-11, 1.33291e-11, 1.325471e-11, 1.311768e-11, 1.298536e-11, 
    1.301456e-11, 1.291615e-11, 1.317359e-11, 1.306683e-11, 1.31083e-11, 
    1.299964e-11, 1.323543e-11, 1.303518e-11, 1.328562e-11, 1.326406e-11, 
    1.319686e-11, 1.305953e-11, 1.302876e-11, 1.299575e-11, 1.301613e-11, 
    1.311416e-11, 1.313008e-11, 1.31985e-11, 1.321727e-11, 1.326876e-11, 
    1.331106e-11, 1.327242e-11, 1.323158e-11, 1.311412e-11, 1.300644e-11, 
    1.288709e-11, 1.285757e-11, 1.271507e-11, 1.283128e-11, 1.26386e-11, 
    1.280272e-11, 1.251652e-11, 1.302338e-11, 1.280749e-11, 1.319379e-11, 
    1.315322e-11, 1.307919e-11, 1.290627e-11, 1.300015e-11, 1.289023e-11, 
    1.313071e-11, 1.325213e-11, 1.328316e-11, 1.334064e-11, 1.328184e-11, 
    1.328664e-11, 1.322988e-11, 1.324818e-11, 1.311018e-11, 1.318468e-11, 
    1.297083e-11, 1.28911e-11, 1.266125e-11, 1.251705e-11, 1.236785e-11, 
    1.230125e-11, 1.22809e-11, 1.227237e-11 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  2.007731e-23, 2.007729e-23, 2.00773e-23, 2.007729e-23, 2.007729e-23, 
    2.007729e-23, 2.00773e-23, 2.007729e-23, 2.00773e-23, 2.00773e-23, 
    2.007727e-23, 2.007729e-23, 2.007726e-23, 2.007727e-23, 2.007724e-23, 
    2.007726e-23, 2.007724e-23, 2.007724e-23, 2.007723e-23, 2.007723e-23, 
    2.007722e-23, 2.007723e-23, 2.007721e-23, 2.007722e-23, 2.007722e-23, 
    2.007723e-23, 2.007728e-23, 2.007728e-23, 2.007729e-23, 2.007728e-23, 
    2.007728e-23, 2.007729e-23, 2.00773e-23, 2.007731e-23, 2.00773e-23, 
    2.00773e-23, 2.007728e-23, 2.007729e-23, 2.007728e-23, 2.007728e-23, 
    2.007726e-23, 2.007727e-23, 2.007725e-23, 2.007725e-23, 2.007723e-23, 
    2.007724e-23, 2.007723e-23, 2.007724e-23, 2.007723e-23, 2.007724e-23, 
    2.007724e-23, 2.007725e-23, 2.007727e-23, 2.007726e-23, 2.007728e-23, 
    2.007729e-23, 2.00773e-23, 2.007731e-23, 2.007731e-23, 2.007731e-23, 
    2.00773e-23, 2.007729e-23, 2.007728e-23, 2.007728e-23, 2.007728e-23, 
    2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007723e-23, 2.007723e-23, 2.007723e-23, 2.007724e-23, 
    2.007724e-23, 2.007725e-23, 2.007725e-23, 2.007728e-23, 2.007729e-23, 
    2.007729e-23, 2.00773e-23, 2.007731e-23, 2.00773e-23, 2.00773e-23, 
    2.00773e-23, 2.007729e-23, 2.007729e-23, 2.007728e-23, 2.007728e-23, 
    2.007726e-23, 2.007727e-23, 2.007724e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007724e-23, 2.007723e-23, 2.007723e-23, 
    2.007723e-23, 2.007722e-23, 2.007724e-23, 2.007723e-23, 2.007729e-23, 
    2.007729e-23, 2.007729e-23, 2.00773e-23, 2.00773e-23, 2.007731e-23, 
    2.00773e-23, 2.00773e-23, 2.007729e-23, 2.007729e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007725e-23, 2.007725e-23, 2.007724e-23, 
    2.007725e-23, 2.007724e-23, 2.007725e-23, 2.007725e-23, 2.007723e-23, 
    2.007724e-23, 2.007722e-23, 2.007722e-23, 2.007723e-23, 2.007722e-23, 
    2.007729e-23, 2.007729e-23, 2.00773e-23, 2.00773e-23, 2.007731e-23, 
    2.00773e-23, 2.00773e-23, 2.007728e-23, 2.007728e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007722e-23, 2.007723e-23, 2.007722e-23, 
    2.007723e-23, 2.007729e-23, 2.007729e-23, 2.007729e-23, 2.007729e-23, 
    2.007729e-23, 2.007728e-23, 2.007728e-23, 2.007726e-23, 2.007727e-23, 
    2.007726e-23, 2.007727e-23, 2.007727e-23, 2.007726e-23, 2.007727e-23, 
    2.007725e-23, 2.007726e-23, 2.007724e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007723e-23, 2.007723e-23, 2.007722e-23, 
    2.007722e-23, 2.007721e-23, 2.007729e-23, 2.007728e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007727e-23, 2.007725e-23, 2.007726e-23, 
    2.007725e-23, 2.007725e-23, 2.007726e-23, 2.007725e-23, 2.007728e-23, 
    2.007728e-23, 2.007728e-23, 2.007728e-23, 2.007726e-23, 2.007727e-23, 
    2.007725e-23, 2.007725e-23, 2.007723e-23, 2.007724e-23, 2.007722e-23, 
    2.007721e-23, 2.00772e-23, 2.007719e-23, 2.007728e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 
    2.007725e-23, 2.007725e-23, 2.007724e-23, 2.007725e-23, 2.007724e-23, 
    2.007727e-23, 2.007726e-23, 2.007728e-23, 2.007728e-23, 2.007727e-23, 
    2.007727e-23, 2.007726e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 
    2.007722e-23, 2.007723e-23, 2.007719e-23, 2.00772e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007727e-23, 2.007725e-23, 2.007725e-23, 
    2.007725e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 
    2.007724e-23, 2.007725e-23, 2.007725e-23, 2.007727e-23, 2.007726e-23, 
    2.007726e-23, 2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 
    2.007725e-23, 2.007724e-23, 2.007725e-23, 2.007721e-23, 2.007724e-23, 
    2.007728e-23, 2.007727e-23, 2.007727e-23, 2.007727e-23, 2.007725e-23, 
    2.007726e-23, 2.007724e-23, 2.007724e-23, 2.007723e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007725e-23, 2.007726e-23, 2.007726e-23, 
    2.007727e-23, 2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007723e-23, 2.007725e-23, 2.007725e-23, 2.007725e-23, 
    2.007724e-23, 2.007726e-23, 2.007724e-23, 2.007726e-23, 2.007726e-23, 
    2.007726e-23, 2.007725e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 
    2.007725e-23, 2.007725e-23, 2.007726e-23, 2.007726e-23, 2.007726e-23, 
    2.007727e-23, 2.007726e-23, 2.007726e-23, 2.007725e-23, 2.007724e-23, 
    2.007723e-23, 2.007723e-23, 2.007722e-23, 2.007723e-23, 2.007721e-23, 
    2.007722e-23, 2.00772e-23, 2.007724e-23, 2.007722e-23, 2.007726e-23, 
    2.007725e-23, 2.007725e-23, 2.007723e-23, 2.007724e-23, 2.007723e-23, 
    2.007725e-23, 2.007726e-23, 2.007726e-23, 2.007727e-23, 2.007726e-23, 
    2.007726e-23, 2.007726e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 
    2.007724e-23, 2.007723e-23, 2.007721e-23, 2.00772e-23, 2.007719e-23, 
    2.007719e-23, 2.007719e-23, 2.007719e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  2.052861e-24, 2.05286e-24, 2.05286e-24, 2.052859e-24, 2.05286e-24, 
    2.052859e-24, 2.052861e-24, 2.05286e-24, 2.052861e-24, 2.052861e-24, 
    2.052857e-24, 2.052859e-24, 2.052855e-24, 2.052856e-24, 2.052853e-24, 
    2.052855e-24, 2.052852e-24, 2.052853e-24, 2.052851e-24, 2.052852e-24, 
    2.05285e-24, 2.052851e-24, 2.052848e-24, 2.05285e-24, 2.05285e-24, 
    2.052851e-24, 2.052859e-24, 2.052857e-24, 2.052859e-24, 2.052858e-24, 
    2.052858e-24, 2.05286e-24, 2.05286e-24, 2.052861e-24, 2.052861e-24, 
    2.05286e-24, 2.052858e-24, 2.052859e-24, 2.052857e-24, 2.052857e-24, 
    2.052855e-24, 2.052856e-24, 2.052853e-24, 2.052854e-24, 2.052852e-24, 
    2.052852e-24, 2.052852e-24, 2.052852e-24, 2.052852e-24, 2.052853e-24, 
    2.052852e-24, 2.052853e-24, 2.052856e-24, 2.052855e-24, 2.052858e-24, 
    2.05286e-24, 2.052861e-24, 2.052862e-24, 2.052862e-24, 2.052861e-24, 
    2.05286e-24, 2.052859e-24, 2.052858e-24, 2.052858e-24, 2.052857e-24, 
    2.052856e-24, 2.052855e-24, 2.052853e-24, 2.052853e-24, 2.052853e-24, 
    2.052852e-24, 2.052851e-24, 2.052851e-24, 2.052851e-24, 2.052853e-24, 
    2.052852e-24, 2.052854e-24, 2.052853e-24, 2.052857e-24, 2.052859e-24, 
    2.052859e-24, 2.05286e-24, 2.052862e-24, 2.052861e-24, 2.052861e-24, 
    2.05286e-24, 2.052859e-24, 2.05286e-24, 2.052858e-24, 2.052859e-24, 
    2.052855e-24, 2.052856e-24, 2.052852e-24, 2.052853e-24, 2.052852e-24, 
    2.052853e-24, 2.052852e-24, 2.052853e-24, 2.052851e-24, 2.052851e-24, 
    2.052851e-24, 2.05285e-24, 2.052853e-24, 2.052852e-24, 2.05286e-24, 
    2.05286e-24, 2.052859e-24, 2.05286e-24, 2.05286e-24, 2.052861e-24, 
    2.052861e-24, 2.05286e-24, 2.052859e-24, 2.052859e-24, 2.052858e-24, 
    2.052857e-24, 2.052856e-24, 2.052855e-24, 2.052853e-24, 2.052852e-24, 
    2.052853e-24, 2.052853e-24, 2.052853e-24, 2.052853e-24, 2.052851e-24, 
    2.052852e-24, 2.05285e-24, 2.05285e-24, 2.052851e-24, 2.05285e-24, 
    2.05286e-24, 2.05286e-24, 2.052861e-24, 2.05286e-24, 2.052861e-24, 
    2.052861e-24, 2.05286e-24, 2.052859e-24, 2.052858e-24, 2.052858e-24, 
    2.052857e-24, 2.052856e-24, 2.052855e-24, 2.052853e-24, 2.052852e-24, 
    2.052852e-24, 2.052852e-24, 2.052852e-24, 2.052853e-24, 2.052852e-24, 
    2.052852e-24, 2.052852e-24, 2.05285e-24, 2.052851e-24, 2.05285e-24, 
    2.05285e-24, 2.05286e-24, 2.052859e-24, 2.05286e-24, 2.052859e-24, 
    2.052859e-24, 2.052858e-24, 2.052857e-24, 2.052855e-24, 2.052856e-24, 
    2.052855e-24, 2.052856e-24, 2.052856e-24, 2.052855e-24, 2.052856e-24, 
    2.052854e-24, 2.052855e-24, 2.052852e-24, 2.052854e-24, 2.052852e-24, 
    2.052852e-24, 2.052852e-24, 2.052851e-24, 2.05285e-24, 2.052849e-24, 
    2.05285e-24, 2.052849e-24, 2.052859e-24, 2.052858e-24, 2.052858e-24, 
    2.052857e-24, 2.052857e-24, 2.052856e-24, 2.052854e-24, 2.052855e-24, 
    2.052854e-24, 2.052854e-24, 2.052855e-24, 2.052854e-24, 2.052858e-24, 
    2.052857e-24, 2.052857e-24, 2.052859e-24, 2.052855e-24, 2.052857e-24, 
    2.052853e-24, 2.052854e-24, 2.052851e-24, 2.052853e-24, 2.05285e-24, 
    2.052848e-24, 2.052847e-24, 2.052846e-24, 2.052858e-24, 2.052858e-24, 
    2.052857e-24, 2.052856e-24, 2.052855e-24, 2.052854e-24, 2.052854e-24, 
    2.052854e-24, 2.052853e-24, 2.052853e-24, 2.052854e-24, 2.052853e-24, 
    2.052857e-24, 2.052855e-24, 2.052858e-24, 2.052857e-24, 2.052856e-24, 
    2.052857e-24, 2.052855e-24, 2.052855e-24, 2.052853e-24, 2.052854e-24, 
    2.052849e-24, 2.052851e-24, 2.052845e-24, 2.052846e-24, 2.052858e-24, 
    2.052858e-24, 2.052856e-24, 2.052857e-24, 2.052854e-24, 2.052854e-24, 
    2.052853e-24, 2.052852e-24, 2.052852e-24, 2.052852e-24, 2.052852e-24, 
    2.052852e-24, 2.052854e-24, 2.052853e-24, 2.052856e-24, 2.052855e-24, 
    2.052856e-24, 2.052856e-24, 2.052855e-24, 2.052854e-24, 2.052854e-24, 
    2.052853e-24, 2.052852e-24, 2.052854e-24, 2.052848e-24, 2.052852e-24, 
    2.052857e-24, 2.052856e-24, 2.052856e-24, 2.052856e-24, 2.052854e-24, 
    2.052855e-24, 2.052852e-24, 2.052853e-24, 2.052851e-24, 2.052852e-24, 
    2.052852e-24, 2.052853e-24, 2.052853e-24, 2.052855e-24, 2.052855e-24, 
    2.052856e-24, 2.052856e-24, 2.052855e-24, 2.052854e-24, 2.052852e-24, 
    2.052853e-24, 2.052851e-24, 2.052854e-24, 2.052853e-24, 2.052854e-24, 
    2.052852e-24, 2.052855e-24, 2.052853e-24, 2.052855e-24, 2.052855e-24, 
    2.052855e-24, 2.052853e-24, 2.052853e-24, 2.052852e-24, 2.052853e-24, 
    2.052854e-24, 2.052854e-24, 2.052855e-24, 2.052855e-24, 2.052855e-24, 
    2.052856e-24, 2.052855e-24, 2.052855e-24, 2.052854e-24, 2.052852e-24, 
    2.052851e-24, 2.052851e-24, 2.052849e-24, 2.052851e-24, 2.052848e-24, 
    2.05285e-24, 2.052847e-24, 2.052853e-24, 2.05285e-24, 2.052855e-24, 
    2.052854e-24, 2.052853e-24, 2.052851e-24, 2.052852e-24, 2.052851e-24, 
    2.052854e-24, 2.052855e-24, 2.052855e-24, 2.052856e-24, 2.052855e-24, 
    2.052855e-24, 2.052855e-24, 2.052855e-24, 2.052854e-24, 2.052855e-24, 
    2.052852e-24, 2.052851e-24, 2.052849e-24, 2.052847e-24, 2.052846e-24, 
    2.052845e-24, 2.052845e-24, 2.052845e-24 ;

 CONC_CH4_SAT =
  7.844502e-08, 7.855568e-08, 7.853413e-08, 7.862337e-08, 7.85738e-08, 
    7.863227e-08, 7.846737e-08, 7.856016e-08, 7.850088e-08, 7.845485e-08, 
    7.87964e-08, 7.862732e-08, 7.897037e-08, 7.886317e-08, 7.913169e-08, 
    7.895385e-08, 7.916742e-08, 7.912632e-08, 7.924933e-08, 7.92141e-08, 
    7.937157e-08, 7.926557e-08, 7.94526e-08, 7.934615e-08, 7.936291e-08, 
    7.926211e-08, 7.866116e-08, 7.877546e-08, 7.865444e-08, 7.867074e-08, 
    7.866337e-08, 7.857491e-08, 7.853042e-08, 7.843639e-08, 7.845343e-08, 
    7.852239e-08, 7.867806e-08, 7.862512e-08, 7.875798e-08, 7.875497e-08, 
    7.890261e-08, 7.88361e-08, 7.908339e-08, 7.901318e-08, 7.921557e-08, 
    7.916479e-08, 7.921323e-08, 7.919851e-08, 7.921342e-08, 7.913891e-08, 
    7.917086e-08, 7.910516e-08, 7.884861e-08, 7.892423e-08, 7.869847e-08, 
    7.856256e-08, 7.847149e-08, 7.840694e-08, 7.841607e-08, 7.843352e-08, 
    7.85228e-08, 7.86064e-08, 7.867007e-08, 7.871266e-08, 7.875455e-08, 
    7.888173e-08, 7.894839e-08, 7.909769e-08, 7.907057e-08, 7.911634e-08, 
    7.915973e-08, 7.923276e-08, 7.922071e-08, 7.925291e-08, 7.911498e-08, 
    7.920676e-08, 7.905517e-08, 7.909671e-08, 7.876675e-08, 7.863937e-08, 
    7.858583e-08, 7.85383e-08, 7.842311e-08, 7.850273e-08, 7.847137e-08, 
    7.854577e-08, 7.85931e-08, 7.856966e-08, 7.871382e-08, 7.865786e-08, 
    7.895234e-08, 7.882571e-08, 7.915467e-08, 7.907612e-08, 7.917345e-08, 
    7.912377e-08, 7.920892e-08, 7.913229e-08, 7.926482e-08, 7.929372e-08, 
    7.927399e-08, 7.934946e-08, 7.912806e-08, 7.921331e-08, 7.856904e-08, 
    7.857287e-08, 7.85906e-08, 7.851261e-08, 7.850779e-08, 7.843596e-08, 
    7.849981e-08, 7.852704e-08, 7.859578e-08, 7.863653e-08, 7.867519e-08, 
    7.876009e-08, 7.885484e-08, 7.898679e-08, 7.908123e-08, 7.914446e-08, 
    7.910565e-08, 7.913993e-08, 7.910163e-08, 7.908364e-08, 7.928295e-08, 
    7.917121e-08, 7.933861e-08, 7.932934e-08, 7.92537e-08, 7.933038e-08, 
    7.857555e-08, 7.855353e-08, 7.847732e-08, 7.853697e-08, 7.842812e-08, 
    7.848919e-08, 7.852432e-08, 7.865921e-08, 7.868859e-08, 7.871608e-08, 
    7.877014e-08, 7.883952e-08, 7.896103e-08, 7.906637e-08, 7.916221e-08, 
    7.915519e-08, 7.915767e-08, 7.917914e-08, 7.912605e-08, 7.918784e-08, 
    7.919828e-08, 7.91711e-08, 7.93281e-08, 7.928329e-08, 7.932914e-08, 
    7.929995e-08, 7.856067e-08, 7.859765e-08, 7.857768e-08, 7.861527e-08, 
    7.858885e-08, 7.870641e-08, 7.87416e-08, 7.890566e-08, 7.88382e-08, 
    7.894531e-08, 7.884903e-08, 7.886614e-08, 7.894914e-08, 7.885418e-08, 
    7.906073e-08, 7.89211e-08, 7.917997e-08, 7.904121e-08, 7.918867e-08, 
    7.91618e-08, 7.92062e-08, 7.924601e-08, 7.92959e-08, 7.938804e-08, 
    7.936669e-08, 7.944351e-08, 7.865265e-08, 7.870059e-08, 7.869622e-08, 
    7.874623e-08, 7.878322e-08, 7.88631e-08, 7.89911e-08, 7.894296e-08, 
    7.903114e-08, 7.904887e-08, 7.89148e-08, 7.899731e-08, 7.873253e-08, 
    7.877557e-08, 7.874984e-08, 7.865652e-08, 7.895427e-08, 7.88018e-08, 
    7.908282e-08, 7.900047e-08, 7.924036e-08, 7.912137e-08, 7.935497e-08, 
    7.945486e-08, 7.954796e-08, 7.965734e-08, 7.872656e-08, 7.869403e-08, 
    7.875213e-08, 7.883268e-08, 7.890685e-08, 7.900552e-08, 7.901552e-08, 
    7.903403e-08, 7.908174e-08, 7.912189e-08, 7.904003e-08, 7.913194e-08, 
    7.878585e-08, 7.896741e-08, 7.868186e-08, 7.876825e-08, 7.882787e-08, 
    7.880156e-08, 7.893741e-08, 7.896943e-08, 7.909937e-08, 7.903215e-08, 
    7.943036e-08, 7.925463e-08, 7.973993e-08, 7.960495e-08, 7.86827e-08, 
    7.872638e-08, 7.887832e-08, 7.880607e-08, 7.901203e-08, 7.906265e-08, 
    7.910364e-08, 7.915622e-08, 7.916179e-08, 7.919289e-08, 7.914193e-08, 
    7.919082e-08, 7.900574e-08, 7.908852e-08, 7.886079e-08, 7.891641e-08, 
    7.889078e-08, 7.886276e-08, 7.89492e-08, 7.904136e-08, 7.904308e-08, 
    7.907263e-08, 7.915625e-08, 7.901285e-08, 7.945344e-08, 7.918227e-08, 
    7.877399e-08, 7.885826e-08, 7.886999e-08, 7.883742e-08, 7.905759e-08, 
    7.897796e-08, 7.91921e-08, 7.913427e-08, 7.922892e-08, 7.918193e-08, 
    7.917502e-08, 7.911454e-08, 7.907691e-08, 7.898166e-08, 7.890395e-08, 
    7.884211e-08, 7.885648e-08, 7.892438e-08, 7.904693e-08, 7.91624e-08, 
    7.913717e-08, 7.922173e-08, 7.899713e-08, 7.909157e-08, 7.905517e-08, 
    7.914997e-08, 7.894173e-08, 7.911986e-08, 7.889618e-08, 7.891578e-08, 
    7.897638e-08, 7.909814e-08, 7.912466e-08, 7.915341e-08, 7.913562e-08, 
    7.904999e-08, 7.903584e-08, 7.897484e-08, 7.895812e-08, 7.89115e-08, 
    7.887299e-08, 7.890824e-08, 7.894528e-08, 7.904993e-08, 7.914417e-08, 
    7.924662e-08, 7.927155e-08, 7.939151e-08, 7.929422e-08, 7.9455e-08, 
    7.931886e-08, 7.955401e-08, 7.91298e-08, 7.931435e-08, 7.897905e-08, 
    7.901523e-08, 7.908086e-08, 7.923051e-08, 7.914952e-08, 7.924411e-08, 
    7.903526e-08, 7.892685e-08, 7.889845e-08, 7.884592e-08, 7.889965e-08, 
    7.889527e-08, 7.894663e-08, 7.893012e-08, 7.905339e-08, 7.898721e-08, 
    7.917492e-08, 7.92433e-08, 7.943555e-08, 7.955316e-08, 7.967216e-08, 
    7.972473e-08, 7.974069e-08, 7.974737e-08,
  2.101887e-10, 2.107804e-10, 2.106652e-10, 2.111435e-10, 2.108775e-10, 
    2.111915e-10, 2.103082e-10, 2.108044e-10, 2.104874e-10, 2.102413e-10, 
    2.120774e-10, 2.111648e-10, 2.130192e-10, 2.124389e-10, 2.138943e-10, 
    2.129296e-10, 2.140884e-10, 2.138653e-10, 2.145337e-10, 2.143423e-10, 
    2.151989e-10, 2.146221e-10, 2.156406e-10, 2.150606e-10, 2.151518e-10, 
    2.146032e-10, 2.113475e-10, 2.119642e-10, 2.113112e-10, 2.113991e-10, 
    2.113594e-10, 2.108833e-10, 2.106452e-10, 2.101427e-10, 2.102337e-10, 
    2.106024e-10, 2.114386e-10, 2.111531e-10, 2.118702e-10, 2.11854e-10, 
    2.126524e-10, 2.122925e-10, 2.136323e-10, 2.132515e-10, 2.143502e-10, 
    2.140742e-10, 2.143375e-10, 2.142575e-10, 2.143385e-10, 2.139336e-10, 
    2.141072e-10, 2.137505e-10, 2.123602e-10, 2.127694e-10, 2.115488e-10, 
    2.108171e-10, 2.103302e-10, 2.099854e-10, 2.100342e-10, 2.101273e-10, 
    2.106045e-10, 2.110521e-10, 2.113956e-10, 2.116254e-10, 2.118517e-10, 
    2.125391e-10, 2.129001e-10, 2.137098e-10, 2.135628e-10, 2.138111e-10, 
    2.140467e-10, 2.144436e-10, 2.143781e-10, 2.145532e-10, 2.138038e-10, 
    2.143023e-10, 2.134792e-10, 2.137046e-10, 2.119171e-10, 2.112299e-10, 
    2.109417e-10, 2.106875e-10, 2.100717e-10, 2.104972e-10, 2.103296e-10, 
    2.107275e-10, 2.109808e-10, 2.108553e-10, 2.116317e-10, 2.113296e-10, 
    2.129216e-10, 2.122362e-10, 2.140192e-10, 2.135929e-10, 2.141213e-10, 
    2.138515e-10, 2.14314e-10, 2.138977e-10, 2.14618e-10, 2.147751e-10, 
    2.146678e-10, 2.150786e-10, 2.138748e-10, 2.143378e-10, 2.10852e-10, 
    2.108725e-10, 2.109675e-10, 2.1055e-10, 2.105243e-10, 2.101404e-10, 
    2.104816e-10, 2.106272e-10, 2.109951e-10, 2.112146e-10, 2.114232e-10, 
    2.118816e-10, 2.123938e-10, 2.131083e-10, 2.136206e-10, 2.139639e-10, 
    2.137531e-10, 2.139392e-10, 2.137313e-10, 2.136337e-10, 2.147165e-10, 
    2.14109e-10, 2.150196e-10, 2.149691e-10, 2.145575e-10, 2.149748e-10, 
    2.108868e-10, 2.107691e-10, 2.103614e-10, 2.106805e-10, 2.100985e-10, 
    2.104248e-10, 2.106126e-10, 2.113368e-10, 2.114955e-10, 2.116439e-10, 
    2.119359e-10, 2.12311e-10, 2.129687e-10, 2.135399e-10, 2.140603e-10, 
    2.140221e-10, 2.140356e-10, 2.141522e-10, 2.138638e-10, 2.141995e-10, 
    2.142562e-10, 2.141085e-10, 2.149624e-10, 2.147185e-10, 2.14968e-10, 
    2.148091e-10, 2.108072e-10, 2.110052e-10, 2.108983e-10, 2.110999e-10, 
    2.10958e-10, 2.115915e-10, 2.117815e-10, 2.126688e-10, 2.123038e-10, 
    2.128835e-10, 2.123624e-10, 2.12455e-10, 2.129041e-10, 2.123903e-10, 
    2.135092e-10, 2.127523e-10, 2.141567e-10, 2.134032e-10, 2.14204e-10, 
    2.14058e-10, 2.142993e-10, 2.145157e-10, 2.147871e-10, 2.152887e-10, 
    2.151724e-10, 2.155911e-10, 2.113015e-10, 2.115602e-10, 2.115367e-10, 
    2.118067e-10, 2.120066e-10, 2.124386e-10, 2.131317e-10, 2.128709e-10, 
    2.133489e-10, 2.13445e-10, 2.127184e-10, 2.131654e-10, 2.117327e-10, 
    2.119651e-10, 2.118262e-10, 2.113224e-10, 2.12932e-10, 2.121068e-10, 
    2.136292e-10, 2.131825e-10, 2.144849e-10, 2.138383e-10, 2.151086e-10, 
    2.156528e-10, 2.16161e-10, 2.167584e-10, 2.117005e-10, 2.115249e-10, 
    2.118386e-10, 2.122739e-10, 2.126753e-10, 2.132099e-10, 2.132642e-10, 
    2.133645e-10, 2.136234e-10, 2.138413e-10, 2.133969e-10, 2.138958e-10, 
    2.120205e-10, 2.130033e-10, 2.114592e-10, 2.119255e-10, 2.122479e-10, 
    2.121057e-10, 2.128409e-10, 2.130143e-10, 2.137189e-10, 2.133543e-10, 
    2.155191e-10, 2.145624e-10, 2.172103e-10, 2.164721e-10, 2.114637e-10, 
    2.116995e-10, 2.125209e-10, 2.121301e-10, 2.132452e-10, 2.135197e-10, 
    2.137422e-10, 2.140277e-10, 2.140579e-10, 2.142269e-10, 2.139501e-10, 
    2.142157e-10, 2.132111e-10, 2.136601e-10, 2.124261e-10, 2.127271e-10, 
    2.125884e-10, 2.124368e-10, 2.129047e-10, 2.134041e-10, 2.134136e-10, 
    2.135739e-10, 2.140274e-10, 2.132497e-10, 2.156447e-10, 2.141688e-10, 
    2.119567e-10, 2.124122e-10, 2.124758e-10, 2.122997e-10, 2.134923e-10, 
    2.130605e-10, 2.142226e-10, 2.139085e-10, 2.144228e-10, 2.141674e-10, 
    2.141299e-10, 2.138014e-10, 2.135971e-10, 2.130806e-10, 2.126597e-10, 
    2.123251e-10, 2.124028e-10, 2.127702e-10, 2.134344e-10, 2.140612e-10, 
    2.139241e-10, 2.143837e-10, 2.131644e-10, 2.136766e-10, 2.134791e-10, 
    2.139937e-10, 2.128642e-10, 2.138298e-10, 2.126176e-10, 2.127238e-10, 
    2.13052e-10, 2.137121e-10, 2.138563e-10, 2.140124e-10, 2.139158e-10, 
    2.13451e-10, 2.133743e-10, 2.130437e-10, 2.12953e-10, 2.127006e-10, 
    2.124921e-10, 2.126829e-10, 2.128834e-10, 2.134507e-10, 2.139622e-10, 
    2.145189e-10, 2.146546e-10, 2.153074e-10, 2.147777e-10, 2.156532e-10, 
    2.149114e-10, 2.161936e-10, 2.13884e-10, 2.148872e-10, 2.130665e-10, 
    2.132626e-10, 2.136184e-10, 2.144313e-10, 2.139913e-10, 2.145052e-10, 
    2.133712e-10, 2.127835e-10, 2.126299e-10, 2.123456e-10, 2.126364e-10, 
    2.126127e-10, 2.128909e-10, 2.128014e-10, 2.134695e-10, 2.131107e-10, 
    2.141292e-10, 2.145008e-10, 2.155476e-10, 2.161892e-10, 2.168396e-10, 
    2.171271e-10, 2.172145e-10, 2.172511e-10,
  1.164426e-13, 1.168784e-13, 1.167935e-13, 1.171459e-13, 1.1695e-13, 
    1.171812e-13, 1.165306e-13, 1.16896e-13, 1.166626e-13, 1.164814e-13, 
    1.178336e-13, 1.171616e-13, 1.185286e-13, 1.181004e-13, 1.191781e-13, 
    1.184624e-13, 1.193254e-13, 1.191563e-13, 1.196635e-13, 1.195181e-13, 
    1.201685e-13, 1.197305e-13, 1.205045e-13, 1.200635e-13, 1.201328e-13, 
    1.197162e-13, 1.172961e-13, 1.177501e-13, 1.172694e-13, 1.173341e-13, 
    1.173049e-13, 1.169543e-13, 1.167787e-13, 1.164088e-13, 1.164758e-13, 
    1.167472e-13, 1.173632e-13, 1.17153e-13, 1.176812e-13, 1.176693e-13, 
    1.182579e-13, 1.179925e-13, 1.189816e-13, 1.187003e-13, 1.195242e-13, 
    1.193147e-13, 1.195145e-13, 1.194538e-13, 1.195152e-13, 1.192081e-13, 
    1.193397e-13, 1.190692e-13, 1.180424e-13, 1.183443e-13, 1.174443e-13, 
    1.169053e-13, 1.165468e-13, 1.16293e-13, 1.163289e-13, 1.163974e-13, 
    1.167488e-13, 1.170787e-13, 1.173316e-13, 1.175008e-13, 1.176676e-13, 
    1.181742e-13, 1.184407e-13, 1.190388e-13, 1.189302e-13, 1.191151e-13, 
    1.192939e-13, 1.19595e-13, 1.195453e-13, 1.196782e-13, 1.191096e-13, 
    1.194877e-13, 1.188686e-13, 1.190351e-13, 1.177154e-13, 1.172096e-13, 
    1.169971e-13, 1.168099e-13, 1.163565e-13, 1.166698e-13, 1.165463e-13, 
    1.168395e-13, 1.170261e-13, 1.169337e-13, 1.175055e-13, 1.17283e-13, 
    1.184565e-13, 1.17951e-13, 1.19273e-13, 1.189525e-13, 1.193504e-13, 
    1.191458e-13, 1.194966e-13, 1.191809e-13, 1.197274e-13, 1.198467e-13, 
    1.197652e-13, 1.200773e-13, 1.191635e-13, 1.195147e-13, 1.169312e-13, 
    1.169463e-13, 1.170163e-13, 1.167087e-13, 1.166897e-13, 1.164071e-13, 
    1.166583e-13, 1.167656e-13, 1.170368e-13, 1.171983e-13, 1.173519e-13, 
    1.176895e-13, 1.180671e-13, 1.185945e-13, 1.189729e-13, 1.192311e-13, 
    1.190712e-13, 1.192124e-13, 1.190548e-13, 1.189827e-13, 1.198022e-13, 
    1.193411e-13, 1.200324e-13, 1.199941e-13, 1.196814e-13, 1.199984e-13, 
    1.169569e-13, 1.168701e-13, 1.165698e-13, 1.168048e-13, 1.163763e-13, 
    1.166165e-13, 1.167548e-13, 1.172882e-13, 1.174052e-13, 1.175144e-13, 
    1.177296e-13, 1.180061e-13, 1.184914e-13, 1.189133e-13, 1.193042e-13, 
    1.192752e-13, 1.192854e-13, 1.193739e-13, 1.191552e-13, 1.194097e-13, 
    1.194527e-13, 1.193407e-13, 1.19989e-13, 1.198037e-13, 1.199933e-13, 
    1.198726e-13, 1.168983e-13, 1.170441e-13, 1.169653e-13, 1.171139e-13, 
    1.170093e-13, 1.174758e-13, 1.176157e-13, 1.1827e-13, 1.180008e-13, 
    1.184285e-13, 1.180441e-13, 1.181123e-13, 1.184435e-13, 1.180647e-13, 
    1.188905e-13, 1.183315e-13, 1.193773e-13, 1.188122e-13, 1.194132e-13, 
    1.193025e-13, 1.194855e-13, 1.196497e-13, 1.198558e-13, 1.202369e-13, 
    1.201486e-13, 1.204669e-13, 1.172623e-13, 1.174527e-13, 1.174355e-13, 
    1.176344e-13, 1.177817e-13, 1.181002e-13, 1.186118e-13, 1.184193e-13, 
    1.187722e-13, 1.188432e-13, 1.183067e-13, 1.186366e-13, 1.175798e-13, 
    1.17751e-13, 1.176487e-13, 1.172776e-13, 1.184643e-13, 1.178555e-13, 
    1.189793e-13, 1.186493e-13, 1.196264e-13, 1.191357e-13, 1.201001e-13, 
    1.205136e-13, 1.209006e-13, 1.213556e-13, 1.175561e-13, 1.174268e-13, 
    1.176579e-13, 1.179787e-13, 1.182749e-13, 1.186695e-13, 1.187097e-13, 
    1.187837e-13, 1.18975e-13, 1.191381e-13, 1.188076e-13, 1.191794e-13, 
    1.177917e-13, 1.185169e-13, 1.173783e-13, 1.177218e-13, 1.179595e-13, 
    1.178548e-13, 1.183971e-13, 1.185252e-13, 1.190456e-13, 1.187763e-13, 
    1.20412e-13, 1.196851e-13, 1.217003e-13, 1.211374e-13, 1.173817e-13, 
    1.175554e-13, 1.181609e-13, 1.178727e-13, 1.186956e-13, 1.188984e-13, 
    1.19063e-13, 1.192794e-13, 1.193024e-13, 1.194305e-13, 1.192206e-13, 
    1.194221e-13, 1.186704e-13, 1.190022e-13, 1.180911e-13, 1.183131e-13, 
    1.182108e-13, 1.180989e-13, 1.184442e-13, 1.188129e-13, 1.1882e-13, 
    1.189384e-13, 1.192787e-13, 1.18699e-13, 1.205073e-13, 1.19386e-13, 
    1.17745e-13, 1.180807e-13, 1.181277e-13, 1.179978e-13, 1.188781e-13, 
    1.185592e-13, 1.194273e-13, 1.19189e-13, 1.195792e-13, 1.193854e-13, 
    1.193569e-13, 1.191078e-13, 1.189556e-13, 1.18574e-13, 1.182633e-13, 
    1.180166e-13, 1.180739e-13, 1.183449e-13, 1.188353e-13, 1.193048e-13, 
    1.192008e-13, 1.195496e-13, 1.18636e-13, 1.190143e-13, 1.188683e-13, 
    1.192537e-13, 1.184143e-13, 1.19129e-13, 1.182324e-13, 1.183107e-13, 
    1.185529e-13, 1.190405e-13, 1.191495e-13, 1.192678e-13, 1.191946e-13, 
    1.188476e-13, 1.18791e-13, 1.185468e-13, 1.184798e-13, 1.182936e-13, 
    1.181397e-13, 1.182805e-13, 1.184284e-13, 1.188474e-13, 1.192297e-13, 
    1.196522e-13, 1.197553e-13, 1.202509e-13, 1.198485e-13, 1.205137e-13, 
    1.199498e-13, 1.209251e-13, 1.191702e-13, 1.199316e-13, 1.185637e-13, 
    1.187085e-13, 1.189713e-13, 1.195855e-13, 1.192518e-13, 1.196417e-13, 
    1.187887e-13, 1.183546e-13, 1.182414e-13, 1.180317e-13, 1.182462e-13, 
    1.182287e-13, 1.18434e-13, 1.18368e-13, 1.188613e-13, 1.185963e-13, 
    1.193564e-13, 1.196384e-13, 1.204338e-13, 1.20922e-13, 1.214177e-13, 
    1.216369e-13, 1.217036e-13, 1.217315e-13,
  1.688094e-17, 1.695295e-17, 1.693892e-17, 1.699712e-17, 1.696478e-17, 
    1.700295e-17, 1.689549e-17, 1.695585e-17, 1.691729e-17, 1.688736e-17, 
    1.711047e-17, 1.699971e-17, 1.722529e-17, 1.715458e-17, 1.733285e-17, 
    1.721434e-17, 1.735807e-17, 1.732912e-17, 1.741603e-17, 1.739112e-17, 
    1.750262e-17, 1.742753e-17, 1.756032e-17, 1.748462e-17, 1.74965e-17, 
    1.742507e-17, 1.702189e-17, 1.709671e-17, 1.701748e-17, 1.702814e-17, 
    1.702333e-17, 1.696549e-17, 1.693645e-17, 1.687537e-17, 1.688644e-17, 
    1.693126e-17, 1.703293e-17, 1.699831e-17, 1.70854e-17, 1.708343e-17, 
    1.718059e-17, 1.713677e-17, 1.730019e-17, 1.725368e-17, 1.739215e-17, 
    1.735627e-17, 1.739049e-17, 1.73801e-17, 1.739062e-17, 1.733799e-17, 
    1.736054e-17, 1.731469e-17, 1.714499e-17, 1.719485e-17, 1.704632e-17, 
    1.695736e-17, 1.689816e-17, 1.685625e-17, 1.686217e-17, 1.687349e-17, 
    1.693153e-17, 1.698606e-17, 1.702774e-17, 1.705565e-17, 1.708315e-17, 
    1.716672e-17, 1.721076e-17, 1.730965e-17, 1.729171e-17, 1.732228e-17, 
    1.73527e-17, 1.740429e-17, 1.739578e-17, 1.741854e-17, 1.732139e-17, 
    1.738589e-17, 1.728151e-17, 1.730904e-17, 1.709097e-17, 1.700763e-17, 
    1.697255e-17, 1.694163e-17, 1.686674e-17, 1.691847e-17, 1.689808e-17, 
    1.694652e-17, 1.697738e-17, 1.69621e-17, 1.705641e-17, 1.701973e-17, 
    1.721338e-17, 1.712989e-17, 1.734912e-17, 1.729539e-17, 1.736238e-17, 
    1.732739e-17, 1.738742e-17, 1.733335e-17, 1.742698e-17, 1.744743e-17, 
    1.743347e-17, 1.748701e-17, 1.733036e-17, 1.739052e-17, 1.696169e-17, 
    1.696418e-17, 1.697576e-17, 1.692489e-17, 1.692177e-17, 1.687509e-17, 
    1.691659e-17, 1.69343e-17, 1.697914e-17, 1.700577e-17, 1.703108e-17, 
    1.708677e-17, 1.714907e-17, 1.723618e-17, 1.729877e-17, 1.734194e-17, 
    1.731504e-17, 1.733873e-17, 1.731232e-17, 1.730039e-17, 1.74398e-17, 
    1.736077e-17, 1.747931e-17, 1.747273e-17, 1.74191e-17, 1.747347e-17, 
    1.696593e-17, 1.695159e-17, 1.690196e-17, 1.69408e-17, 1.687e-17, 
    1.690966e-17, 1.69325e-17, 1.702057e-17, 1.703987e-17, 1.705788e-17, 
    1.709338e-17, 1.713901e-17, 1.721915e-17, 1.72889e-17, 1.735446e-17, 
    1.73495e-17, 1.735125e-17, 1.73664e-17, 1.732894e-17, 1.737254e-17, 
    1.73799e-17, 1.736072e-17, 1.747185e-17, 1.744008e-17, 1.747259e-17, 
    1.745189e-17, 1.695624e-17, 1.698035e-17, 1.696733e-17, 1.699185e-17, 
    1.697459e-17, 1.705149e-17, 1.707457e-17, 1.718256e-17, 1.713813e-17, 
    1.720875e-17, 1.714528e-17, 1.715654e-17, 1.721121e-17, 1.714868e-17, 
    1.728512e-17, 1.719272e-17, 1.736698e-17, 1.727214e-17, 1.737313e-17, 
    1.735417e-17, 1.738553e-17, 1.741367e-17, 1.744901e-17, 1.751439e-17, 
    1.749923e-17, 1.755387e-17, 1.701632e-17, 1.70477e-17, 1.704487e-17, 
    1.707768e-17, 1.710196e-17, 1.715455e-17, 1.723905e-17, 1.720724e-17, 
    1.726558e-17, 1.727732e-17, 1.718866e-17, 1.724315e-17, 1.706866e-17, 
    1.709689e-17, 1.708003e-17, 1.701883e-17, 1.721466e-17, 1.711413e-17, 
    1.729982e-17, 1.724526e-17, 1.740966e-17, 1.732569e-17, 1.74909e-17, 
    1.756187e-17, 1.76284e-17, 1.770661e-17, 1.706476e-17, 1.704344e-17, 
    1.708156e-17, 1.713446e-17, 1.718339e-17, 1.72486e-17, 1.725524e-17, 
    1.726748e-17, 1.729912e-17, 1.732611e-17, 1.727142e-17, 1.73331e-17, 
    1.710357e-17, 1.722337e-17, 1.703544e-17, 1.709206e-17, 1.713131e-17, 
    1.711403e-17, 1.720359e-17, 1.722474e-17, 1.731078e-17, 1.726625e-17, 
    1.754441e-17, 1.741971e-17, 1.776597e-17, 1.766909e-17, 1.703601e-17, 
    1.706465e-17, 1.716455e-17, 1.711699e-17, 1.725292e-17, 1.728645e-17, 
    1.731367e-17, 1.73502e-17, 1.735415e-17, 1.73761e-17, 1.734014e-17, 
    1.737466e-17, 1.724874e-17, 1.730361e-17, 1.715305e-17, 1.71897e-17, 
    1.717281e-17, 1.715434e-17, 1.721137e-17, 1.727229e-17, 1.727348e-17, 
    1.729305e-17, 1.735001e-17, 1.725347e-17, 1.756072e-17, 1.736841e-17, 
    1.709591e-17, 1.71513e-17, 1.715909e-17, 1.713765e-17, 1.728309e-17, 
    1.723037e-17, 1.737555e-17, 1.733475e-17, 1.740159e-17, 1.736837e-17, 
    1.73635e-17, 1.732109e-17, 1.729591e-17, 1.72328e-17, 1.718147e-17, 
    1.714074e-17, 1.71502e-17, 1.719495e-17, 1.727599e-17, 1.735456e-17, 
    1.733674e-17, 1.739651e-17, 1.724306e-17, 1.730561e-17, 1.728146e-17, 
    1.734581e-17, 1.720642e-17, 1.732453e-17, 1.717638e-17, 1.718931e-17, 
    1.722932e-17, 1.730992e-17, 1.732799e-17, 1.734822e-17, 1.73357e-17, 
    1.727803e-17, 1.726867e-17, 1.722832e-17, 1.721724e-17, 1.718648e-17, 
    1.716108e-17, 1.718432e-17, 1.720875e-17, 1.727801e-17, 1.734169e-17, 
    1.741408e-17, 1.743177e-17, 1.751674e-17, 1.744771e-17, 1.756181e-17, 
    1.746502e-17, 1.763254e-17, 1.733147e-17, 1.746196e-17, 1.723111e-17, 
    1.725505e-17, 1.729848e-17, 1.740263e-17, 1.734549e-17, 1.741227e-17, 
    1.72683e-17, 1.719655e-17, 1.717786e-17, 1.714324e-17, 1.717866e-17, 
    1.717577e-17, 1.720969e-17, 1.719878e-17, 1.728031e-17, 1.72365e-17, 
    1.73634e-17, 1.741171e-17, 1.754818e-17, 1.763204e-17, 1.771733e-17, 
    1.775507e-17, 1.776655e-17, 1.777135e-17,
  7.070315e-22, 7.104262e-22, 7.097647e-22, 7.125093e-22, 7.109846e-22, 
    7.12784e-22, 7.077174e-22, 7.105626e-22, 7.087447e-22, 7.073345e-22, 
    7.178561e-22, 7.126314e-22, 7.232842e-22, 7.199418e-22, 7.283669e-22, 
    7.227659e-22, 7.2956e-22, 7.28192e-22, 7.323026e-22, 7.311237e-22, 
    7.364208e-22, 7.328469e-22, 7.392375e-22, 7.355493e-22, 7.361228e-22, 
    7.327304e-22, 7.136777e-22, 7.172059e-22, 7.134698e-22, 7.139722e-22, 
    7.137459e-22, 7.110175e-22, 7.096474e-22, 7.067697e-22, 7.07291e-22, 
    7.094033e-22, 7.14198e-22, 7.125658e-22, 7.166749e-22, 7.165819e-22, 
    7.211712e-22, 7.191005e-22, 7.268302e-22, 7.246287e-22, 7.311728e-22, 
    7.294754e-22, 7.310937e-22, 7.306023e-22, 7.311001e-22, 7.286112e-22, 
    7.296774e-22, 7.275162e-22, 7.194889e-22, 7.21845e-22, 7.1483e-22, 
    7.106331e-22, 7.078428e-22, 7.058688e-22, 7.061477e-22, 7.066804e-22, 
    7.094157e-22, 7.119885e-22, 7.13954e-22, 7.152707e-22, 7.165685e-22, 
    7.205138e-22, 7.22597e-22, 7.272778e-22, 7.264287e-22, 7.278709e-22, 
    7.293064e-22, 7.317467e-22, 7.313442e-22, 7.32421e-22, 7.278298e-22, 
    7.30876e-22, 7.25946e-22, 7.272494e-22, 7.169351e-22, 7.130054e-22, 
    7.113498e-22, 7.098923e-22, 7.063625e-22, 7.088e-22, 7.07839e-22, 
    7.101235e-22, 7.115787e-22, 7.108583e-22, 7.153067e-22, 7.135761e-22, 
    7.227207e-22, 7.187754e-22, 7.291374e-22, 7.266026e-22, 7.297646e-22, 
    7.281108e-22, 7.309485e-22, 7.283919e-22, 7.328208e-22, 7.337883e-22, 
    7.331274e-22, 7.35663e-22, 7.282506e-22, 7.310951e-22, 7.108387e-22, 
    7.109563e-22, 7.115026e-22, 7.09103e-22, 7.089556e-22, 7.067561e-22, 
    7.087118e-22, 7.095465e-22, 7.116621e-22, 7.129178e-22, 7.141115e-22, 
    7.167391e-22, 7.19681e-22, 7.237997e-22, 7.267628e-22, 7.28798e-22, 
    7.275325e-22, 7.286465e-22, 7.274047e-22, 7.268397e-22, 7.334267e-22, 
    7.296881e-22, 7.35298e-22, 7.349866e-22, 7.324471e-22, 7.350217e-22, 
    7.110386e-22, 7.103626e-22, 7.080221e-22, 7.098534e-22, 7.065166e-22, 
    7.083852e-22, 7.094616e-22, 7.136152e-22, 7.145262e-22, 7.153757e-22, 
    7.170515e-22, 7.192065e-22, 7.229943e-22, 7.26295e-22, 7.293902e-22, 
    7.291557e-22, 7.292383e-22, 7.299543e-22, 7.281834e-22, 7.30245e-22, 
    7.305926e-22, 7.29686e-22, 7.34945e-22, 7.334407e-22, 7.349801e-22, 
    7.340001e-22, 7.10582e-22, 7.117192e-22, 7.111048e-22, 7.122612e-22, 
    7.114474e-22, 7.150736e-22, 7.161625e-22, 7.212636e-22, 7.191647e-22, 
    7.225025e-22, 7.195024e-22, 7.200344e-22, 7.226172e-22, 7.196635e-22, 
    7.261155e-22, 7.217436e-22, 7.299821e-22, 7.255006e-22, 7.302728e-22, 
    7.293764e-22, 7.308595e-22, 7.321903e-22, 7.338635e-22, 7.369958e-22, 
    7.362565e-22, 7.389234e-22, 7.134154e-22, 7.14895e-22, 7.147623e-22, 
    7.163102e-22, 7.174566e-22, 7.199409e-22, 7.239362e-22, 7.224318e-22, 
    7.251918e-22, 7.257473e-22, 7.215531e-22, 7.241295e-22, 7.158841e-22, 
    7.172161e-22, 7.164211e-22, 7.135335e-22, 7.227819e-22, 7.180306e-22, 
    7.268123e-22, 7.242299e-22, 7.320009e-22, 7.280306e-22, 7.358503e-22, 
    7.393122e-22, 7.425642e-22, 7.463871e-22, 7.157004e-22, 7.146947e-22, 
    7.164937e-22, 7.189907e-22, 7.213037e-22, 7.243878e-22, 7.247023e-22, 
    7.252815e-22, 7.267797e-22, 7.280506e-22, 7.254672e-22, 7.283801e-22, 
    7.175303e-22, 7.231938e-22, 7.143169e-22, 7.169883e-22, 7.188423e-22, 
    7.180261e-22, 7.222593e-22, 7.232595e-22, 7.27331e-22, 7.252236e-22, 
    7.384594e-22, 7.324753e-22, 7.492945e-22, 7.445523e-22, 7.14344e-22, 
    7.156958e-22, 7.204128e-22, 7.181663e-22, 7.245925e-22, 7.261793e-22, 
    7.274684e-22, 7.291882e-22, 7.293753e-22, 7.304132e-22, 7.287132e-22, 
    7.30345e-22, 7.243944e-22, 7.269919e-22, 7.198699e-22, 7.216021e-22, 
    7.208041e-22, 7.199312e-22, 7.226271e-22, 7.255084e-22, 7.255658e-22, 
    7.264915e-22, 7.29176e-22, 7.246185e-22, 7.392538e-22, 7.300465e-22, 
    7.171713e-22, 7.197862e-22, 7.20155e-22, 7.191423e-22, 7.260203e-22, 
    7.235253e-22, 7.303873e-22, 7.284579e-22, 7.316192e-22, 7.300479e-22, 
    7.298171e-22, 7.27816e-22, 7.266273e-22, 7.236405e-22, 7.21213e-22, 
    7.192886e-22, 7.197355e-22, 7.218501e-22, 7.256838e-22, 7.293942e-22, 
    7.285515e-22, 7.313787e-22, 7.241259e-22, 7.270863e-22, 7.259428e-22, 
    7.289808e-22, 7.223928e-22, 7.279742e-22, 7.209725e-22, 7.215837e-22, 
    7.234758e-22, 7.272901e-22, 7.281391e-22, 7.290944e-22, 7.28503e-22, 
    7.257805e-22, 7.253378e-22, 7.234288e-22, 7.229042e-22, 7.214503e-22, 
    7.202495e-22, 7.213476e-22, 7.225024e-22, 7.2578e-22, 7.287859e-22, 
    7.3221e-22, 7.330473e-22, 7.371089e-22, 7.338003e-22, 7.39307e-22, 
    7.346176e-22, 7.427635e-22, 7.283013e-22, 7.344744e-22, 7.235606e-22, 
    7.246932e-22, 7.267481e-22, 7.316672e-22, 7.289658e-22, 7.321234e-22, 
    7.253201e-22, 7.219252e-22, 7.210428e-22, 7.194063e-22, 7.210803e-22, 
    7.209438e-22, 7.225474e-22, 7.220317e-22, 7.258888e-22, 7.238157e-22, 
    7.298124e-22, 7.320973e-22, 7.386452e-22, 7.42741e-22, 7.469134e-22, 
    7.487609e-22, 7.493232e-22, 7.495585e-22,
  9.118946e-27, 9.168647e-27, 9.15896e-27, 9.19917e-27, 9.176834e-27, 
    9.203197e-27, 9.128988e-27, 9.170642e-27, 9.144026e-27, 9.123385e-27, 
    9.277584e-27, 9.200962e-27, 9.357393e-27, 9.308254e-27, 9.432116e-27, 
    9.349764e-27, 9.449389e-27, 9.429596e-27, 9.489122e-27, 9.472042e-27, 
    9.548921e-27, 9.497009e-27, 9.590268e-27, 9.53618e-27, 9.544556e-27, 
    9.49532e-27, 9.216305e-27, 9.268039e-27, 9.213257e-27, 9.220618e-27, 
    9.217304e-27, 9.177311e-27, 9.15723e-27, 9.115123e-27, 9.12275e-27, 
    9.153663e-27, 9.223929e-27, 9.200007e-27, 9.260279e-27, 9.258914e-27, 
    9.326327e-27, 9.295895e-27, 9.409612e-27, 9.377195e-27, 9.472754e-27, 
    9.448174e-27, 9.471607e-27, 9.464491e-27, 9.4717e-27, 9.435662e-27, 
    9.451095e-27, 9.419713e-27, 9.301599e-27, 9.33623e-27, 9.233202e-27, 
    9.171664e-27, 9.130821e-27, 9.101943e-27, 9.106022e-27, 9.11381e-27, 
    9.153845e-27, 9.191547e-27, 9.22036e-27, 9.239672e-27, 9.258719e-27, 
    9.316641e-27, 9.347285e-27, 9.416199e-27, 9.403699e-27, 9.424896e-27, 
    9.445728e-27, 9.481064e-27, 9.475236e-27, 9.490833e-27, 9.424302e-27, 
    9.468449e-27, 9.396593e-27, 9.41579e-27, 9.26406e-27, 9.20645e-27, 
    9.182168e-27, 9.160828e-27, 9.109162e-27, 9.144831e-27, 9.130763e-27, 
    9.164219e-27, 9.185541e-27, 9.174985e-27, 9.2402e-27, 9.214818e-27, 
    9.349103e-27, 9.291114e-27, 9.443281e-27, 9.40626e-27, 9.452361e-27, 
    9.428415e-27, 9.469501e-27, 9.432492e-27, 9.496628e-27, 9.510647e-27, 
    9.501069e-27, 9.537835e-27, 9.430448e-27, 9.471623e-27, 9.174697e-27, 
    9.176419e-27, 9.184426e-27, 9.149267e-27, 9.14711e-27, 9.114922e-27, 
    9.143545e-27, 9.155764e-27, 9.186765e-27, 9.205165e-27, 9.222666e-27, 
    9.261218e-27, 9.304416e-27, 9.364985e-27, 9.40862e-27, 9.438369e-27, 
    9.419955e-27, 9.436178e-27, 9.41808e-27, 9.409757e-27, 9.505403e-27, 
    9.451249e-27, 9.532542e-27, 9.528027e-27, 9.49121e-27, 9.528536e-27, 
    9.177625e-27, 9.167723e-27, 9.133446e-27, 9.160264e-27, 9.111418e-27, 
    9.138759e-27, 9.154515e-27, 9.215382e-27, 9.228752e-27, 9.24121e-27, 
    9.265806e-27, 9.297452e-27, 9.353136e-27, 9.401726e-27, 9.446943e-27, 
    9.443548e-27, 9.444744e-27, 9.455106e-27, 9.429474e-27, 9.459317e-27, 
    9.464346e-27, 9.451223e-27, 9.527424e-27, 9.505614e-27, 9.527931e-27, 
    9.513723e-27, 9.170937e-27, 9.187599e-27, 9.178596e-27, 9.19554e-27, 
    9.183613e-27, 9.236769e-27, 9.252744e-27, 9.327674e-27, 9.296837e-27, 
    9.345899e-27, 9.301802e-27, 9.309615e-27, 9.34757e-27, 9.304171e-27, 
    9.399074e-27, 9.334728e-27, 9.455509e-27, 9.390009e-27, 9.45972e-27, 
    9.446743e-27, 9.468217e-27, 9.487492e-27, 9.511744e-27, 9.557368e-27, 
    9.546527e-27, 9.585663e-27, 9.212462e-27, 9.234155e-27, 9.232214e-27, 
    9.254925e-27, 9.27175e-27, 9.308246e-27, 9.366998e-27, 9.344868e-27, 
    9.385486e-27, 9.393663e-27, 9.331947e-27, 9.369839e-27, 9.248667e-27, 
    9.26821e-27, 9.256549e-27, 9.214189e-27, 9.350006e-27, 9.28017e-27, 
    9.409348e-27, 9.371323e-27, 9.484747e-27, 9.427231e-27, 9.540569e-27, 
    9.591353e-27, 9.64032e-27, 9.698113e-27, 9.245974e-27, 9.231223e-27, 
    9.257619e-27, 9.294273e-27, 9.328276e-27, 9.373646e-27, 9.378278e-27, 
    9.386805e-27, 9.408873e-27, 9.427534e-27, 9.38953e-27, 9.432323e-27, 
    9.272806e-27, 9.35607e-27, 9.225677e-27, 9.264863e-27, 9.292097e-27, 
    9.280113e-27, 9.342333e-27, 9.357046e-27, 9.416985e-27, 9.385954e-27, 
    9.578832e-27, 9.49161e-27, 9.742149e-27, 9.670359e-27, 9.22608e-27, 
    9.24591e-27, 9.315174e-27, 9.282173e-27, 9.376663e-27, 9.400024e-27, 
    9.419017e-27, 9.444012e-27, 9.446726e-27, 9.461749e-27, 9.437143e-27, 
    9.460765e-27, 9.373742e-27, 9.411997e-27, 9.307204e-27, 9.332662e-27, 
    9.320935e-27, 9.308104e-27, 9.347742e-27, 9.390135e-27, 9.390992e-27, 
    9.404619e-27, 9.443798e-27, 9.377046e-27, 9.59047e-27, 9.456405e-27, 
    9.267566e-27, 9.305958e-27, 9.311391e-27, 9.296512e-27, 9.397682e-27, 
    9.360954e-27, 9.461377e-27, 9.433448e-27, 9.479221e-27, 9.456463e-27, 
    9.453121e-27, 9.424101e-27, 9.406623e-27, 9.362645e-27, 9.326941e-27, 
    9.298662e-27, 9.30523e-27, 9.336307e-27, 9.39272e-27, 9.446995e-27, 
    9.434795e-27, 9.475736e-27, 9.369793e-27, 9.413382e-27, 9.396536e-27, 
    9.441014e-27, 9.344291e-27, 9.426377e-27, 9.323411e-27, 9.332396e-27, 
    9.360225e-27, 9.416375e-27, 9.428828e-27, 9.442655e-27, 9.434101e-27, 
    9.394145e-27, 9.38763e-27, 9.359537e-27, 9.351813e-27, 9.330436e-27, 
    9.312783e-27, 9.328923e-27, 9.345901e-27, 9.394142e-27, 9.438188e-27, 
    9.487774e-27, 9.499912e-27, 9.559007e-27, 9.510807e-27, 9.591249e-27, 
    9.522627e-27, 9.643291e-27, 9.43116e-27, 9.520574e-27, 9.361476e-27, 
    9.378146e-27, 9.408394e-27, 9.479899e-27, 9.440798e-27, 9.486512e-27, 
    9.387372e-27, 9.337405e-27, 9.324444e-27, 9.30039e-27, 9.324994e-27, 
    9.322989e-27, 9.34657e-27, 9.338986e-27, 9.395746e-27, 9.365229e-27, 
    9.45305e-27, 9.486137e-27, 9.581575e-27, 9.642976e-27, 9.706098e-27, 
    9.734071e-27, 9.74259e-27, 9.746156e-27,
  3.690674e-32, 3.714632e-32, 3.709961e-32, 3.729364e-32, 3.718585e-32, 
    3.731309e-32, 3.695514e-32, 3.715592e-32, 3.70276e-32, 3.692816e-32, 
    3.767701e-32, 3.73023e-32, 3.807498e-32, 3.782991e-32, 3.844818e-32, 
    3.803685e-32, 3.85333e-32, 3.843583e-32, 3.872932e-32, 3.864505e-32, 
    3.902418e-32, 3.876826e-32, 3.922683e-32, 3.896174e-32, 3.900285e-32, 
    3.875991e-32, 3.737644e-32, 3.76295e-32, 3.736171e-32, 3.739727e-32, 
    3.738127e-32, 3.718813e-32, 3.709121e-32, 3.688837e-32, 3.69251e-32, 
    3.707405e-32, 3.741326e-32, 3.729772e-32, 3.75911e-32, 3.758431e-32, 
    3.792001e-32, 3.776835e-32, 3.833605e-32, 3.817397e-32, 3.864856e-32, 
    3.852736e-32, 3.864289e-32, 3.860781e-32, 3.864335e-32, 3.84657e-32, 
    3.854175e-32, 3.838658e-32, 3.779675e-32, 3.796939e-32, 3.74581e-32, 
    3.71608e-32, 3.696396e-32, 3.682491e-32, 3.684454e-32, 3.688202e-32, 
    3.707492e-32, 3.725687e-32, 3.739605e-32, 3.748942e-32, 3.758333e-32, 
    3.78716e-32, 3.802451e-32, 3.836897e-32, 3.830648e-32, 3.841238e-32, 
    3.851531e-32, 3.868954e-32, 3.86608e-32, 3.873774e-32, 3.840947e-32, 
    3.862729e-32, 3.827095e-32, 3.836697e-32, 3.76097e-32, 3.732884e-32, 
    3.721151e-32, 3.710861e-32, 3.685965e-32, 3.703147e-32, 3.696367e-32, 
    3.712499e-32, 3.722787e-32, 3.717694e-32, 3.749197e-32, 3.736927e-32, 
    3.803359e-32, 3.774451e-32, 3.850324e-32, 3.831929e-32, 3.8548e-32, 
    3.842998e-32, 3.863249e-32, 3.845011e-32, 3.876636e-32, 3.883556e-32, 
    3.878827e-32, 3.896997e-32, 3.844004e-32, 3.864295e-32, 3.717554e-32, 
    3.718385e-32, 3.72225e-32, 3.705285e-32, 3.704246e-32, 3.688739e-32, 
    3.702529e-32, 3.708419e-32, 3.72338e-32, 3.732263e-32, 3.740719e-32, 
    3.759574e-32, 3.781076e-32, 3.811292e-32, 3.833109e-32, 3.847906e-32, 
    3.838781e-32, 3.846826e-32, 3.837844e-32, 3.83368e-32, 3.880966e-32, 
    3.854249e-32, 3.894379e-32, 3.892148e-32, 3.87396e-32, 3.892399e-32, 
    3.718967e-32, 3.71419e-32, 3.697662e-32, 3.710592e-32, 3.687053e-32, 
    3.700221e-32, 3.707814e-32, 3.737195e-32, 3.743661e-32, 3.749683e-32, 
    3.761858e-32, 3.777611e-32, 3.805376e-32, 3.829657e-32, 3.852131e-32, 
    3.850458e-32, 3.851047e-32, 3.856153e-32, 3.843524e-32, 3.858228e-32, 
    3.860706e-32, 3.854239e-32, 3.89185e-32, 3.881075e-32, 3.892101e-32, 
    3.885081e-32, 3.715741e-32, 3.723782e-32, 3.719436e-32, 3.727614e-32, 
    3.721856e-32, 3.747532e-32, 3.755354e-32, 3.792668e-32, 3.777303e-32, 
    3.801763e-32, 3.779778e-32, 3.783669e-32, 3.802588e-32, 3.780959e-32, 
    3.828327e-32, 3.796184e-32, 3.856351e-32, 3.82379e-32, 3.858427e-32, 
    3.852032e-32, 3.862619e-32, 3.872126e-32, 3.884101e-32, 3.906561e-32, 
    3.901254e-32, 3.920427e-32, 3.735788e-32, 3.74627e-32, 3.745335e-32, 
    3.756446e-32, 3.764814e-32, 3.782989e-32, 3.8123e-32, 3.801253e-32, 
    3.821541e-32, 3.825628e-32, 3.794807e-32, 3.813717e-32, 3.753332e-32, 
    3.763047e-32, 3.757252e-32, 3.736621e-32, 3.803812e-32, 3.768999e-32, 
    3.833472e-32, 3.814462e-32, 3.870771e-32, 3.842401e-32, 3.898337e-32, 
    3.923209e-32, 3.947455e-32, 3.976141e-32, 3.751995e-32, 3.744856e-32, 
    3.757787e-32, 3.776022e-32, 3.792973e-32, 3.815621e-32, 3.817938e-32, 
    3.822198e-32, 3.833237e-32, 3.842558e-32, 3.823557e-32, 3.844928e-32, 
    3.765325e-32, 3.80684e-32, 3.742173e-32, 3.761381e-32, 3.77494e-32, 
    3.768976e-32, 3.799989e-32, 3.807332e-32, 3.837292e-32, 3.821775e-32, 
    3.917069e-32, 3.874152e-32, 3.998392e-32, 3.962356e-32, 3.74237e-32, 
    3.751964e-32, 3.786438e-32, 3.770002e-32, 3.817131e-32, 3.828808e-32, 
    3.838313e-32, 3.850684e-32, 3.852023e-32, 3.859427e-32, 3.847302e-32, 
    3.858943e-32, 3.815669e-32, 3.834798e-32, 3.782472e-32, 3.795161e-32, 
    3.789316e-32, 3.78292e-32, 3.802688e-32, 3.823858e-32, 3.824293e-32, 
    3.831105e-32, 3.850557e-32, 3.817322e-32, 3.922762e-32, 3.856774e-32, 
    3.762734e-32, 3.781842e-32, 3.784555e-32, 3.777144e-32, 3.827637e-32, 
    3.809282e-32, 3.859244e-32, 3.845482e-32, 3.868046e-32, 3.856822e-32, 
    3.855174e-32, 3.840847e-32, 3.83211e-32, 3.810125e-32, 3.792307e-32, 
    3.778216e-32, 3.781487e-32, 3.796979e-32, 3.825152e-32, 3.852153e-32, 
    3.846141e-32, 3.866327e-32, 3.813698e-32, 3.835489e-32, 3.827061e-32, 
    3.849208e-32, 3.800964e-32, 3.841961e-32, 3.79055e-32, 3.795031e-32, 
    3.808918e-32, 3.836983e-32, 3.843204e-32, 3.850015e-32, 3.845804e-32, 
    3.825866e-32, 3.822611e-32, 3.808576e-32, 3.804717e-32, 3.794054e-32, 
    3.785252e-32, 3.793298e-32, 3.801765e-32, 3.825867e-32, 3.847814e-32, 
    3.872264e-32, 3.878259e-32, 3.907353e-32, 3.883628e-32, 3.923143e-32, 
    3.889452e-32, 3.948911e-32, 3.844343e-32, 3.88845e-32, 3.809545e-32, 
    3.817872e-32, 3.832991e-32, 3.868372e-32, 3.849102e-32, 3.871637e-32, 
    3.822482e-32, 3.797523e-32, 3.791065e-32, 3.779075e-32, 3.791339e-32, 
    3.79034e-32, 3.802104e-32, 3.798319e-32, 3.826669e-32, 3.811419e-32, 
    3.855137e-32, 3.871454e-32, 3.918421e-32, 3.948766e-32, 3.98012e-32, 
    3.994274e-32, 3.998621e-32, 4.00044e-32,
  4.88481e-38, 4.927285e-38, 4.918992e-38, 4.953486e-38, 4.934312e-38, 
    4.956951e-38, 4.893381e-38, 4.928987e-38, 4.90622e-38, 4.888606e-38, 
    5.02214e-38, 4.955029e-38, 5.094197e-38, 5.049783e-38, 5.163779e-38, 
    5.08727e-38, 5.179611e-38, 5.161495e-38, 5.216181e-38, 5.200446e-38, 
    5.271312e-38, 5.223461e-38, 5.308996e-38, 5.25971e-38, 5.267359e-38, 
    5.221899e-38, 4.968249e-38, 5.013575e-38, 4.965621e-38, 4.971959e-38, 
    4.96911e-38, 4.934715e-38, 4.917492e-38, 4.881566e-38, 4.888064e-38, 
    4.914452e-38, 4.974811e-38, 4.95422e-38, 5.006687e-38, 5.005464e-38, 
    5.066094e-38, 5.03866e-38, 5.142774e-38, 5.112413e-38, 5.201102e-38, 
    5.178515e-38, 5.200042e-38, 5.193501e-38, 5.200127e-38, 5.167045e-38, 
    5.181191e-38, 5.152262e-38, 5.043789e-38, 5.075041e-38, 4.98282e-38, 
    4.929845e-38, 4.894941e-38, 4.870346e-38, 4.873816e-38, 4.88044e-38, 
    4.914608e-38, 4.946947e-38, 4.97175e-38, 4.988419e-38, 5.005289e-38, 
    5.05731e-38, 5.085034e-38, 5.148949e-38, 5.137229e-38, 5.157093e-38, 
    5.176273e-38, 5.208747e-38, 5.203383e-38, 5.217751e-38, 5.156554e-38, 
    5.197127e-38, 5.130571e-38, 5.14858e-38, 5.010004e-38, 4.959763e-38, 
    4.93886e-38, 4.920588e-38, 4.876486e-38, 4.9069e-38, 4.894889e-38, 
    4.923503e-38, 4.941787e-38, 4.932731e-38, 4.988876e-38, 4.96697e-38, 
    5.086683e-38, 5.034346e-38, 5.174028e-38, 5.13963e-38, 5.182358e-38, 
    5.160403e-38, 5.198098e-38, 5.164151e-38, 5.223103e-38, 5.23605e-38, 
    5.2272e-38, 5.261262e-38, 5.162279e-38, 5.200049e-38, 4.932481e-38, 
    4.933957e-38, 4.940832e-38, 4.910692e-38, 4.908851e-38, 4.881391e-38, 
    4.90581e-38, 4.916253e-38, 4.942843e-38, 4.958657e-38, 4.973734e-38, 
    5.00752e-38, 5.046317e-38, 5.101097e-38, 5.141844e-38, 5.169533e-38, 
    5.152495e-38, 5.167525e-38, 5.150737e-38, 5.14292e-38, 5.2312e-38, 
    5.181328e-38, 5.256347e-38, 5.252161e-38, 5.218096e-38, 5.252633e-38, 
    4.934993e-38, 4.926506e-38, 4.897183e-38, 4.920115e-38, 4.87841e-38, 
    4.901717e-38, 4.915177e-38, 4.967442e-38, 4.978988e-38, 4.989742e-38, 
    5.011637e-38, 5.04006e-38, 5.09035e-38, 5.135367e-38, 5.177391e-38, 
    5.174278e-38, 5.175375e-38, 5.184876e-38, 5.161387e-38, 5.188743e-38, 
    5.193357e-38, 5.181313e-38, 5.251601e-38, 5.23141e-38, 5.252072e-38, 
    5.238912e-38, 4.929261e-38, 4.943556e-38, 4.935827e-38, 4.950374e-38, 
    4.940126e-38, 4.98589e-38, 4.999911e-38, 5.067293e-38, 5.039503e-38, 
    5.08379e-38, 5.043977e-38, 5.051011e-38, 5.085272e-38, 5.046114e-38, 
    5.132865e-38, 5.073661e-38, 5.185245e-38, 5.124356e-38, 5.189113e-38, 
    5.177207e-38, 5.196928e-38, 5.214671e-38, 5.237076e-38, 5.279011e-38, 
    5.269164e-38, 5.304801e-38, 4.964941e-38, 4.98364e-38, 4.981978e-38, 
    5.001889e-38, 5.016962e-38, 5.049785e-38, 5.102934e-38, 5.082872e-38, 
    5.120167e-38, 5.127819e-38, 5.071183e-38, 5.105526e-38, 4.99628e-38, 
    5.013768e-38, 5.003338e-38, 4.966421e-38, 5.087506e-38, 5.024502e-38, 
    5.142525e-38, 5.106922e-38, 5.212139e-38, 5.159272e-38, 5.263756e-38, 
    5.309967e-38, 5.35482e-38, 5.408624e-38, 4.993877e-38, 4.981123e-38, 
    5.004305e-38, 5.037181e-38, 5.067856e-38, 5.109088e-38, 5.113425e-38, 
    5.121396e-38, 5.142089e-38, 5.159577e-38, 5.123932e-38, 5.163997e-38, 
    5.01786e-38, 5.093009e-38, 4.976327e-38, 5.010764e-38, 5.035231e-38, 
    5.024468e-38, 5.080581e-38, 5.09391e-38, 5.149693e-38, 5.120606e-38, 
    5.298531e-38, 5.218447e-38, 5.451356e-38, 5.382426e-38, 4.976683e-38, 
    4.993825e-38, 5.056018e-38, 5.026321e-38, 5.111915e-38, 5.133779e-38, 
    5.151618e-38, 5.174693e-38, 5.17719e-38, 5.190975e-38, 5.16841e-38, 
    5.190075e-38, 5.109178e-38, 5.145017e-38, 5.048851e-38, 5.071822e-38, 
    5.061236e-38, 5.049661e-38, 5.085478e-38, 5.124494e-38, 5.125321e-38, 
    5.138082e-38, 5.17442e-38, 5.112273e-38, 5.30911e-38, 5.185997e-38, 
    5.013217e-38, 5.047697e-38, 5.052616e-38, 5.03922e-38, 5.131582e-38, 
    5.09745e-38, 5.190635e-38, 5.165026e-38, 5.207054e-38, 5.186124e-38, 
    5.183054e-38, 5.156367e-38, 5.139971e-38, 5.09898e-38, 5.066649e-38, 
    5.041158e-38, 5.047071e-38, 5.075115e-38, 5.126919e-38, 5.177427e-38, 
    5.166243e-38, 5.203846e-38, 5.105498e-38, 5.146308e-38, 5.130498e-38, 
    5.171951e-38, 5.082345e-38, 5.158419e-38, 5.063471e-38, 5.071589e-38, 
    5.096789e-38, 5.149104e-38, 5.160788e-38, 5.173448e-38, 5.165624e-38, 
    5.128259e-38, 5.122166e-38, 5.096169e-38, 5.089156e-38, 5.069819e-38, 
    5.05388e-38, 5.068446e-38, 5.083796e-38, 5.128266e-38, 5.169355e-38, 
    5.214928e-38, 5.22614e-38, 5.280464e-38, 5.236169e-38, 5.309817e-38, 
    5.247057e-38, 5.357482e-38, 5.162889e-38, 5.245201e-38, 5.097931e-38, 
    5.113303e-38, 5.141613e-38, 5.207647e-38, 5.171754e-38, 5.213748e-38, 
    5.121925e-38, 5.076096e-38, 5.064403e-38, 5.042708e-38, 5.064899e-38, 
    5.06309e-38, 5.084418e-38, 5.077552e-38, 5.129769e-38, 5.101337e-38, 
    5.182983e-38, 5.213409e-38, 5.301062e-38, 5.357233e-38, 5.416249e-38, 
    5.44343e-38, 5.451802e-38, 5.455309e-38,
  2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 
    2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.522337e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  6.828931e-06, 7.09688e-06, 7.044445e-06, 7.263109e-06, 7.141474e-06, 
    7.285154e-06, 6.882906e-06, 7.107592e-06, 6.963802e-06, 6.852895e-06, 
    7.695298e-06, 7.272935e-06, 8.139269e-06, 7.86367e-06, 8.562467e-06, 
    8.096115e-06, 8.657519e-06, 8.548946e-06, 8.877004e-06, 8.782683e-06, 
    9.205468e-06, 8.920621e-06, 9.426185e-06, 9.137308e-06, 9.182381e-06, 
    8.911248e-06, 7.3572e-06, 7.64218e-06, 7.340442e-06, 7.380776e-06, 
    7.362678e-06, 7.143961e-06, 7.034781e-06, 6.808674e-06, 6.849487e-06, 
    7.015694e-06, 7.398944e-06, 7.26791e-06, 7.600076e-06, 7.59251e-06, 
    7.964835e-06, 7.794836e-06, 8.435532e-06, 8.251588e-06, 8.786616e-06, 
    8.651105e-06, 8.780228e-06, 8.741026e-06, 8.780739e-06, 8.582241e-06, 
    8.667129e-06, 8.493069e-06, 7.826554e-06, 8.020339e-06, 7.450112e-06, 
    7.112852e-06, 6.892685e-06, 6.73829e-06, 6.760021e-06, 6.801526e-06, 
    7.01667e-06, 7.221674e-06, 7.379572e-06, 7.485974e-06, 7.591422e-06, 
    7.910005e-06, 8.082303e-06, 8.472864e-06, 8.401962e-06, 8.522219e-06, 
    8.637658e-06, 8.832397e-06, 8.800271e-06, 8.886335e-06, 8.51907e-06, 
    8.762669e-06, 8.361651e-06, 8.470756e-06, 7.620021e-06, 7.303172e-06, 
    7.170046e-06, 7.054505e-06, 6.776748e-06, 6.968023e-06, 6.892332e-06, 
    7.073038e-06, 7.188899e-06, 7.131501e-06, 7.488893e-06, 7.349076e-06, 
    8.092559e-06, 7.768052e-06, 8.624171e-06, 8.416502e-06, 8.674177e-06, 
    8.542404e-06, 8.768523e-06, 8.564942e-06, 8.918434e-06, 8.995864e-06, 
    8.94293e-06, 9.146693e-06, 8.553692e-06, 8.780211e-06, 7.129888e-06, 
    7.139234e-06, 7.182863e-06, 6.991939e-06, 6.980342e-06, 6.807549e-06, 
    6.961221e-06, 7.027109e-06, 7.195653e-06, 7.29612e-06, 7.392177e-06, 
    7.60518e-06, 7.842126e-06, 8.182285e-06, 8.429914e-06, 8.597241e-06, 
    8.494529e-06, 8.585189e-06, 8.483854e-06, 8.436496e-06, 8.966822e-06, 
    8.66791e-06, 9.117327e-06, 9.09233e-06, 8.888377e-06, 9.095147e-06, 
    7.145802e-06, 7.092067e-06, 6.906829e-06, 7.051612e-06, 6.788851e-06, 
    6.935364e-06, 7.020226e-06, 7.351951e-06, 7.425738e-06, 7.494374e-06, 
    7.630715e-06, 7.803501e-06, 8.115467e-06, 8.390591e-06, 8.644395e-06, 
    8.625725e-06, 8.632295e-06, 8.689261e-06, 8.54833e-06, 8.712462e-06, 
    8.740077e-06, 8.667897e-06, 9.088983e-06, 8.9682e-06, 9.091799e-06, 
    9.013116e-06, 7.109519e-06, 7.200139e-06, 7.151108e-06, 7.243418e-06, 
    7.178319e-06, 7.469624e-06, 7.557887e-06, 7.972122e-06, 7.800018e-06, 
    8.074658e-06, 7.827758e-06, 7.871277e-06, 8.083604e-06, 7.841034e-06, 
    8.375306e-06, 8.011585e-06, 8.691477e-06, 8.323595e-06, 8.714684e-06, 
    8.643293e-06, 8.761598e-06, 8.867898e-06, 9.002106e-06, 9.250795e-06, 
    9.193102e-06, 9.401781e-06, 7.336156e-06, 7.45533e-06, 7.444837e-06, 
    7.570338e-06, 7.663682e-06, 7.863761e-06, 8.193791e-06, 8.069095e-06, 
    8.298578e-06, 8.344908e-06, 7.996512e-06, 8.209759e-06, 7.535547e-06, 
    7.643722e-06, 7.579265e-06, 7.345509e-06, 8.097723e-06, 7.710307e-06, 
    8.434021e-06, 8.218295e-06, 8.852718e-06, 8.535373e-06, 9.161362e-06, 
    9.431678e-06, 9.6871e-06, 9.985784e-06, 7.520735e-06, 7.439379e-06, 
    7.585328e-06, 7.785528e-06, 7.975787e-06, 8.231393e-06, 8.257727e-06, 
    8.305979e-06, 8.431448e-06, 8.537393e-06, 8.321224e-06, 8.564019e-06, 
    7.668831e-06, 8.131994e-06, 7.408686e-06, 7.62508e-06, 7.773523e-06, 
    7.710236e-06, 8.054897e-06, 8.137734e-06, 8.477406e-06, 8.301242e-06, 
    9.364824e-06, 8.890345e-06, 1.021309e-05, 9.842374e-06, 7.411031e-06, 
    7.520468e-06, 7.902274e-06, 7.721746e-06, 8.248578e-06, 8.381015e-06, 
    8.489219e-06, 8.628111e-06, 8.64317e-06, 8.725819e-06, 8.590499e-06, 
    8.720475e-06, 8.231939e-06, 8.449159e-06, 7.858005e-06, 8.000407e-06, 
    7.934785e-06, 7.863021e-06, 8.085312e-06, 8.324606e-06, 8.329797e-06, 
    8.407044e-06, 8.625844e-06, 8.250752e-06, 9.426265e-06, 8.695398e-06, 
    7.64053e-06, 7.850601e-06, 7.881277e-06, 7.798351e-06, 8.367703e-06, 
    8.159692e-06, 8.72381e-06, 8.570196e-06, 8.822296e-06, 8.696764e-06, 
    8.678335e-06, 8.517961e-06, 8.418563e-06, 8.169179e-06, 7.968275e-06, 
    7.810363e-06, 7.846973e-06, 8.020822e-06, 8.339333e-06, 8.644511e-06, 
    8.577364e-06, 8.803068e-06, 8.209697e-06, 8.456905e-06, 8.361048e-06, 
    8.611716e-06, 8.065779e-06, 8.52978e-06, 7.94866e-06, 7.999027e-06, 
    8.155582e-06, 8.473724e-06, 8.544726e-06, 8.620641e-06, 8.573785e-06, 
    8.347486e-06, 8.310623e-06, 8.151776e-06, 8.108087e-06, 7.988055e-06, 
    7.889175e-06, 7.979485e-06, 8.074742e-06, 8.347603e-06, 8.596068e-06, 
    8.869406e-06, 8.936654e-06, 9.258983e-06, 8.996341e-06, 9.430353e-06, 
    9.061007e-06, 9.7016e-06, 8.557005e-06, 9.050297e-06, 8.16275e-06, 
    8.256999e-06, 8.428357e-06, 8.825592e-06, 8.610533e-06, 8.862208e-06, 
    8.309185e-06, 8.026821e-06, 7.954419e-06, 7.819917e-06, 7.957505e-06, 
    7.946281e-06, 8.078734e-06, 8.036082e-06, 8.356717e-06, 8.183931e-06, 
    8.677857e-06, 8.860226e-06, 9.379859e-06, 9.700511e-06, 1.002748e-05, 
    1.017166e-05, 1.021551e-05, 1.023383e-05,
  7.384479e-06, 7.256267e-06, 7.28086e-06, 7.179917e-06, 7.235556e-06, 
    7.169977e-06, 7.35815e-06, 7.251264e-06, 7.319156e-06, 7.372768e-06, 
    6.992725e-06, 7.175483e-06, 6.518623e-06, 6.590724e-06, 6.418115e-06, 
    6.529555e-06, 6.39721e-06, 6.42115e-06, 6.351246e-06, 6.37061e-06, 
    6.288383e-06, 6.34249e-06, 6.250149e-06, 6.300848e-06, 6.292573e-06, 
    6.34436e-06, 7.137797e-06, 7.014844e-06, 7.145243e-06, 7.127351e-06, 
    7.135367e-06, 7.234397e-06, 7.285394e-06, 7.39445e-06, 7.374432e-06, 
    7.294438e-06, 7.119339e-06, 7.177767e-06, 7.032629e-06, 7.035828e-06, 
    6.563645e-06, 6.609568e-06, 6.446995e-06, 6.490772e-06, 6.369791e-06, 
    6.398612e-06, 6.37112e-06, 6.37935e-06, 6.371014e-06, 6.413726e-06, 
    6.395137e-06, 6.433776e-06, 6.600842e-06, 6.549089e-06, 7.096947e-06, 
    7.248791e-06, 7.353399e-06, 7.429317e-06, 7.418502e-06, 7.39796e-06, 
    7.293975e-06, 7.198737e-06, 7.127901e-06, 7.081395e-06, 7.036288e-06, 
    6.578208e-06, 6.53309e-06, 6.438386e-06, 6.454815e-06, 6.427158e-06, 
    6.401539e-06, 6.360327e-06, 6.366954e-06, 6.349358e-06, 6.427876e-06, 
    6.374789e-06, 6.464305e-06, 6.438877e-06, 7.024141e-06, 7.161899e-06, 
    7.222336e-06, 7.27612e-06, 7.410205e-06, 7.317127e-06, 7.353567e-06, 
    7.267431e-06, 7.213715e-06, 7.240182e-06, 7.080134e-06, 7.141408e-06, 
    6.530469e-06, 6.616982e-06, 6.404486e-06, 6.451419e-06, 6.393619e-06, 
    6.422621e-06, 6.373564e-06, 6.417578e-06, 6.342924e-06, 6.327675e-06, 
    6.338056e-06, 6.299121e-06, 6.42009e-06, 6.37112e-06, 7.240926e-06, 
    7.236595e-06, 7.216488e-06, 7.305718e-06, 7.311247e-06, 7.395e-06, 
    7.320392e-06, 7.28904e-06, 7.210627e-06, 7.165062e-06, 7.122333e-06, 
    7.030465e-06, 6.596579e-06, 6.507854e-06, 6.448299e-06, 6.410411e-06, 
    6.433447e-06, 6.413077e-06, 6.435881e-06, 6.446777e-06, 6.333346e-06, 
    6.394966e-06, 6.304564e-06, 6.309243e-06, 6.348945e-06, 6.308713e-06, 
    7.233557e-06, 7.25853e-06, 7.346555e-06, 7.277495e-06, 7.404224e-06, 
    7.332791e-06, 7.292285e-06, 7.140113e-06, 7.107601e-06, 7.07776e-06, 
    7.019723e-06, 6.607177e-06, 6.524648e-06, 6.457475e-06, 6.400073e-06, 
    6.404149e-06, 6.402711e-06, 6.390372e-06, 6.42129e-06, 6.38541e-06, 
    6.379546e-06, 6.394974e-06, 6.309872e-06, 6.333082e-06, 6.309342e-06, 
    6.324339e-06, 7.250394e-06, 7.208569e-06, 7.231108e-06, 7.188846e-06, 
    7.218565e-06, 7.088452e-06, 7.050497e-06, 6.561711e-06, 6.608135e-06, 
    6.535055e-06, 6.600515e-06, 6.588662e-06, 6.532744e-06, 6.596889e-06, 
    6.461063e-06, 6.551357e-06, 6.389896e-06, 6.473338e-06, 6.384937e-06, 
    6.400313e-06, 6.375021e-06, 6.353086e-06, 6.326469e-06, 6.280277e-06, 
    6.290632e-06, 6.254224e-06, 7.147158e-06, 7.094673e-06, 7.099259e-06, 
    7.045226e-06, 7.005926e-06, 6.590705e-06, 6.504999e-06, 6.536492e-06, 
    6.479371e-06, 6.468275e-06, 6.555319e-06, 6.50104e-06, 7.060055e-06, 
    7.014244e-06, 7.041429e-06, 7.142984e-06, 6.529155e-06, 6.986564e-06, 
    6.447345e-06, 6.498939e-06, 6.356172e-06, 6.42419e-06, 6.29642e-06, 
    6.24923e-06, 6.209082e-06, 6.167578e-06, 7.066413e-06, 7.10164e-06, 
    7.038869e-06, 6.612129e-06, 6.560757e-06, 6.495714e-06, 6.489274e-06, 
    6.477586e-06, 6.447947e-06, 6.423747e-06, 6.473919e-06, 6.417784e-06, 
    7.003725e-06, 6.520465e-06, 7.115067e-06, 7.022059e-06, 6.615462e-06, 
    6.986612e-06, 6.540148e-06, 6.519027e-06, 6.437348e-06, 6.47873e-06, 
    6.260449e-06, 6.348541e-06, 6.140008e-06, 6.186763e-06, 7.114048e-06, 
    7.066534e-06, 6.580302e-06, 6.981868e-06, 6.491508e-06, 6.459729e-06, 
    6.434657e-06, 6.40362e-06, 6.400338e-06, 6.382567e-06, 6.411901e-06, 
    6.383705e-06, 6.49558e-06, 6.443846e-06, 6.59227e-06, 6.554294e-06, 
    6.57162e-06, 6.590908e-06, 6.532337e-06, 6.473108e-06, 6.471879e-06, 
    6.453621e-06, 6.404078e-06, 6.490976e-06, 6.250109e-06, 6.38902e-06, 
    7.01561e-06, 6.594264e-06, 6.585962e-06, 6.608601e-06, 6.462869e-06, 
    6.513505e-06, 6.382996e-06, 6.416407e-06, 6.362405e-06, 6.388764e-06, 
    6.392722e-06, 6.428128e-06, 6.450939e-06, 6.511128e-06, 6.562736e-06, 
    6.605293e-06, 6.595271e-06, 6.548966e-06, 6.469593e-06, 6.400041e-06, 
    6.414805e-06, 6.366375e-06, 6.501063e-06, 6.442055e-06, 6.464438e-06, 
    6.407219e-06, 6.537341e-06, 6.425422e-06, 6.567933e-06, 6.554661e-06, 
    6.514535e-06, 6.438183e-06, 6.422099e-06, 6.405256e-06, 6.415609e-06, 
    6.467656e-06, 6.476468e-06, 6.515493e-06, 6.526525e-06, 6.557538e-06, 
    6.583837e-06, 6.559786e-06, 6.535035e-06, 6.467633e-06, 6.410663e-06, 
    6.352779e-06, 6.339303e-06, 6.27881e-06, 6.32757e-06, 6.249429e-06, 
    6.315119e-06, 6.206908e-06, 6.419327e-06, 6.317179e-06, 6.512743e-06, 
    6.489453e-06, 6.448651e-06, 6.361712e-06, 6.407479e-06, 6.354232e-06, 
    6.476815e-06, 6.547399e-06, 6.566406e-06, 6.602666e-06, 6.565589e-06, 
    6.568564e-06, 6.534021e-06, 6.545012e-06, 6.46547e-06, 6.507455e-06, 
    6.392821e-06, 6.354638e-06, 6.257912e-06, 6.207083e-06, 6.162269e-06, 
    6.144776e-06, 6.139736e-06, 6.137668e-06,
  9.865213e-06, 9.872855e-06, 9.871599e-06, 9.876066e-06, 9.873833e-06, 
    9.876403e-06, 9.866996e-06, 9.873097e-06, 9.86944e-06, 9.86602e-06, 
    9.878866e-06, 9.876218e-06, 1.019468e-05, 1.024287e-05, 1.01198e-05, 
    1.020225e-05, 1.01028e-05, 1.012222e-05, 1.006329e-05, 1.008033e-05, 
    1.000328e-05, 1.005538e-05, 9.962342e-06, 1.001583e-05, 1.000754e-05, 
    1.005708e-05, 9.877361e-06, 9.878955e-06, 9.877158e-06, 9.877625e-06, 
    9.877424e-06, 9.873884e-06, 9.871354e-06, 9.864511e-06, 9.865907e-06, 
    9.870861e-06, 9.877813e-06, 9.876142e-06, 9.878948e-06, 9.878937e-06, 
    1.022524e-05, 1.025485e-05, 1.01424e-05, 1.017494e-05, 1.007962e-05, 
    1.010397e-05, 1.008077e-05, 1.008783e-05, 1.008068e-05, 1.011628e-05, 
    1.010109e-05, 1.013218e-05, 1.024933e-05, 1.021554e-05, 9.878267e-06, 
    9.873213e-06, 9.867306e-06, 9.861941e-06, 9.862757e-06, 9.86426e-06, 
    9.870886e-06, 9.875376e-06, 9.877614e-06, 9.878519e-06, 9.878935e-06, 
    1.023478e-05, 1.020468e-05, 1.013576e-05, 1.014836e-05, 1.012698e-05, 
    1.010638e-05, 1.007135e-05, 1.007715e-05, 1.006159e-05, 1.012755e-05, 
    1.008392e-05, 1.015551e-05, 1.013615e-05, 9.878956e-06, 9.876664e-06, 
    9.874412e-06, 9.871849e-06, 9.863372e-06, 9.869559e-06, 9.867295e-06, 
    9.872299e-06, 9.874779e-06, 9.873622e-06, 9.878537e-06, 9.877264e-06, 
    1.020288e-05, 1.025949e-05, 1.010879e-05, 1.014578e-05, 1.009983e-05, 
    1.01234e-05, 1.008287e-05, 1.011937e-05, 1.005578e-05, 1.004169e-05, 
    1.005133e-05, 1.001412e-05, 1.012138e-05, 1.008077e-05, 9.873587e-06, 
    9.873786e-06, 9.874664e-06, 9.870224e-06, 9.869905e-06, 9.864472e-06, 
    9.869366e-06, 9.871158e-06, 9.874906e-06, 9.876564e-06, 9.877745e-06, 
    9.878953e-06, 1.024662e-05, 1.018713e-05, 1.01434e-05, 1.011361e-05, 
    1.013192e-05, 1.011576e-05, 1.013382e-05, 1.014224e-05, 1.004698e-05, 
    1.010095e-05, 1.00195e-05, 1.002408e-05, 1.006122e-05, 1.002357e-05, 
    9.873923e-06, 9.872746e-06, 9.867747e-06, 9.871778e-06, 9.863809e-06, 
    9.868612e-06, 9.870979e-06, 9.877298e-06, 9.878066e-06, 9.878569e-06, 
    9.878967e-06, 1.025334e-05, 1.019887e-05, 1.015037e-05, 1.010517e-05, 
    1.010851e-05, 1.010734e-05, 1.009713e-05, 1.012234e-05, 1.009296e-05, 
    1.008799e-05, 1.010096e-05, 1.00247e-05, 1.004674e-05, 1.002418e-05, 
    1.003856e-05, 9.873142e-06, 9.874989e-06, 9.874033e-06, 9.875747e-06, 
    9.874576e-06, 9.878408e-06, 9.878851e-06, 1.022395e-05, 1.025395e-05, 
    1.020602e-05, 1.024913e-05, 1.024155e-05, 1.020443e-05, 1.024682e-05, 
    1.015307e-05, 1.021705e-05, 1.009673e-05, 1.01622e-05, 1.009256e-05, 
    1.010537e-05, 1.008413e-05, 1.006493e-05, 1.004057e-05, 9.994927e-06, 
    1.000557e-05, 9.966906e-06, 9.877104e-06, 9.878307e-06, 9.878227e-06, 
    9.87889e-06, 9.878941e-06, 1.024286e-05, 1.018512e-05, 1.020701e-05, 
    1.016665e-05, 1.015846e-05, 1.021971e-05, 1.01823e-05, 9.878772e-06, 
    9.87896e-06, 9.878911e-06, 9.877221e-06, 1.020198e-05, 9.878824e-06, 
    1.014267e-05, 1.018081e-05, 1.006768e-05, 1.012463e-05, 1.001141e-05, 
    9.961301e-06, 9.913195e-06, 9.855741e-06, 9.878708e-06, 9.878182e-06, 
    9.878924e-06, 1.025645e-05, 1.022333e-05, 1.01785e-05, 1.017386e-05, 
    1.016534e-05, 1.014313e-05, 1.012429e-05, 1.016264e-05, 1.011954e-05, 
    9.878927e-06, 1.019597e-05, 9.877908e-06, 9.878962e-06, 1.025854e-05, 
    9.878827e-06, 1.02095e-05, 1.019497e-05, 1.013496e-05, 1.016618e-05, 
    9.973762e-06, 1.006085e-05, 9.811118e-06, 9.883485e-06, 9.877932e-06, 
    9.878708e-06, 1.023615e-05, 9.878784e-06, 1.017547e-05, 1.015207e-05, 
    1.013287e-05, 1.010808e-05, 1.010539e-05, 1.009056e-05, 1.011481e-05, 
    1.009152e-05, 1.01784e-05, 1.013999e-05, 1.024387e-05, 1.021903e-05, 
    1.023049e-05, 1.0243e-05, 1.020417e-05, 1.016204e-05, 1.016114e-05, 
    1.014745e-05, 1.010843e-05, 1.017509e-05, 9.962274e-06, 1.009597e-05, 
    9.878965e-06, 1.024514e-05, 1.023981e-05, 1.025424e-05, 1.015443e-05, 
    1.019111e-05, 1.009092e-05, 1.011844e-05, 1.007318e-05, 1.009578e-05, 
    1.009909e-05, 1.012775e-05, 1.014542e-05, 1.018944e-05, 1.022464e-05, 
    1.025216e-05, 1.024579e-05, 1.021545e-05, 1.015944e-05, 1.010514e-05, 
    1.011715e-05, 1.007665e-05, 1.018232e-05, 1.01386e-05, 1.01556e-05, 
    1.011102e-05, 1.020759e-05, 1.012559e-05, 1.022807e-05, 1.021927e-05, 
    1.019183e-05, 1.01356e-05, 1.012298e-05, 1.010941e-05, 1.01178e-05, 
    1.0158e-05, 1.016452e-05, 1.019251e-05, 1.020017e-05, 1.022119e-05, 
    1.023844e-05, 1.022268e-05, 1.020601e-05, 1.015799e-05, 1.011381e-05, 
    1.006466e-05, 1.005247e-05, 9.993385e-06, 1.004159e-05, 9.961507e-06, 
    1.002974e-05, 9.910386e-06, 1.012076e-05, 1.003174e-05, 1.019058e-05, 
    1.017399e-05, 1.014366e-05, 1.007256e-05, 1.011123e-05, 1.006595e-05, 
    1.016478e-05, 1.02144e-05, 1.022706e-05, 1.025049e-05, 1.022652e-05, 
    1.022848e-05, 1.020532e-05, 1.021279e-05, 1.015637e-05, 1.018686e-05, 
    1.009917e-05, 1.006631e-05, 9.970985e-06, 9.910624e-06, 9.847644e-06, 
    9.819327e-06, 9.810647e-06, 9.807009e-06,
  4.318736e-06, 4.232435e-06, 4.249199e-06, 4.179705e-06, 4.218241e-06, 
    4.172759e-06, 4.301227e-06, 4.22901e-06, 4.275098e-06, 4.310964e-06, 
    4.04526e-06, 4.176609e-06, 3.909788e-06, 3.993093e-06, 3.784401e-06, 
    3.922728e-06, 3.756619e-06, 3.788389e-06, 3.692944e-06, 3.72024e-06, 
    3.598665e-06, 3.680359e-06, 3.535988e-06, 3.618145e-06, 3.605263e-06, 
    3.683059e-06, 4.150139e-06, 4.061578e-06, 4.155392e-06, 4.142746e-06, 
    4.148422e-06, 4.217442e-06, 4.25227e-06, 4.325345e-06, 4.31207e-06, 
    4.258407e-06, 4.137061e-06, 4.178209e-06, 4.074629e-06, 4.076964e-06, 
    3.962363e-06, 4.014122e-06, 3.821739e-06, 3.87626e-06, 3.719101e-06, 
    3.758511e-06, 3.720948e-06, 3.732332e-06, 3.7208e-06, 3.778632e-06, 
    3.753833e-06, 3.804799e-06, 4.004419e-06, 3.945576e-06, 4.121103e-06, 
    4.22731e-06, 4.298056e-06, 4.348329e-06, 4.341218e-06, 4.327664e-06, 
    4.258093e-06, 4.192809e-06, 4.14314e-06, 4.109958e-06, 4.0773e-06, 
    3.97895e-06, 3.926892e-06, 3.810727e-06, 3.831654e-06, 3.79622e-06, 
    3.762436e-06, 3.705833e-06, 3.715139e-06, 3.69024e-06, 3.79716e-06, 
    3.726033e-06, 3.843581e-06, 3.811364e-06, 4.068397e-06, 4.167105e-06, 
    4.209127e-06, 4.245975e-06, 4.335751e-06, 4.273729e-06, 4.298166e-06, 
    4.240062e-06, 4.203185e-06, 4.22142e-06, 4.109051e-06, 4.152689e-06, 
    3.923809e-06, 4.022314e-06, 3.766374e-06, 3.827357e-06, 3.751784e-06, 
    3.790315e-06, 3.724338e-06, 3.783707e-06, 3.680984e-06, 3.658685e-06, 
    3.67392e-06, 3.615479e-06, 3.787002e-06, 3.720946e-06, 4.221929e-06, 
    4.218955e-06, 4.205102e-06, 4.266034e-06, 4.269767e-06, 4.325708e-06, 
    4.27593e-06, 4.25475e-06, 4.201051e-06, 4.169322e-06, 4.139191e-06, 
    4.073046e-06, 3.999653e-06, 3.896923e-06, 3.823399e-06, 3.774252e-06, 
    3.804377e-06, 3.777778e-06, 3.807513e-06, 3.821466e-06, 3.667035e-06, 
    3.7536e-06, 3.623873e-06, 3.631028e-06, 3.689647e-06, 3.630222e-06, 
    4.216867e-06, 4.233987e-06, 4.293482e-06, 4.246914e-06, 4.331805e-06, 
    4.28426e-06, 4.256946e-06, 4.15177e-06, 4.128714e-06, 4.107341e-06, 
    4.065181e-06, 4.01147e-06, 3.916943e-06, 3.835003e-06, 3.760474e-06, 
    3.765926e-06, 3.764006e-06, 3.747387e-06, 3.788573e-06, 3.740634e-06, 
    3.732596e-06, 3.753614e-06, 3.631987e-06, 3.666654e-06, 3.631181e-06, 
    3.653745e-06, 4.228422e-06, 4.199625e-06, 4.215182e-06, 4.185932e-06, 
    4.206534e-06, 4.115017e-06, 4.08763e-06, 3.960136e-06, 4.012531e-06, 
    3.929203e-06, 4.004057e-06, 3.990775e-06, 3.926476e-06, 4.000008e-06, 
    3.839507e-06, 3.948194e-06, 3.746742e-06, 3.854808e-06, 3.739988e-06, 
    3.760795e-06, 3.72636e-06, 3.695567e-06, 3.656904e-06, 3.585775e-06, 
    3.602222e-06, 3.54291e-06, 4.156743e-06, 4.119476e-06, 4.122761e-06, 
    4.083809e-06, 4.055033e-06, 3.993076e-06, 3.893494e-06, 3.930895e-06, 
    3.862284e-06, 3.848533e-06, 3.95279e-06, 3.888717e-06, 4.094564e-06, 
    4.061149e-06, 4.081044e-06, 4.153798e-06, 3.922263e-06, 4.040705e-06, 
    3.822185e-06, 3.88618e-06, 3.699953e-06, 3.792354e-06, 3.611281e-06, 
    3.534411e-06, 3.462423e-06, 3.378697e-06, 4.099162e-06, 4.124462e-06, 
    4.079182e-06, 4.01695e-06, 3.959049e-06, 3.882271e-06, 3.874432e-06, 
    3.86008e-06, 3.822953e-06, 3.791784e-06, 3.855538e-06, 3.783978e-06, 
    4.053394e-06, 3.911984e-06, 4.134027e-06, 4.066886e-06, 4.020637e-06, 
    4.040746e-06, 3.935175e-06, 3.910281e-06, 3.809394e-06, 3.861493e-06, 
    3.553345e-06, 3.689061e-06, 3.315298e-06, 3.418828e-06, 4.133305e-06, 
    4.099251e-06, 3.981337e-06, 4.037222e-06, 3.877157e-06, 3.837842e-06, 
    3.805938e-06, 3.765216e-06, 3.760829e-06, 3.736745e-06, 3.776224e-06, 
    3.738305e-06, 3.882108e-06, 3.817726e-06, 3.994835e-06, 3.951604e-06, 
    3.971484e-06, 3.993305e-06, 3.926019e-06, 3.854532e-06, 3.853016e-06, 
    3.830141e-06, 3.765795e-06, 3.87651e-06, 3.535889e-06, 3.745522e-06, 
    4.062162e-06, 3.997058e-06, 3.987736e-06, 4.013053e-06, 3.84178e-06, 
    3.903695e-06, 3.737333e-06, 3.782168e-06, 3.708762e-06, 3.745204e-06, 
    3.750571e-06, 3.797488e-06, 3.826749e-06, 3.900851e-06, 3.961321e-06, 
    4.009381e-06, 3.998198e-06, 3.945433e-06, 3.850168e-06, 3.760427e-06, 
    3.780051e-06, 3.714331e-06, 3.888751e-06, 3.815433e-06, 3.843739e-06, 
    3.770014e-06, 3.931887e-06, 3.793939e-06, 3.967276e-06, 3.95203e-06, 
    3.904926e-06, 3.810463e-06, 3.789633e-06, 3.767398e-06, 3.781117e-06, 
    3.847757e-06, 3.858698e-06, 3.906072e-06, 3.919165e-06, 3.955349e-06, 
    3.985342e-06, 3.957934e-06, 3.929183e-06, 3.847732e-06, 3.774581e-06, 
    3.695127e-06, 3.675737e-06, 3.583403e-06, 3.658517e-06, 3.534727e-06, 
    3.639896e-06, 3.458278e-06, 3.785985e-06, 3.643018e-06, 3.902788e-06, 
    3.874651e-06, 3.823837e-06, 3.707774e-06, 3.77036e-06, 3.697191e-06, 
    3.859127e-06, 3.94361e-06, 3.965529e-06, 4.006454e-06, 3.964594e-06, 
    3.967996e-06, 3.927999e-06, 3.940846e-06, 3.845033e-06, 3.896451e-06, 
    3.750703e-06, 3.69777e-06, 3.549113e-06, 3.458626e-06, 3.367085e-06, 
    3.326855e-06, 3.314635e-06, 3.309529e-06,
  4.426445e-07, 4.259535e-07, 4.291688e-07, 4.159239e-07, 4.23241e-07, 
    4.146122e-07, 4.392305e-07, 4.252981e-07, 4.341618e-07, 4.411273e-07, 
    3.909277e-07, 4.15339e-07, 3.665235e-07, 3.81396e-07, 3.447263e-07, 
    3.688131e-07, 3.399918e-07, 3.454086e-07, 3.292705e-07, 3.338444e-07, 
    3.137266e-07, 3.271728e-07, 3.036103e-07, 3.169061e-07, 3.148017e-07, 
    3.276223e-07, 4.103561e-07, 3.939177e-07, 4.113424e-07, 4.089701e-07, 
    4.100339e-07, 4.230885e-07, 4.297592e-07, 4.439371e-07, 4.413431e-07, 
    4.309403e-07, 4.079061e-07, 4.156412e-07, 3.963176e-07, 3.967479e-07, 
    3.758733e-07, 3.852e-07, 3.511434e-07, 3.606259e-07, 3.336528e-07, 
    3.403131e-07, 3.339635e-07, 3.358812e-07, 3.339386e-07, 3.437402e-07, 
    3.395189e-07, 3.482242e-07, 3.834423e-07, 3.728744e-07, 4.049271e-07, 
    4.24973e-07, 4.386135e-07, 4.484475e-07, 4.470494e-07, 4.443909e-07, 
    4.308799e-07, 4.184044e-07, 4.090439e-07, 4.028534e-07, 3.968098e-07, 
    3.788491e-07, 3.695514e-07, 3.492443e-07, 3.528579e-07, 3.467508e-07, 
    3.409803e-07, 3.314261e-07, 3.329871e-07, 3.288191e-07, 3.46912e-07, 
    3.348194e-07, 3.549263e-07, 3.49354e-07, 3.951707e-07, 4.135461e-07, 
    4.215043e-07, 4.285494e-07, 4.45976e-07, 4.338971e-07, 4.386351e-07, 
    4.274146e-07, 4.203741e-07, 4.238477e-07, 4.026849e-07, 4.108347e-07, 
    3.690048e-07, 3.866872e-07, 3.416502e-07, 3.521144e-07, 3.391715e-07, 
    3.457384e-07, 3.345339e-07, 3.446075e-07, 3.272768e-07, 3.235767e-07, 
    3.261022e-07, 3.164699e-07, 3.451713e-07, 3.339631e-07, 4.23945e-07, 
    4.233772e-07, 4.207386e-07, 4.324109e-07, 4.331314e-07, 4.440081e-07, 
    4.343227e-07, 4.302364e-07, 4.199686e-07, 4.13964e-07, 4.083045e-07, 
    3.960261e-07, 3.825805e-07, 3.642545e-07, 3.514301e-07, 3.429926e-07, 
    3.481516e-07, 3.435944e-07, 3.48691e-07, 3.510962e-07, 3.249596e-07, 
    3.394794e-07, 3.178441e-07, 3.19018e-07, 3.287202e-07, 3.188856e-07, 
    4.229789e-07, 4.262505e-07, 4.377247e-07, 4.287297e-07, 4.452023e-07, 
    4.359355e-07, 4.306591e-07, 4.106622e-07, 4.063464e-07, 4.023673e-07, 
    3.945794e-07, 3.847192e-07, 3.677885e-07, 3.534381e-07, 3.406466e-07, 
    3.41574e-07, 3.412473e-07, 3.384262e-07, 3.454402e-07, 3.372834e-07, 
    3.359258e-07, 3.394817e-07, 3.191754e-07, 3.248965e-07, 3.19043e-07, 
    3.227599e-07, 4.251855e-07, 4.196977e-07, 4.226577e-07, 4.171015e-07, 
    4.210109e-07, 4.037939e-07, 3.987162e-07, 3.754747e-07, 3.849115e-07, 
    3.699616e-07, 3.833768e-07, 3.80978e-07, 3.694778e-07, 3.826447e-07, 
    3.542191e-07, 3.733412e-07, 3.383169e-07, 3.56879e-07, 3.371741e-07, 
    3.407013e-07, 3.348744e-07, 3.297085e-07, 3.232821e-07, 3.116319e-07, 
    3.143058e-07, 3.04719e-07, 4.115963e-07, 4.046239e-07, 4.052359e-07, 
    3.980104e-07, 3.92717e-07, 3.813929e-07, 3.636509e-07, 3.702621e-07, 
    3.581824e-07, 3.557869e-07, 3.741616e-07, 3.628112e-07, 3.999986e-07, 
    3.93839e-07, 3.975002e-07, 4.11043e-07, 3.687307e-07, 3.900954e-07, 
    3.512203e-07, 3.623656e-07, 3.304418e-07, 3.460878e-07, 3.157837e-07, 
    3.033579e-07, 2.919569e-07, 2.789823e-07, 4.008501e-07, 4.055531e-07, 
    3.971567e-07, 3.857132e-07, 3.752802e-07, 3.616794e-07, 3.603058e-07, 
    3.577979e-07, 3.513531e-07, 3.459901e-07, 3.570062e-07, 3.446539e-07, 
    3.924167e-07, 3.669115e-07, 4.073388e-07, 3.948927e-07, 3.863825e-07, 
    3.901029e-07, 3.710227e-07, 3.666105e-07, 3.490148e-07, 3.580444e-07, 
    3.063944e-07, 3.286225e-07, 2.693609e-07, 2.85163e-07, 4.072039e-07, 
    4.008668e-07, 3.792782e-07, 3.894595e-07, 3.60783e-07, 3.539301e-07, 
    3.484201e-07, 3.414531e-07, 3.407069e-07, 3.366262e-07, 3.433292e-07, 
    3.368897e-07, 3.616508e-07, 3.504507e-07, 3.817103e-07, 3.739497e-07, 
    3.775081e-07, 3.814343e-07, 3.693967e-07, 3.568308e-07, 3.565669e-07, 
    3.52596e-07, 3.415518e-07, 3.606696e-07, 3.035945e-07, 3.381104e-07, 
    3.940249e-07, 3.821117e-07, 3.804304e-07, 3.85006e-07, 3.546135e-07, 
    3.65448e-07, 3.367255e-07, 3.443444e-07, 3.319171e-07, 3.380566e-07, 
    3.389657e-07, 3.469684e-07, 3.520092e-07, 3.649465e-07, 3.756867e-07, 
    3.843406e-07, 3.823177e-07, 3.72849e-07, 3.560713e-07, 3.406387e-07, 
    3.439826e-07, 3.328515e-07, 3.62817e-07, 3.500552e-07, 3.549536e-07, 
    3.422702e-07, 3.704384e-07, 3.463595e-07, 3.767534e-07, 3.740257e-07, 
    3.656651e-07, 3.491988e-07, 3.456216e-07, 3.418246e-07, 3.441648e-07, 
    3.556518e-07, 3.575569e-07, 3.658673e-07, 3.681818e-07, 3.746187e-07, 
    3.799989e-07, 3.75081e-07, 3.699581e-07, 3.556476e-07, 3.430488e-07, 
    3.296351e-07, 3.264041e-07, 3.112472e-07, 3.23549e-07, 3.034085e-07, 
    3.204761e-07, 2.913074e-07, 3.449972e-07, 3.209901e-07, 3.65288e-07, 
    3.603441e-07, 3.515059e-07, 3.317514e-07, 3.423292e-07, 3.299799e-07, 
    3.576318e-07, 3.725241e-07, 3.764403e-07, 3.838107e-07, 3.762728e-07, 
    3.768826e-07, 3.69748e-07, 3.720317e-07, 3.551785e-07, 3.641714e-07, 
    3.389881e-07, 3.300767e-07, 3.057144e-07, 2.913619e-07, 2.77207e-07, 
    2.711018e-07, 2.692612e-07, 2.684941e-07,
  1.244258e-08, 1.172508e-08, 1.186215e-08, 1.130106e-08, 1.160987e-08, 
    1.1246e-08, 1.229463e-08, 1.169721e-08, 1.207609e-08, 1.237675e-08, 
    1.026804e-08, 1.12765e-08, 9.292962e-09, 9.883202e-09, 8.4509e-09, 
    9.383009e-09, 8.271684e-09, 8.476838e-09, 7.870791e-09, 8.040978e-09, 
    7.301955e-09, 7.793165e-09, 6.944861e-09, 7.417106e-09, 7.340821e-09, 
    7.809774e-09, 1.106801e-08, 1.03898e-08, 1.110917e-08, 1.101025e-08, 
    1.105457e-08, 1.160341e-08, 1.188738e-08, 1.249876e-08, 1.238611e-08, 
    1.193791e-08, 1.096599e-08, 1.128919e-08, 1.048789e-08, 1.050551e-08, 
    9.66256e-09, 1.003617e-08, 8.695928e-09, 9.062407e-09, 8.033821e-09, 
    8.283805e-09, 8.045425e-09, 8.117164e-09, 8.044493e-09, 8.413467e-09, 
    8.253857e-09, 8.584163e-09, 9.96539e-09, 9.54347e-09, 1.084239e-08, 
    1.168339e-08, 1.226795e-08, 1.269546e-08, 1.263438e-08, 1.25185e-08, 
    1.193532e-08, 1.140543e-08, 1.101333e-08, 1.075663e-08, 1.050804e-08, 
    9.781234e-09, 9.412111e-09, 8.623161e-09, 8.761801e-09, 8.527942e-09, 
    8.308992e-09, 7.950838e-09, 8.008983e-09, 7.854067e-09, 8.534089e-09, 
    8.077415e-09, 8.8415e-09, 8.627358e-09, 1.044097e-08, 1.120133e-08, 
    1.153632e-08, 1.18357e-08, 1.258755e-08, 1.206472e-08, 1.226889e-08, 
    1.17873e-08, 1.148854e-08, 1.163561e-08, 1.074967e-08, 1.108798e-08, 
    9.390562e-09, 1.00962e-08, 8.33431e-09, 8.733214e-09, 8.240767e-09, 
    8.489389e-09, 8.06674e-09, 8.446391e-09, 7.797005e-09, 7.660708e-09, 
    7.753649e-09, 7.40127e-09, 8.467816e-09, 8.045407e-09, 1.163974e-08, 
    1.161565e-08, 1.150394e-08, 1.200092e-08, 1.203184e-08, 1.250185e-08, 
    1.208301e-08, 1.190778e-08, 1.147141e-08, 1.121883e-08, 1.098256e-08, 
    1.047596e-08, 9.93075e-09, 9.204024e-09, 8.70693e-09, 8.385124e-09, 
    8.581389e-09, 8.407936e-09, 8.602003e-09, 8.694115e-09, 7.711553e-09, 
    8.252369e-09, 7.451194e-09, 7.493934e-09, 7.850403e-09, 7.48911e-09, 
    1.159876e-08, 1.173772e-08, 1.222957e-08, 1.18434e-08, 1.255383e-08, 
    1.215241e-08, 1.192587e-08, 1.108077e-08, 1.090121e-08, 1.073656e-08, 
    1.041681e-08, 1.00168e-08, 9.342679e-09, 8.784132e-09, 8.296393e-09, 
    8.331428e-09, 8.31908e-09, 8.212715e-09, 8.478042e-09, 8.169759e-09, 
    8.118837e-09, 8.252457e-09, 7.499672e-09, 7.70923e-09, 7.494845e-09, 
    7.630733e-09, 1.169242e-08, 1.145997e-08, 1.158515e-08, 1.135057e-08, 
    1.151545e-08, 1.079549e-08, 1.058624e-08, 9.646701e-09, 1.002455e-08, 
    9.428294e-09, 9.962755e-09, 9.866443e-09, 9.409209e-09, 9.933327e-09, 
    8.814223e-09, 9.561977e-09, 8.208601e-09, 8.916971e-09, 8.165657e-09, 
    8.298457e-09, 8.079472e-09, 7.887035e-09, 7.649894e-09, 7.226439e-09, 
    7.322887e-09, 6.979157e-09, 1.111977e-08, 1.082983e-08, 1.085518e-08, 
    1.055727e-08, 1.034084e-08, 9.883078e-09, 9.180416e-09, 9.440153e-09, 
    8.967472e-09, 8.874734e-09, 9.594524e-09, 9.147604e-09, 1.063895e-08, 
    1.038659e-08, 1.053634e-08, 1.109667e-08, 9.379765e-09, 1.023423e-08, 
    8.698879e-09, 9.13021e-09, 7.914255e-09, 8.502687e-09, 7.376386e-09, 
    6.935881e-09, 6.534466e-09, 6.088046e-09, 1.067401e-08, 1.086832e-08, 
    1.052226e-08, 1.005687e-08, 9.638969e-09, 9.103446e-09, 9.049954e-09, 
    8.952562e-09, 8.703975e-09, 8.498969e-09, 8.921894e-09, 8.448152e-09, 
    1.032861e-08, 9.308201e-09, 1.094241e-08, 1.042961e-08, 1.008389e-08, 
    1.023453e-08, 9.470193e-09, 9.29638e-09, 8.614384e-09, 8.962121e-09, 
    7.038812e-09, 7.846783e-09, 5.764294e-09, 6.299311e-09, 1.093681e-08, 
    1.067469e-08, 9.798391e-09, 1.020843e-08, 9.068525e-09, 8.803086e-09, 
    8.591647e-09, 8.32686e-09, 8.29867e-09, 8.145093e-09, 8.397881e-09, 
    8.154983e-09, 9.10233e-09, 8.669361e-09, 9.89581e-09, 9.586113e-09, 
    9.727693e-09, 9.884737e-09, 9.40601e-09, 8.915107e-09, 8.904894e-09, 
    8.751726e-09, 8.330587e-09, 9.064109e-09, 6.9443e-09, 8.200836e-09, 
    1.039417e-08, 9.911921e-09, 9.844498e-09, 1.002836e-08, 8.829431e-09, 
    9.25077e-09, 8.148819e-09, 8.436398e-09, 7.969109e-09, 8.198812e-09, 
    8.233019e-09, 8.536236e-09, 8.72917e-09, 9.231117e-09, 9.655136e-09, 
    1.000154e-08, 9.920192e-09, 9.542465e-09, 8.885727e-09, 8.296093e-09, 
    8.422664e-09, 8.003925e-09, 9.147833e-09, 8.654206e-09, 8.842555e-09, 
    8.357763e-09, 9.447114e-09, 8.513033e-09, 9.697608e-09, 9.589132e-09, 
    9.259282e-09, 8.621421e-09, 8.484944e-09, 8.340905e-09, 8.42958e-09, 
    8.869518e-09, 8.943223e-09, 9.267214e-09, 9.358154e-09, 9.612678e-09, 
    9.827223e-09, 9.631046e-09, 9.428154e-09, 8.869354e-09, 8.387253e-09, 
    7.884312e-09, 7.764785e-09, 7.212599e-09, 7.659689e-09, 6.937682e-09, 
    7.547137e-09, 6.511855e-09, 8.461198e-09, 7.565925e-09, 9.244499e-09, 
    9.051442e-09, 8.70984e-09, 7.962944e-09, 8.359996e-09, 7.897103e-09, 
    8.946125e-09, 9.529593e-09, 9.685133e-09, 9.980211e-09, 9.678463e-09, 
    9.702752e-09, 9.419866e-09, 9.510098e-09, 8.851235e-09, 9.200773e-09, 
    8.233863e-09, 7.900696e-09, 7.014576e-09, 6.51375e-09, 6.027837e-09, 
    5.822407e-09, 5.760973e-09, 5.735437e-09,
  8.582678e-11, 7.828047e-11, 7.970476e-11, 7.392763e-11, 7.708981e-11, 
    7.336845e-11, 8.425249e-11, 7.799186e-11, 8.194435e-11, 8.51252e-11, 
    6.367281e-11, 7.367799e-11, 5.447788e-11, 5.998542e-11, 4.694775e-11, 
    5.530623e-11, 4.53973e-11, 4.71737e-11, 4.199856e-11, 4.342949e-11, 
    3.734755e-11, 4.13518e-11, 3.139601e-11, 3.827231e-11, 3.76587e-11, 
    4.148987e-11, 7.157008e-11, 6.485486e-11, 7.198465e-11, 7.098976e-11, 
    7.143496e-11, 7.702316e-11, 7.996785e-11, 8.642695e-11, 8.522481e-11, 
    8.049552e-11, 7.054601e-11, 7.380693e-11, 6.581241e-11, 6.598491e-11, 
    5.790527e-11, 6.144223e-11, 4.909776e-11, 5.237694e-11, 4.336896e-11, 
    4.550157e-11, 4.346712e-11, 4.407578e-11, 4.345924e-11, 4.662235e-11, 
    4.524412e-11, 4.811279e-11, 6.076665e-11, 5.679303e-11, 6.931181e-11, 
    7.784891e-11, 8.396967e-11, 8.853893e-11, 8.78813e-11, 8.66382e-11, 
    8.046846e-11, 7.499148e-11, 7.102061e-11, 6.845973e-11, 6.600975e-11, 
    5.902097e-11, 5.557487e-11, 4.845566e-11, 4.968162e-11, 4.762003e-11, 
    4.571851e-11, 4.266939e-11, 4.315913e-11, 4.185889e-11, 4.767381e-11, 
    4.373816e-11, 5.039131e-11, 4.849262e-11, 6.535383e-11, 7.291567e-11, 
    7.63327e-11, 7.94293e-11, 8.737826e-11, 8.182478e-11, 8.397955e-11, 
    7.892596e-11, 7.584219e-11, 7.735525e-11, 6.839077e-11, 7.177111e-11, 
    5.537591e-11, 6.201713e-11, 4.593695e-11, 4.942794e-11, 4.513175e-11, 
    4.728318e-11, 4.364765e-11, 4.690851e-11, 4.138371e-11, 4.025689e-11, 
    4.1024e-11, 3.814463e-11, 4.709506e-11, 4.346698e-11, 7.739787e-11, 
    7.714935e-11, 7.600019e-11, 8.115515e-11, 8.147943e-11, 8.645996e-11, 
    8.201711e-11, 8.018079e-11, 7.566663e-11, 7.309298e-11, 7.0712e-11, 
    6.56957e-11, 6.043695e-11, 5.366401e-11, 4.919511e-11, 4.637651e-11, 
    4.808843e-11, 4.657434e-11, 4.826953e-11, 4.908172e-11, 4.067588e-11, 
    4.523133e-11, 3.854773e-11, 3.889411e-11, 4.182833e-11, 3.885495e-11, 
    7.697526e-11, 7.841147e-11, 8.356318e-11, 7.950945e-11, 8.701659e-11, 
    8.274808e-11, 8.036972e-11, 7.16986e-11, 6.989832e-11, 6.826086e-11, 
    6.511811e-11, 6.125702e-11, 5.493469e-11, 4.988011e-11, 4.560994e-11, 
    4.591206e-11, 4.58055e-11, 4.489129e-11, 4.71842e-11, 4.4524e-11, 
    4.409002e-11, 4.523209e-11, 3.89407e-11, 4.06567e-11, 3.89015e-11, 
    4.001065e-11, 7.794237e-11, 7.554946e-11, 7.683507e-11, 7.443168e-11, 
    7.611833e-11, 6.884544e-11, 6.677724e-11, 5.775673e-11, 6.133107e-11, 
    5.572445e-11, 6.074154e-11, 5.982654e-11, 5.554806e-11, 6.046146e-11, 
    5.014802e-11, 5.696539e-11, 4.485607e-11, 5.106664e-11, 4.448899e-11, 
    4.562772e-11, 4.375561e-11, 4.213437e-11, 4.016799e-11, 3.674581e-11, 
    3.7515e-11, 3.480201e-11, 7.209158e-11, 6.918685e-11, 6.943919e-11, 
    6.649253e-11, 6.437874e-11, 5.998425e-11, 5.344869e-11, 5.583415e-11, 
    5.15203e-11, 5.06883e-11, 5.726894e-11, 5.314993e-11, 6.729627e-11, 
    6.48236e-11, 6.628713e-11, 7.185869e-11, 5.527632e-11, 6.33459e-11, 
    4.912387e-11, 5.299179e-11, 4.236232e-11, 4.739926e-11, 3.79443e-11, 
    3.134359e-11, 2.901295e-11, 2.645106e-11, 6.764215e-11, 6.957015e-11, 
    6.614904e-11, 6.164026e-11, 5.768435e-11, 5.274879e-11, 5.226428e-11, 
    5.138621e-11, 4.916896e-11, 4.73668e-11, 5.11108e-11, 4.692384e-11, 
    6.425994e-11, 5.461776e-11, 7.031006e-11, 6.524296e-11, 6.189911e-11, 
    6.334884e-11, 5.611237e-11, 5.450924e-11, 4.837842e-11, 5.147216e-11, 
    3.526716e-11, 4.179812e-11, 2.461437e-11, 2.765936e-11, 7.025399e-11, 
    6.764892e-11, 5.918287e-11, 6.309679e-11, 5.243231e-11, 5.004881e-11, 
    4.817852e-11, 4.587263e-11, 4.562956e-11, 4.43136e-11, 4.64871e-11, 
    4.439791e-11, 5.273867e-11, 4.886298e-11, 6.010504e-11, 5.719045e-11, 
    5.851671e-11, 5.999998e-11, 5.551852e-11, 5.104991e-11, 5.095836e-11, 
    4.959217e-11, 4.59048e-11, 5.239235e-11, 3.139274e-11, 4.478961e-11, 
    6.489746e-11, 6.025801e-11, 5.961871e-11, 6.136749e-11, 5.028361e-11, 
    5.409125e-11, 4.434536e-11, 4.682159e-11, 4.282306e-11, 4.47723e-11, 
    4.506529e-11, 4.769261e-11, 4.939209e-11, 5.391149e-11, 5.783572e-11, 
    6.111138e-11, 6.03366e-11, 5.678368e-11, 5.078667e-11, 4.560736e-11, 
    4.670223e-11, 4.311644e-11, 5.315201e-11, 4.872924e-11, 5.040073e-11, 
    4.613964e-11, 5.589858e-11, 4.748966e-11, 5.823401e-11, 5.721862e-11, 
    5.416917e-11, 4.844034e-11, 4.72444e-11, 4.599391e-11, 4.676231e-11, 
    5.064164e-11, 5.130229e-11, 5.424182e-11, 5.507715e-11, 5.743849e-11, 
    5.94553e-11, 5.761023e-11, 5.572316e-11, 5.064018e-11, 4.639495e-11, 
    4.211159e-11, 4.111628e-11, 3.663593e-11, 4.024851e-11, 3.13541e-11, 
    3.932692e-11, 2.888241e-11, 4.703741e-11, 3.94802e-11, 5.403386e-11, 
    5.227774e-11, 4.922086e-11, 4.277118e-11, 4.615896e-11, 4.221863e-11, 
    5.132836e-11, 5.666392e-11, 5.811693e-11, 6.090789e-11, 5.805436e-11, 
    5.828232e-11, 5.564653e-11, 5.64827e-11, 5.047825e-11, 5.363433e-11, 
    4.507253e-11, 4.224871e-11, 3.507789e-11, 2.889335e-11, 2.610809e-11, 
    2.494268e-11, 2.459563e-11, 2.445157e-11,
  8.2723e-14, 7.054447e-14, 7.281189e-14, 6.371174e-14, 6.866073e-14, 
    6.284501e-14, 8.014966e-14, 7.008687e-14, 7.640725e-14, 8.157414e-14, 
    4.825941e-14, 6.332449e-14, 3.5329e-14, 4.295663e-14, 2.556488e-14, 
    3.645209e-14, 2.366503e-14, 2.584516e-14, 1.965235e-14, 2.131524e-14, 
    1.454314e-14, 1.891407e-14, 1.164344e-14, 1.552043e-14, 1.48697e-14, 
    1.907097e-14, 6.007536e-14, 4.998971e-14, 6.07114e-14, 5.918752e-14, 
    5.986838e-14, 6.855561e-14, 7.323237e-14, 8.370835e-14, 8.173707e-14, 
    7.407721e-14, 5.851062e-14, 6.352444e-14, 5.140173e-14, 5.165706e-14, 
    4.003241e-14, 4.503399e-14, 2.826554e-14, 3.252167e-14, 2.124409e-14, 
    2.379149e-14, 2.13595e-14, 2.207914e-14, 2.135022e-14, 2.516274e-14, 
    2.34796e-14, 2.701905e-14, 4.406769e-14, 3.848998e-14, 5.663715e-14, 
    6.986045e-14, 7.968913e-14, 8.719429e-14, 8.610579e-14, 8.405573e-14, 
    7.403384e-14, 6.53678e-14, 5.923463e-14, 5.535177e-14, 5.169384e-14, 
    4.159456e-14, 3.681823e-14, 2.745121e-14, 2.901158e-14, 2.640129e-14, 
    2.405521e-14, 2.042695e-14, 2.099801e-14, 1.949221e-14, 2.646852e-14, 
    2.16791e-14, 2.992542e-14, 2.74979e-14, 5.072436e-14, 6.214511e-14, 
    6.746859e-14, 7.237219e-14, 8.5275e-14, 7.621438e-14, 7.97052e-14, 
    7.15702e-14, 6.669865e-14, 6.907974e-14, 5.524803e-14, 6.038359e-14, 
    3.654697e-14, 4.586022e-14, 2.43216e-14, 2.868679e-14, 2.334384e-14, 
    2.598126e-14, 2.157221e-14, 2.551629e-14, 1.895029e-14, 1.76839e-14, 
    1.854315e-14, 1.53843e-14, 2.574752e-14, 2.135932e-14, 6.914708e-14, 
    6.875467e-14, 6.694645e-14, 7.513619e-14, 7.565793e-14, 8.376261e-14, 
    7.652465e-14, 7.357306e-14, 6.642351e-14, 6.241899e-14, 5.876362e-14, 
    5.122914e-14, 4.359796e-14, 3.423437e-14, 2.838956e-14, 2.486011e-14, 
    2.698842e-14, 2.510356e-14, 2.721637e-14, 2.824512e-14, 1.815168e-14, 
    2.346414e-14, 1.581537e-14, 1.618878e-14, 1.945721e-14, 1.614643e-14, 
    6.848009e-14, 7.075239e-14, 7.902817e-14, 7.250008e-14, 8.46787e-14, 
    7.770624e-14, 7.387562e-14, 6.027236e-14, 5.752573e-14, 5.505273e-14, 
    5.037699e-14, 4.476858e-14, 3.594725e-14, 2.926639e-14, 2.392314e-14, 
    2.429121e-14, 2.416119e-14, 2.305407e-14, 2.58582e-14, 2.261348e-14, 
    2.209606e-14, 2.346506e-14, 1.623921e-14, 1.813018e-14, 1.619678e-14, 
    1.741074e-14, 7.000847e-14, 6.624005e-14, 6.825913e-14, 6.449523e-14, 
    6.713187e-14, 5.59328e-14, 5.283358e-14, 3.982556e-14, 4.487465e-14, 
    3.70225e-14, 4.403189e-14, 4.273151e-14, 3.678165e-14, 4.363285e-14, 
    2.961128e-14, 3.872802e-14, 2.301172e-14, 3.080198e-14, 2.257161e-14, 
    2.394476e-14, 2.169972e-14, 1.980845e-14, 1.758512e-14, 1.391827e-14, 
    1.47186e-14, 1.19624e-14, 6.087569e-14, 5.644823e-14, 5.682987e-14, 
    5.241011e-14, 4.929106e-14, 4.295497e-14, 3.394626e-14, 3.717249e-14, 
    3.13946e-14, 3.031007e-14, 3.914812e-14, 3.354755e-14, 5.360756e-14, 
    4.994378e-14, 5.210509e-14, 6.051798e-14, 3.641138e-14, 4.778343e-14, 
    2.829878e-14, 3.3337e-14, 2.007127e-14, 2.61258e-14, 1.517148e-14, 
    1.157616e-14, 8.760279e-15, 6.080912e-15, 5.412476e-14, 5.702817e-14, 
    5.190026e-14, 4.531819e-14, 3.972485e-14, 3.301414e-14, 3.237286e-14, 
    3.121913e-14, 2.835623e-14, 2.608536e-14, 3.085954e-14, 2.553527e-14, 
    4.911708e-14, 3.551802e-14, 5.81514e-14, 5.056091e-14, 4.569031e-14, 
    4.778769e-14, 3.755357e-14, 3.537136e-14, 2.735369e-14, 3.133157e-14, 
    1.242146e-14, 1.942265e-14, 4.446216e-15, 7.288357e-15, 5.806611e-14, 
    5.41349e-14, 4.182246e-14, 4.742145e-14, 3.259488e-14, 2.948344e-14, 
    2.710175e-14, 2.424307e-14, 2.394698e-14, 2.236219e-14, 2.499612e-14, 
    2.246279e-14, 3.300072e-14, 2.796704e-14, 4.31263e-14, 3.903938e-14, 
    4.08867e-14, 4.297727e-14, 3.674135e-14, 3.07802e-14, 3.066099e-14, 
    2.889694e-14, 2.428234e-14, 3.254204e-14, 1.163922e-14, 2.293185e-14, 
    5.005235e-14, 4.334353e-14, 4.243748e-14, 4.492684e-14, 2.978625e-14, 
    3.480789e-14, 2.240007e-14, 2.540876e-14, 2.060564e-14, 2.291106e-14, 
    2.326364e-14, 2.649203e-14, 2.864098e-14, 3.456628e-14, 3.993552e-14, 
    4.456014e-14, 4.345522e-14, 3.847708e-14, 3.043777e-14, 2.392e-14, 
    2.526129e-14, 2.094805e-14, 3.355032e-14, 2.779737e-14, 2.993759e-14, 
    2.456951e-14, 3.726065e-14, 2.62385e-14, 4.049117e-14, 3.90784e-14, 
    3.491276e-14, 2.743186e-14, 2.593302e-14, 2.439119e-14, 2.533549e-14, 
    3.024955e-14, 3.110944e-14, 3.50106e-14, 3.614061e-14, 3.938326e-14, 
    4.220663e-14, 3.962179e-14, 3.702073e-14, 3.024766e-14, 2.488279e-14, 
    1.978224e-14, 1.864734e-14, 1.380513e-14, 1.767458e-14, 1.158963e-14, 
    1.665917e-14, 8.612961e-15, 2.5676e-14, 1.682676e-14, 3.473071e-14, 
    3.239063e-14, 2.842239e-14, 2.054526e-14, 2.459317e-14, 1.990548e-14, 
    3.11435e-14, 3.831191e-14, 4.032763e-14, 4.42693e-14, 4.024032e-14, 
    4.05587e-14, 3.691606e-14, 3.806233e-14, 3.003788e-14, 3.419462e-14, 
    2.327238e-14, 1.994016e-14, 1.223397e-14, 8.625269e-15, 5.757012e-15, 
    4.720195e-15, 4.430813e-15, 4.313349e-15,
  2.795984e-19, 2.389544e-19, 2.465295e-19, 2.161035e-19, 2.326581e-19, 
    2.132022e-19, 2.710187e-19, 2.374251e-19, 2.585334e-19, 2.757686e-19, 
    1.642776e-19, 2.148073e-19, 1.207162e-19, 1.464373e-19, 8.767294e-20, 
    1.245082e-19, 8.122402e-20, 8.86237e-20, 6.757771e-20, 7.323728e-20, 
    5.014306e-20, 6.506282e-20, 4.024981e-20, 5.348385e-20, 5.125973e-20, 
    6.559737e-20, 2.039268e-19, 1.700923e-19, 2.060575e-19, 2.009522e-19, 
    2.032334e-19, 2.323067e-19, 2.479338e-19, 2.828825e-19, 2.763118e-19, 
    2.507551e-19, 1.986837e-19, 2.154766e-19, 1.748351e-19, 1.756925e-19, 
    1.365854e-19, 1.5343e-19, 9.682819e-20, 1.112307e-19, 7.299526e-20, 
    8.16535e-20, 7.338784e-20, 7.583507e-20, 7.33563e-20, 8.63085e-20, 
    8.059417e-20, 9.260425e-20, 1.501779e-19, 1.313845e-19, 1.924032e-19, 
    2.366684e-19, 2.694828e-19, 2.944958e-19, 2.908703e-19, 2.840401e-19, 
    2.506103e-19, 2.216452e-19, 2.0111e-19, 1.880924e-19, 1.75816e-19, 
    1.418497e-19, 1.25744e-19, 9.4069e-20, 9.935494e-20, 9.05098e-20, 
    8.254905e-20, 7.021485e-20, 7.215811e-20, 6.703231e-20, 9.07378e-20, 
    7.447481e-20, 1.024487e-19, 9.422726e-20, 1.725601e-19, 2.108589e-19, 
    2.286721e-19, 2.450608e-19, 2.881027e-19, 2.578897e-19, 2.695364e-19, 
    2.423816e-19, 2.260972e-19, 2.340589e-19, 1.877444e-19, 2.049594e-19, 
    1.248285e-19, 1.562098e-19, 8.34535e-20, 9.825504e-20, 8.013299e-20, 
    8.908536e-20, 7.411132e-20, 8.750808e-20, 6.518623e-20, 6.086921e-20, 
    6.379878e-20, 5.301866e-20, 8.82925e-20, 7.338724e-20, 2.34284e-19, 
    2.329722e-19, 2.26926e-19, 2.542907e-19, 2.560324e-19, 2.830633e-19, 
    2.589252e-19, 2.490716e-19, 2.251769e-19, 2.117759e-19, 1.995316e-19, 
    1.742555e-19, 1.485967e-19, 1.170186e-19, 9.724828e-20, 8.528148e-20, 
    9.250042e-20, 8.610767e-20, 9.327311e-20, 9.675901e-20, 6.246432e-20, 
    8.054165e-20, 5.44915e-20, 5.576684e-20, 6.69131e-20, 5.56222e-20, 
    2.320542e-19, 2.396491e-19, 2.672782e-19, 2.454879e-19, 2.86116e-19, 
    2.628681e-19, 2.500819e-19, 2.045868e-19, 1.953825e-19, 1.870893e-19, 
    1.713933e-19, 1.525369e-19, 1.228039e-19, 1.002177e-19, 8.210056e-20, 
    8.335032e-20, 8.290891e-20, 7.914858e-20, 8.866795e-20, 7.765139e-20, 
    7.589257e-20, 8.054479e-20, 5.593904e-20, 6.239103e-20, 5.579415e-20, 
    5.993746e-20, 2.371631e-19, 2.245633e-19, 2.313155e-19, 2.187256e-19, 
    2.275461e-19, 1.900412e-19, 1.796425e-19, 1.358881e-19, 1.528938e-19, 
    1.264334e-19, 1.500574e-19, 1.456792e-19, 1.256206e-19, 1.487141e-19, 
    1.013854e-19, 1.321873e-19, 7.900467e-20, 1.054149e-19, 7.750906e-20, 
    8.217398e-20, 7.454495e-20, 6.810926e-20, 6.053232e-20, 4.800538e-20, 
    5.074307e-20, 4.130545e-20, 2.066078e-19, 1.917698e-19, 1.930495e-19, 
    1.782209e-19, 1.677448e-19, 1.464317e-19, 1.160451e-19, 1.269396e-19, 
    1.074196e-19, 1.037505e-19, 1.33604e-19, 1.146978e-19, 1.822403e-19, 
    1.69938e-19, 1.771969e-19, 2.054096e-19, 1.243708e-19, 1.626775e-19, 
    9.694079e-20, 1.139864e-19, 6.900412e-20, 8.957556e-20, 5.229133e-20, 
    4.001881e-20, 3.033257e-20, 2.107736e-20, 1.839759e-19, 1.937143e-19, 
    1.765091e-19, 1.543863e-19, 1.355486e-19, 1.128953e-19, 1.107276e-19, 
    1.068261e-19, 9.713539e-20, 8.943841e-20, 1.056097e-19, 8.757247e-20, 
    1.671602e-19, 1.213546e-19, 1.974798e-19, 1.720111e-19, 1.556382e-19, 
    1.626918e-19, 1.282255e-19, 1.208593e-19, 9.373849e-20, 1.072064e-19, 
    4.287924e-20, 6.679538e-20, 1.540594e-20, 2.525344e-20, 1.971939e-19, 
    1.840099e-19, 1.426174e-19, 1.614605e-19, 1.114781e-19, 1.009526e-19, 
    9.288458e-20, 8.31869e-20, 8.218154e-20, 7.679727e-20, 8.574306e-20, 
    7.713923e-20, 1.128499e-19, 9.581691e-20, 1.470087e-19, 1.332374e-19, 
    1.394647e-19, 1.465068e-19, 1.254846e-19, 1.053412e-19, 1.049379e-19, 
    9.896672e-20, 8.332021e-20, 1.112995e-19, 4.023534e-20, 7.873328e-20, 
    1.703027e-19, 1.477401e-19, 1.44689e-19, 1.530694e-19, 1.019776e-19, 
    1.189562e-19, 7.692603e-20, 8.714326e-20, 7.082299e-20, 7.866265e-20, 
    7.986057e-20, 9.08175e-20, 9.809986e-20, 1.1814e-19, 1.362588e-19, 
    1.518354e-19, 1.481161e-19, 1.31341e-19, 1.041826e-19, 8.20899e-20, 
    8.664288e-20, 7.198813e-20, 1.147072e-19, 9.524205e-20, 1.024899e-19, 
    8.429511e-20, 1.272371e-19, 8.995779e-20, 1.381317e-19, 1.333689e-19, 
    1.193104e-19, 9.400343e-20, 8.892175e-20, 8.368978e-20, 8.689466e-20, 
    1.035457e-19, 1.064551e-19, 1.196409e-19, 1.234567e-19, 1.343969e-19, 
    1.439115e-19, 1.352011e-19, 1.264275e-19, 1.035393e-19, 8.535843e-20, 
    6.802002e-20, 6.415389e-20, 4.76182e-20, 6.083743e-20, 4.006507e-20, 
    5.737281e-20, 2.982477e-20, 8.804988e-20, 5.794484e-20, 1.186955e-19, 
    1.107876e-19, 9.73595e-20, 7.061751e-20, 8.437541e-20, 6.843964e-20, 
    1.065703e-19, 1.307838e-19, 1.375805e-19, 1.508565e-19, 1.372862e-19, 
    1.383592e-19, 1.260742e-19, 1.29942e-19, 1.028293e-19, 1.168843e-19, 
    7.989026e-20, 6.855773e-20, 4.223658e-20, 2.98672e-20, 1.995537e-20, 
    1.635812e-20, 1.535239e-20, 1.494392e-20,
  2.052293e-25, 1.75542e-25, 1.810767e-25, 1.588413e-25, 1.709412e-25, 
    1.567203e-25, 1.989642e-25, 1.744246e-25, 1.898456e-25, 2.024328e-25, 
    1.209308e-25, 1.578937e-25, 8.901889e-26, 1.078676e-25, 6.476819e-26, 
    9.179894e-26, 6.002975e-26, 6.546661e-26, 4.999551e-26, 5.415835e-26, 
    3.715747e-26, 4.814505e-26, 2.987048e-26, 3.961935e-26, 3.798048e-26, 
    4.853842e-26, 1.499385e-25, 1.251869e-25, 1.514965e-25, 1.477633e-25, 
    1.494315e-25, 1.706843e-25, 1.821027e-25, 2.076272e-25, 2.028294e-25, 
    1.841637e-25, 1.461044e-25, 1.58383e-25, 1.286578e-25, 1.292853e-25, 
    1.006503e-25, 1.129888e-25, 7.149181e-26, 8.206204e-26, 5.398038e-26, 
    6.034538e-26, 5.426907e-26, 5.606849e-26, 5.424587e-26, 6.376581e-26, 
    5.956684e-26, 6.83902e-26, 1.106073e-25, 9.68391e-26, 1.415109e-25, 
    1.738717e-25, 1.978426e-25, 2.161057e-25, 2.13459e-25, 2.084724e-25, 
    1.84058e-25, 1.628923e-25, 1.478787e-25, 1.383576e-25, 1.293756e-25, 
    1.045071e-25, 9.270489e-26, 6.946585e-26, 7.334683e-26, 6.685199e-26, 
    6.10035e-26, 5.193548e-26, 5.336473e-26, 4.959424e-26, 6.701944e-26, 
    5.506835e-26, 7.561774e-26, 6.958206e-26, 1.26993e-25, 1.550071e-25, 
    1.680282e-25, 1.800037e-25, 2.114385e-25, 1.893754e-25, 1.978818e-25, 
    1.780462e-25, 1.661462e-25, 1.719648e-25, 1.38103e-25, 1.506936e-25, 
    9.203373e-26, 1.150243e-25, 6.166813e-26, 7.253937e-26, 5.922789e-26, 
    6.580571e-26, 5.480107e-26, 6.464708e-26, 4.823587e-26, 4.505843e-26, 
    4.721481e-26, 3.92766e-26, 6.522332e-26, 5.426863e-26, 1.721293e-25, 
    1.711707e-25, 1.66752e-25, 1.867465e-25, 1.880188e-25, 2.077592e-25, 
    1.901318e-25, 1.829339e-25, 1.654736e-25, 1.556775e-25, 1.467244e-25, 
    1.282337e-25, 1.094492e-25, 8.630758e-26, 7.180023e-26, 6.301127e-26, 
    6.831396e-26, 6.361827e-26, 6.888139e-26, 7.144102e-26, 4.623263e-26, 
    5.952825e-26, 4.036171e-26, 4.130116e-26, 4.950653e-26, 4.119463e-26, 
    1.704998e-25, 1.760497e-25, 1.962326e-25, 1.803158e-25, 2.09988e-25, 
    1.930117e-25, 1.83672e-25, 1.504211e-25, 1.4369e-25, 1.376238e-25, 
    1.261391e-25, 1.123348e-25, 9.05495e-26, 7.398018e-26, 6.067392e-26, 
    6.159231e-26, 6.126795e-26, 5.850433e-26, 6.549911e-26, 5.740379e-26, 
    5.611076e-26, 5.953055e-26, 4.1428e-26, 4.617868e-26, 4.132128e-26, 
    4.437246e-26, 1.742332e-25, 1.650251e-25, 1.6996e-25, 1.607581e-25, 
    1.672052e-25, 1.397832e-25, 1.321756e-25, 1.001393e-25, 1.125962e-25, 
    9.321025e-26, 1.10519e-25, 1.073124e-25, 9.261439e-26, 1.095352e-25, 
    7.483727e-26, 9.742745e-26, 5.839856e-26, 7.779473e-26, 5.729916e-26, 
    6.072787e-26, 5.511992e-26, 5.038657e-26, 4.481041e-26, 3.558164e-26, 
    3.75997e-26, 3.063965e-26, 1.518989e-25, 1.410475e-25, 1.419836e-25, 
    1.311354e-25, 1.234687e-25, 1.078635e-25, 8.559366e-26, 9.358128e-26, 
    7.92658e-26, 7.657321e-26, 9.846566e-26, 8.460549e-26, 1.340763e-25, 
    1.250739e-25, 1.303861e-25, 1.510228e-25, 9.169822e-26, 1.197595e-25, 
    7.157448e-26, 8.408362e-26, 5.104488e-26, 6.616579e-26, 3.874068e-26, 
    2.969992e-26, 2.254176e-26, 1.568702e-26, 1.353461e-25, 1.424699e-25, 
    1.298829e-25, 1.13689e-25, 9.989056e-26, 8.328323e-26, 8.169294e-26, 
    7.88303e-26, 7.171735e-26, 6.606505e-26, 7.793764e-26, 6.469438e-26, 
    1.230408e-25, 8.948692e-26, 1.452238e-25, 1.265912e-25, 1.146058e-25, 
    1.1977e-25, 9.452383e-26, 8.912378e-26, 6.922315e-26, 7.910938e-26, 
    3.180095e-26, 4.941992e-26, 1.147616e-26, 1.878227e-26, 1.450148e-25, 
    1.35371e-25, 1.050696e-25, 1.188685e-25, 8.224361e-26, 7.451959e-26, 
    6.859607e-26, 6.147223e-26, 6.073343e-26, 5.677589e-26, 6.33504e-26, 
    5.702728e-26, 8.324993e-26, 7.07493e-26, 1.082861e-25, 9.819695e-26, 
    1.027598e-25, 1.079186e-25, 9.25147e-26, 7.774065e-26, 7.744464e-26, 
    7.306183e-26, 6.157019e-26, 8.211256e-26, 2.98598e-26, 5.819908e-26, 
    1.253409e-25, 1.088218e-25, 1.06587e-25, 1.127248e-25, 7.5272e-26, 
    8.772835e-26, 5.687054e-26, 6.437907e-26, 5.238279e-26, 5.814716e-26, 
    5.902766e-26, 6.707798e-26, 7.242544e-26, 8.712988e-26, 1.00411e-25, 
    1.118211e-25, 1.090972e-25, 9.680719e-26, 7.689035e-26, 6.066608e-26, 
    6.401148e-26, 5.323972e-26, 8.461236e-26, 7.032721e-26, 7.564798e-26, 
    6.228653e-26, 9.379935e-26, 6.644654e-26, 1.017832e-25, 9.829336e-26, 
    8.798811e-26, 6.94177e-26, 6.568554e-26, 6.184175e-26, 6.419645e-26, 
    7.64229e-26, 7.855802e-26, 8.823041e-26, 9.10281e-26, 9.904666e-26, 
    1.060175e-25, 9.963597e-26, 9.320588e-26, 7.64182e-26, 6.30678e-26, 
    5.032092e-26, 4.747616e-26, 3.529618e-26, 4.503504e-26, 2.973408e-26, 
    4.248398e-26, 2.21661e-26, 6.504509e-26, 4.290524e-26, 8.753718e-26, 
    8.173703e-26, 7.188189e-26, 5.223165e-26, 6.234554e-26, 5.062963e-26, 
    7.864257e-26, 9.63989e-26, 1.013794e-25, 1.111042e-25, 1.011637e-25, 
    1.0195e-25, 9.294693e-26, 9.578188e-26, 7.589712e-26, 8.620909e-26, 
    5.904949e-26, 5.07165e-26, 3.132677e-26, 2.219749e-26, 1.485471e-26, 
    1.218381e-26, 1.143635e-26, 1.113267e-26,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.01045852, 0.01047329, 0.01047041, 0.01048232, 0.0104757, 0.01048351, 
    0.0104615, 0.01047388, 0.01046597, 0.01045983, 0.01050541, 0.01048285, 
    0.01052862, 0.01051432, 0.01055015, 0.01052642, 0.01055492, 0.01054943, 
    0.01056585, 0.01056115, 0.01058216, 0.01056802, 0.01059297, 0.01057877, 
    0.010581, 0.01056755, 0.01048736, 0.01050261, 0.01048646, 0.01048864, 
    0.01048766, 0.01047585, 0.01046992, 0.01045737, 0.01045964, 0.01046884, 
    0.01048962, 0.01048255, 0.01050028, 0.01049988, 0.01051958, 0.01051071, 
    0.0105437, 0.01053434, 0.01056134, 0.01055457, 0.01056103, 0.01055907, 
    0.01056106, 0.01055111, 0.01055538, 0.01054661, 0.01051238, 0.01052247, 
    0.01049234, 0.0104742, 0.01046205, 0.01045344, 0.01045466, 0.01045698, 
    0.0104689, 0.01048005, 0.01048855, 0.01049423, 0.01049982, 0.01051679, 
    0.01052569, 0.01054561, 0.010542, 0.0105481, 0.01055389, 0.01056364, 
    0.01056203, 0.01056632, 0.01054792, 0.01056017, 0.01053994, 0.01054548, 
    0.01050145, 0.01048446, 0.01047731, 0.01047097, 0.0104556, 0.01046622, 
    0.01046204, 0.01047196, 0.01047828, 0.01047515, 0.01049439, 0.01048692, 
    0.01052622, 0.01050932, 0.01055322, 0.01054274, 0.01055572, 0.01054909, 
    0.01056046, 0.01055023, 0.01056791, 0.01057177, 0.01056914, 0.01057921, 
    0.01054967, 0.01056104, 0.01047507, 0.01047558, 0.01047795, 0.01046754, 
    0.0104669, 0.01045731, 0.01046583, 0.01046946, 0.01047864, 0.01048408, 
    0.01048924, 0.01050056, 0.01051321, 0.01053081, 0.01054342, 0.01055186, 
    0.01054668, 0.01055125, 0.01054614, 0.01054374, 0.01057033, 0.01055542, 
    0.01057776, 0.01057652, 0.01056643, 0.01057666, 0.01047594, 0.010473, 
    0.01046283, 0.01047079, 0.01045626, 0.01046441, 0.0104691, 0.0104871, 
    0.01049102, 0.01049469, 0.01050191, 0.01051116, 0.01052738, 0.01054143, 
    0.01055422, 0.01055329, 0.01055362, 0.01055648, 0.0105494, 0.01055764, 
    0.01055904, 0.01055541, 0.01057636, 0.01057038, 0.0105765, 0.0105726, 
    0.01047395, 0.01047889, 0.01047622, 0.01048124, 0.01047771, 0.0104934, 
    0.0104981, 0.01051999, 0.01051099, 0.01052528, 0.01051243, 0.01051472, 
    0.01052579, 0.01051312, 0.01054068, 0.01052205, 0.01055659, 0.01053808, 
    0.01055775, 0.01055417, 0.01056009, 0.0105654, 0.01057206, 0.01058436, 
    0.01058151, 0.01059176, 0.01048623, 0.01049262, 0.01049204, 0.01049871, 
    0.01050365, 0.01051431, 0.01053139, 0.01052497, 0.01053673, 0.0105391, 
    0.01052121, 0.01053222, 0.01049689, 0.01050263, 0.0104992, 0.01048674, 
    0.01052647, 0.01050613, 0.01054363, 0.01053264, 0.01056465, 0.01054877, 
    0.01057994, 0.01059327, 0.0106057, 0.01062029, 0.01049609, 0.01049175, 
    0.0104995, 0.01051025, 0.01052015, 0.01053332, 0.01053465, 0.01053712, 
    0.01054349, 0.01054884, 0.01053792, 0.01055018, 0.010504, 0.01052823, 
    0.01049013, 0.01050165, 0.01050961, 0.0105061, 0.01052423, 0.0105285, 
    0.01054584, 0.01053687, 0.01059, 0.01056655, 0.01063131, 0.0106133, 
    0.01049024, 0.01049607, 0.01051634, 0.0105067, 0.01053418, 0.01054094, 
    0.01054641, 0.01055342, 0.01055417, 0.01055832, 0.01055152, 0.01055804, 
    0.01053334, 0.01054439, 0.010514, 0.01052142, 0.010518, 0.01051427, 
    0.0105258, 0.0105381, 0.01053833, 0.01054227, 0.01055343, 0.01053429, 
    0.01059308, 0.0105569, 0.01050242, 0.01051366, 0.01051523, 0.01051088, 
    0.01054026, 0.01052964, 0.01055821, 0.0105505, 0.01056312, 0.01055685, 
    0.01055593, 0.01054786, 0.01054284, 0.01053013, 0.01051976, 0.01051151, 
    0.01051343, 0.01052249, 0.01053884, 0.01055425, 0.01055088, 0.01056217, 
    0.01053219, 0.0105448, 0.01053994, 0.01055259, 0.0105248, 0.01054857, 
    0.01051873, 0.01052134, 0.01052943, 0.01054567, 0.01054921, 0.01055305, 
    0.01055067, 0.01053925, 0.01053736, 0.01052922, 0.01052699, 0.01052077, 
    0.01051563, 0.01052033, 0.01052528, 0.01053924, 0.01055182, 0.01056549, 
    0.01056881, 0.01058482, 0.01057184, 0.01059329, 0.01057512, 0.0106065, 
    0.0105499, 0.01057452, 0.01052978, 0.01053461, 0.01054337, 0.01056334, 
    0.01055253, 0.01056515, 0.01053728, 0.01052282, 0.01051903, 0.01051202, 
    0.01051919, 0.0105186, 0.01052546, 0.01052325, 0.0105397, 0.01053087, 
    0.01055592, 0.01056504, 0.0105907, 0.01060639, 0.01062227, 0.01062928, 
    0.01063141, 0.0106323,
  3.330992e-05, 3.340029e-05, 3.338268e-05, 3.345574e-05, 3.34151e-05, 
    3.346307e-05, 3.332817e-05, 3.340394e-05, 3.335553e-05, 3.331795e-05, 
    3.359839e-05, 3.345899e-05, 3.37422e-05, 3.365358e-05, 3.387577e-05, 
    3.372852e-05, 3.390539e-05, 3.387134e-05, 3.397334e-05, 3.394412e-05, 
    3.407483e-05, 3.398682e-05, 3.414221e-05, 3.405372e-05, 3.406765e-05, 
    3.398395e-05, 3.348689e-05, 3.358111e-05, 3.348134e-05, 3.349478e-05, 
    3.348871e-05, 3.3416e-05, 3.337963e-05, 3.330289e-05, 3.331679e-05, 
    3.337309e-05, 3.350081e-05, 3.345719e-05, 3.356673e-05, 3.356425e-05, 
    3.368618e-05, 3.363123e-05, 3.383577e-05, 3.377764e-05, 3.394534e-05, 
    3.390322e-05, 3.394339e-05, 3.393119e-05, 3.394355e-05, 3.388177e-05, 
    3.390825e-05, 3.385381e-05, 3.364156e-05, 3.370405e-05, 3.351764e-05, 
    3.340589e-05, 3.333152e-05, 3.327885e-05, 3.328631e-05, 3.330054e-05, 
    3.337342e-05, 3.344176e-05, 3.349423e-05, 3.352934e-05, 3.35639e-05, 
    3.366889e-05, 3.372401e-05, 3.384761e-05, 3.382516e-05, 3.386306e-05, 
    3.389902e-05, 3.395959e-05, 3.39496e-05, 3.397631e-05, 3.386194e-05, 
    3.393802e-05, 3.38124e-05, 3.384681e-05, 3.357392e-05, 3.346893e-05, 
    3.342491e-05, 3.338609e-05, 3.329204e-05, 3.335703e-05, 3.333143e-05, 
    3.33922e-05, 3.343087e-05, 3.341172e-05, 3.35303e-05, 3.348416e-05, 
    3.372728e-05, 3.362264e-05, 3.389483e-05, 3.382975e-05, 3.39104e-05, 
    3.386923e-05, 3.393981e-05, 3.387629e-05, 3.398619e-05, 3.401018e-05, 
    3.399381e-05, 3.405648e-05, 3.387278e-05, 3.394345e-05, 3.341121e-05, 
    3.341434e-05, 3.342884e-05, 3.33651e-05, 3.336117e-05, 3.330253e-05, 
    3.335465e-05, 3.337689e-05, 3.343307e-05, 3.346659e-05, 3.349845e-05, 
    3.356847e-05, 3.364669e-05, 3.375579e-05, 3.383398e-05, 3.388638e-05, 
    3.385421e-05, 3.388262e-05, 3.385089e-05, 3.383598e-05, 3.400123e-05, 
    3.390854e-05, 3.404747e-05, 3.403976e-05, 3.397696e-05, 3.404063e-05, 
    3.341653e-05, 3.339854e-05, 3.333629e-05, 3.338501e-05, 3.329614e-05, 
    3.334598e-05, 3.337466e-05, 3.348527e-05, 3.35095e-05, 3.353217e-05, 
    3.357677e-05, 3.363405e-05, 3.373448e-05, 3.382167e-05, 3.390109e-05, 
    3.389526e-05, 3.389732e-05, 3.391512e-05, 3.387111e-05, 3.392233e-05, 
    3.393099e-05, 3.390845e-05, 3.403874e-05, 3.400153e-05, 3.40396e-05, 
    3.401536e-05, 3.340438e-05, 3.34346e-05, 3.341828e-05, 3.344907e-05, 
    3.34274e-05, 3.352417e-05, 3.355319e-05, 3.368869e-05, 3.363295e-05, 
    3.372147e-05, 3.36419e-05, 3.365604e-05, 3.372462e-05, 3.364616e-05, 
    3.381698e-05, 3.370144e-05, 3.391581e-05, 3.380082e-05, 3.392302e-05, 
    3.390075e-05, 3.393756e-05, 3.397059e-05, 3.4012e-05, 3.408853e-05, 
    3.407079e-05, 3.413465e-05, 3.347987e-05, 3.351938e-05, 3.351579e-05, 
    3.355704e-05, 3.358756e-05, 3.365353e-05, 3.375936e-05, 3.371954e-05, 
    3.37925e-05, 3.380719e-05, 3.369626e-05, 3.37645e-05, 3.354573e-05, 
    3.358123e-05, 3.356001e-05, 3.348305e-05, 3.372888e-05, 3.360288e-05, 
    3.383529e-05, 3.376712e-05, 3.396589e-05, 3.386722e-05, 3.406105e-05, 
    3.414407e-05, 3.422157e-05, 3.431267e-05, 3.354081e-05, 3.351398e-05, 
    3.356191e-05, 3.362838e-05, 3.368968e-05, 3.37713e-05, 3.377958e-05, 
    3.379489e-05, 3.38344e-05, 3.386767e-05, 3.379985e-05, 3.387599e-05, 
    3.358969e-05, 3.373976e-05, 3.350395e-05, 3.357518e-05, 3.362441e-05, 
    3.36027e-05, 3.371496e-05, 3.374144e-05, 3.3849e-05, 3.379334e-05, 
    3.412369e-05, 3.397773e-05, 3.438157e-05, 3.426901e-05, 3.350464e-05, 
    3.354066e-05, 3.36661e-05, 3.360642e-05, 3.377668e-05, 3.381859e-05, 
    3.385255e-05, 3.389612e-05, 3.390073e-05, 3.392652e-05, 3.388427e-05, 
    3.392481e-05, 3.377147e-05, 3.384001e-05, 3.365163e-05, 3.369759e-05, 
    3.367641e-05, 3.365326e-05, 3.37247e-05, 3.380095e-05, 3.380239e-05, 
    3.382685e-05, 3.389609e-05, 3.377737e-05, 3.414286e-05, 3.391767e-05, 
    3.357994e-05, 3.364952e-05, 3.365922e-05, 3.363232e-05, 3.38144e-05, 
    3.374849e-05, 3.392587e-05, 3.387793e-05, 3.395641e-05, 3.391744e-05, 
    3.391171e-05, 3.386158e-05, 3.383041e-05, 3.375155e-05, 3.368729e-05, 
    3.36362e-05, 3.364807e-05, 3.370417e-05, 3.380557e-05, 3.390124e-05, 
    3.388031e-05, 3.395044e-05, 3.376435e-05, 3.384254e-05, 3.381239e-05, 
    3.389094e-05, 3.371852e-05, 3.386594e-05, 3.368087e-05, 3.369707e-05, 
    3.374718e-05, 3.384797e-05, 3.386996e-05, 3.389379e-05, 3.387905e-05, 
    3.38081e-05, 3.379639e-05, 3.374592e-05, 3.373207e-05, 3.369353e-05, 
    3.36617e-05, 3.369083e-05, 3.372145e-05, 3.380805e-05, 3.388612e-05, 
    3.397109e-05, 3.399179e-05, 3.409139e-05, 3.401058e-05, 3.414415e-05, 
    3.4031e-05, 3.422656e-05, 3.387419e-05, 3.402729e-05, 3.37494e-05, 
    3.377934e-05, 3.383366e-05, 3.395771e-05, 3.389057e-05, 3.396899e-05, 
    3.379592e-05, 3.37062e-05, 3.368274e-05, 3.363934e-05, 3.368373e-05, 
    3.368011e-05, 3.372259e-05, 3.370893e-05, 3.381092e-05, 3.375615e-05, 
    3.391162e-05, 3.396833e-05, 3.412803e-05, 3.422588e-05, 3.432505e-05, 
    3.436888e-05, 3.438221e-05, 3.438778e-05,
  7.917382e-10, 7.943943e-10, 7.938767e-10, 7.960262e-10, 7.9483e-10, 
    7.962423e-10, 7.922744e-10, 7.945017e-10, 7.930785e-10, 7.919743e-10, 
    8.002336e-10, 7.961221e-10, 8.044827e-10, 8.018642e-10, 8.084563e-10, 
    8.040782e-10, 8.093605e-10, 8.083215e-10, 8.114356e-10, 8.105431e-10, 
    8.145371e-10, 8.118474e-10, 8.165987e-10, 8.13892e-10, 8.143174e-10, 
    8.117595e-10, 7.969447e-10, 7.997234e-10, 7.967812e-10, 7.971772e-10, 
    7.969984e-10, 7.948563e-10, 7.937869e-10, 7.915318e-10, 7.919402e-10, 
    7.935946e-10, 7.973551e-10, 7.960692e-10, 7.993001e-10, 7.99227e-10, 
    8.028272e-10, 8.01204e-10, 8.07251e-10, 8.055313e-10, 8.105803e-10, 
    8.092945e-10, 8.105208e-10, 8.101483e-10, 8.105257e-10, 8.086396e-10, 
    8.09448e-10, 8.077867e-10, 8.01509e-10, 8.033553e-10, 7.978515e-10, 
    7.945586e-10, 7.923731e-10, 7.90826e-10, 7.910447e-10, 7.914627e-10, 
    7.936044e-10, 7.956146e-10, 7.971614e-10, 7.98197e-10, 7.992165e-10, 
    8.02316e-10, 8.039451e-10, 8.076012e-10, 8.069371e-10, 8.080687e-10, 
    8.091664e-10, 8.110154e-10, 8.107104e-10, 8.115261e-10, 8.080349e-10, 
    8.103568e-10, 8.065598e-10, 8.075777e-10, 7.995111e-10, 7.964153e-10, 
    7.951182e-10, 7.939768e-10, 7.912132e-10, 7.931226e-10, 7.923703e-10, 
    7.941566e-10, 7.95294e-10, 7.947307e-10, 7.982253e-10, 7.968645e-10, 
    8.040418e-10, 8.009501e-10, 8.090384e-10, 8.07073e-10, 8.095136e-10, 
    8.082571e-10, 8.104114e-10, 8.084725e-10, 8.118282e-10, 8.125609e-10, 
    8.120606e-10, 8.139765e-10, 8.083655e-10, 8.105225e-10, 7.947157e-10, 
    7.948077e-10, 7.952343e-10, 7.933598e-10, 7.932442e-10, 7.915214e-10, 
    7.930528e-10, 7.937063e-10, 7.953586e-10, 7.963464e-10, 7.972858e-10, 
    7.993511e-10, 8.016606e-10, 8.048848e-10, 8.071981e-10, 8.087805e-10, 
    8.07799e-10, 8.086657e-10, 8.076986e-10, 8.072575e-10, 8.122876e-10, 
    8.094566e-10, 8.137009e-10, 8.134655e-10, 8.115462e-10, 8.134919e-10, 
    7.948721e-10, 7.943433e-10, 7.925132e-10, 7.939454e-10, 7.913336e-10, 
    7.927977e-10, 7.936408e-10, 7.968967e-10, 7.976116e-10, 7.982801e-10, 
    7.995961e-10, 8.012872e-10, 8.042547e-10, 8.068337e-10, 8.092295e-10, 
    8.090517e-10, 8.091144e-10, 8.096576e-10, 8.083146e-10, 8.098779e-10, 
    8.10142e-10, 8.094542e-10, 8.13434e-10, 8.122968e-10, 8.134605e-10, 
    8.127196e-10, 7.945147e-10, 7.954036e-10, 7.949236e-10, 7.958298e-10, 
    7.951919e-10, 7.980441e-10, 7.989002e-10, 8.029012e-10, 8.012549e-10, 
    8.038702e-10, 8.015192e-10, 8.019368e-10, 8.039629e-10, 8.016451e-10, 
    8.066949e-10, 8.032779e-10, 8.096787e-10, 8.062163e-10, 8.098989e-10, 
    8.092191e-10, 8.103429e-10, 8.113514e-10, 8.126167e-10, 8.149565e-10, 
    8.144139e-10, 8.163677e-10, 7.967379e-10, 7.979029e-10, 7.977971e-10, 
    7.99014e-10, 7.999146e-10, 8.018626e-10, 8.049906e-10, 8.038133e-10, 
    8.05971e-10, 8.064053e-10, 8.031253e-10, 8.051423e-10, 7.986801e-10, 
    7.997276e-10, 7.991015e-10, 7.968317e-10, 8.040892e-10, 8.003667e-10, 
    8.07237e-10, 8.052199e-10, 8.11208e-10, 8.081956e-10, 8.141161e-10, 
    8.166554e-10, 8.190293e-10, 8.218214e-10, 7.985352e-10, 7.977439e-10, 
    7.991577e-10, 8.011197e-10, 8.029308e-10, 8.053436e-10, 8.055887e-10, 
    8.060416e-10, 8.072108e-10, 8.082096e-10, 8.06188e-10, 8.084636e-10, 
    7.99977e-10, 8.044108e-10, 7.974478e-10, 7.99549e-10, 8.010026e-10, 
    8.003617e-10, 8.03678e-10, 8.044607e-10, 8.076424e-10, 8.059958e-10, 
    8.160316e-10, 8.11569e-10, 8.239357e-10, 8.204828e-10, 7.974683e-10, 
    7.985309e-10, 8.022338e-10, 8.004715e-10, 8.055029e-10, 8.067428e-10, 
    8.077483e-10, 8.090775e-10, 8.092185e-10, 8.100056e-10, 8.087162e-10, 
    8.099534e-10, 8.053487e-10, 8.073768e-10, 8.018066e-10, 8.031644e-10, 
    8.025386e-10, 8.018547e-10, 8.039659e-10, 8.062204e-10, 8.062633e-10, 
    8.069871e-10, 8.090754e-10, 8.055231e-10, 8.166176e-10, 8.097342e-10, 
    7.996899e-10, 8.017438e-10, 8.020308e-10, 8.012363e-10, 8.066187e-10, 
    8.046692e-10, 8.099857e-10, 8.085226e-10, 8.109184e-10, 8.097283e-10, 
    8.095535e-10, 8.080238e-10, 8.070923e-10, 8.047596e-10, 8.0286e-10, 
    8.013508e-10, 8.017014e-10, 8.033589e-10, 8.063571e-10, 8.092337e-10, 
    8.085951e-10, 8.107363e-10, 8.051383e-10, 8.074513e-10, 8.06559e-10, 
    8.089195e-10, 8.037832e-10, 8.081556e-10, 8.026705e-10, 8.031493e-10, 
    8.046304e-10, 8.076118e-10, 8.082796e-10, 8.090064e-10, 8.085568e-10, 
    8.064322e-10, 8.060858e-10, 8.045932e-10, 8.041837e-10, 8.030447e-10, 
    8.021042e-10, 8.029648e-10, 8.038696e-10, 8.064309e-10, 8.087725e-10, 
    8.113666e-10, 8.119992e-10, 8.150432e-10, 8.125726e-10, 8.166569e-10, 
    8.131957e-10, 8.191812e-10, 8.084079e-10, 8.130832e-10, 8.046961e-10, 
    8.055814e-10, 8.071884e-10, 8.109577e-10, 8.089082e-10, 8.113024e-10, 
    8.060718e-10, 8.034187e-10, 8.027258e-10, 8.014436e-10, 8.027551e-10, 
    8.026482e-10, 8.039034e-10, 8.034998e-10, 8.065159e-10, 8.048956e-10, 
    8.095506e-10, 8.112821e-10, 8.161649e-10, 8.19161e-10, 8.222016e-10, 
    8.235466e-10, 8.239554e-10, 8.241267e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  0.8262706, 0.8578012, 0.8516332, 0.8773481, 0.8630461, 0.8799395, 
    0.8326243, 0.8590612, 0.8421448, 0.8290916, 0.9281192, 0.8785033, 
    0.9800585, 0.9477273, 1.029649, 0.9749979, 1.040778, 1.028065, 1.066462, 
    1.055427, 1.104865, 1.071564, 1.130647, 1.096899, 1.102167, 1.070467, 
    0.8884075, 0.9218832, 0.8864381, 0.8911781, 0.8890513, 0.8633385, 
    0.8504964, 0.8238857, 0.8286904, 0.8482506, 0.8933131, 0.8779125, 
    0.9169393, 0.9160509, 0.9595985, 0.9396477, 1.014782, 0.9932266, 
    1.055887, 1.040027, 1.055139, 1.050552, 1.055199, 1.031964, 1.041902, 
    1.021521, 0.9433708, 0.9661101, 0.899325, 0.8596799, 0.8337753, 
    0.8155981, 0.8181571, 0.8230441, 0.8483655, 0.8724767, 0.8910366, 
    0.9035381, 0.915923, 0.953165, 0.9733779, 1.019155, 1.010849, 1.024935, 
    1.038452, 1.061243, 1.057485, 1.067554, 1.024567, 1.053084, 1.006126, 
    1.018908, 0.9192813, 0.8820574, 0.8664061, 0.8528166, 0.8201267, 
    0.8426416, 0.8337337, 0.8549968, 0.868623, 0.8618732, 0.903881, 
    0.8874528, 0.9745809, 0.9365033, 1.036873, 1.012552, 1.042727, 1.027299, 
    1.05377, 1.029938, 1.071308, 1.080363, 1.074173, 1.097996, 1.028621, 
    1.055137, 0.8616835, 0.8627826, 0.8679133, 0.8454557, 0.8440912, 
    0.8237532, 0.8418411, 0.8495937, 0.8694172, 0.8812286, 0.8925179, 
    0.9175386, 0.9451986, 0.9851022, 1.014123, 1.03372, 1.021692, 1.032309, 
    1.020442, 1.014894, 1.076967, 1.041994, 1.094564, 1.091642, 1.067792, 
    1.091971, 0.8635551, 0.8572351, 0.83544, 0.8524762, 0.8215517, 0.8387983, 
    0.8487839, 0.8877906, 0.8964612, 0.9045248, 0.9205369, 0.9406648, 
    0.9772673, 1.009516, 1.039241, 1.037055, 1.037825, 1.044493, 1.027993, 
    1.047209, 1.050441, 1.041992, 1.09125, 1.077128, 1.09158, 1.082381, 
    0.8592878, 0.8699447, 0.864179, 0.8750332, 0.867379, 0.9016173, 
    0.9119847, 0.9604535, 0.9402559, 0.9724813, 0.9435121, 0.9486201, 
    0.9735306, 0.9450704, 1.007726, 0.9650831, 1.044752, 1.001666, 1.047469, 
    1.039112, 1.052959, 1.065397, 1.081093, 1.110161, 1.10342, 1.127797, 
    0.8859342, 0.899938, 0.8987052, 0.913447, 0.9244075, 0.9477379, 
    0.9864512, 0.9718289, 0.9987342, 1.004164, 0.9633149, 0.9883232, 
    0.9093609, 0.9220641, 0.9144955, 0.8870336, 0.9751865, 0.9298811, 
    1.014605, 0.9893239, 1.063621, 1.026476, 1.09971, 1.131288, 1.1611, 
    1.195929, 0.9076212, 0.898064, 0.9152073, 0.938555, 0.9608834, 0.9908593, 
    0.9939462, 0.9996017, 1.014303, 1.026712, 1.001388, 1.02983, 0.9250122, 
    0.9792054, 0.8944576, 0.9198753, 0.9371457, 0.9298727, 0.9701636, 
    0.9798784, 1.019687, 0.9990464, 1.123481, 1.068022, 1.222411, 1.179211, 
    0.8947333, 0.9075899, 0.9522578, 0.9312239, 0.9928737, 1.008394, 1.02107, 
    1.037335, 1.039098, 1.048772, 1.032931, 1.048147, 0.9909233, 1.016378, 
    0.9470624, 0.9637719, 0.9560726, 0.9476511, 0.973731, 1.001785, 1.002393, 
    1.011444, 1.037069, 0.9931286, 1.130656, 1.045211, 0.9216895, 0.9461933, 
    0.9497936, 0.9400603, 1.006835, 0.9824532, 1.048537, 1.030554, 1.060062, 
    1.045371, 1.043214, 1.024437, 1.012794, 0.9835655, 0.9600021, 0.9414703, 
    0.9457675, 0.9661667, 1.00351, 1.039255, 1.031393, 1.057812, 0.9883159, 
    1.017285, 1.006055, 1.035415, 0.97144, 1.025821, 0.9577007, 0.9636099, 
    0.9819713, 1.019255, 1.027571, 1.03646, 1.030974, 1.004466, 1.000146, 
    0.9815251, 0.9764018, 0.9623227, 0.9507205, 0.9613174, 0.9724913, 
    1.00448, 1.033583, 1.065573, 1.073439, 1.111118, 1.080419, 1.131134, 
    1.08798, 1.162792, 1.029009, 1.086728, 0.9828117, 0.9938608, 1.013941, 
    1.060447, 1.035277, 1.064731, 0.9999773, 0.9668703, 0.9583764, 0.9425918, 
    0.9587384, 0.9574215, 0.9729594, 0.9679568, 1.005548, 0.9852951, 
    1.043158, 1.064499, 1.125237, 1.162665, 1.200788, 1.217586, 1.222693, 
    1.224826,
  0.8832567, 0.8685132, 0.8713382, 0.859753, 0.8661355, 0.8586136, 0.8802259, 
    0.8679388, 0.8757402, 0.8819085, 0.8383449, 0.8592446, 0.7816319, 
    0.7895164, 0.7707522, 0.7828236, 0.7685093, 0.7710784, 0.7636082, 
    0.7656676, 0.7569872, 0.7626798, 0.7530208, 0.7582913, 0.757425, 
    0.7628779, 0.8549269, 0.8408688, 0.8557796, 0.8537307, 0.8546486, 
    0.8660024, 0.8718591, 0.884405, 0.8821, 0.8728986, 0.8528135, 0.8595064, 
    0.8428994, 0.8432647, 0.7865486, 0.7915862, 0.773863, 0.7786027, 
    0.7655804, 0.7686595, 0.765722, 0.7665998, 0.7657106, 0.7702807, 
    0.7682874, 0.7724374, 0.7906274, 0.7849565, 0.850251, 0.8676548, 
    0.8796793, 0.8884217, 0.8871755, 0.8848091, 0.8728453, 0.8619109, 
    0.8537936, 0.8484724, 0.8433173, 0.7881437, 0.7832091, 0.7729341, 
    0.7747076, 0.7717246, 0.7689731, 0.764573, 0.765278, 0.7634078, 0.771802, 
    0.7661131, 0.7757338, 0.7729871, 0.8419301, 0.8576879, 0.8646181, 
    0.8707936, 0.8862196, 0.8755069, 0.8796985, 0.8697955, 0.863629, 
    0.8666664, 0.8483281, 0.8553404, 0.7829232, 0.7924016, 0.7692891, 
    0.7743406, 0.7681249, 0.7712366, 0.7659824, 0.7706944, 0.7627257, 
    0.7611132, 0.7622103, 0.7581103, 0.7709644, 0.765722, 0.8667518, 
    0.8662546, 0.8639472, 0.8741951, 0.8748308, 0.8844683, 0.8758823, 
    0.8722782, 0.8632748, 0.8580503, 0.8531563, 0.8426524, 0.7901592, 
    0.7804595, 0.7740037, 0.7699247, 0.7724019, 0.7702109, 0.7726641, 
    0.7738394, 0.7617122, 0.7682691, 0.7586809, 0.7591721, 0.763364, 
    0.7591165, 0.8659059, 0.8687732, 0.8788918, 0.8709516, 0.8855307, 
    0.8773083, 0.8726511, 0.855192, 0.8514701, 0.8480566, 0.8414258, 
    0.7913235, 0.7822885, 0.774995, 0.768816, 0.7692528, 0.7690988, 
    0.7677775, 0.7710935, 0.767247, 0.7666207, 0.7682699, 0.7592382, 
    0.7616843, 0.7591826, 0.7607612, 0.8678389, 0.8630387, 0.8656248, 
    0.8607767, 0.8641855, 0.8492793, 0.8449404, 0.7863368, 0.7914287, 
    0.7834235, 0.7905915, 0.7892902, 0.7831714, 0.7901933, 0.7753831, 
    0.7852044, 0.7677266, 0.7767118, 0.7671964, 0.7688417, 0.7661378, 
    0.7638035, 0.7609859, 0.756142, 0.7572222, 0.753441, 0.855999, 0.8499909, 
    0.8505156, 0.8443382, 0.8398511, 0.7895144, 0.7801488, 0.7835804, 
    0.7773657, 0.7761635, 0.7856376, 0.7797184, 0.8460327, 0.8408003, 
    0.8439046, 0.8555209, 0.7827799, 0.8376423, 0.7739007, 0.7794899, 
    0.7641312, 0.7714053, 0.7578275, 0.7529262, 0.74883, 0.7446977, 
    0.8467593, 0.8507881, 0.8436121, 0.7918679, 0.7862325, 0.7791396, 
    0.7784401, 0.7771721, 0.7739657, 0.7713577, 0.7767748, 0.7707166, 
    0.8395999, 0.7818326, 0.8523245, 0.8416925, 0.7922344, 0.8376477, 
    0.7839796, 0.7816759, 0.7728222, 0.7772961, 0.7540839, 0.7633212, 
    0.7420376, 0.7465922, 0.8522078, 0.8467733, 0.7883733, 0.8371067, 
    0.7786826, 0.7752388, 0.7725323, 0.7691962, 0.7688444, 0.7669433, 
    0.7700847, 0.7670648, 0.779125, 0.7735231, 0.7896861, 0.7855255, 
    0.7874219, 0.7895367, 0.783127, 0.7766868, 0.7765538, 0.7745785, 
    0.7692453, 0.778625, 0.7530167, 0.7676329, 0.8409563, 0.7899051, 
    0.788994, 0.7914799, 0.7755784, 0.7810744, 0.766989, 0.7705687, 0.764794, 
    0.7676055, 0.7680289, 0.7718291, 0.7742887, 0.7808157, 0.7864491, 
    0.7911164, 0.7900156, 0.7849429, 0.7763062, 0.7688127, 0.7703965, 
    0.7652165, 0.7797208, 0.7733299, 0.7757481, 0.7695822, 0.7836731, 
    0.771538, 0.787018, 0.7855656, 0.7811866, 0.7729123, 0.7711805, 
    0.7693716, 0.7704828, 0.7760964, 0.777051, 0.781291, 0.7824931, 
    0.7858803, 0.7887609, 0.7861263, 0.7834215, 0.776094, 0.7699518, 
    0.7637709, 0.7623423, 0.7559892, 0.7611021, 0.7529466, 0.7597899, 
    0.7486107, 0.7708824, 0.7600067, 0.7809915, 0.7784595, 0.7740417, 
    0.7647203, 0.7696101, 0.7639252, 0.7770886, 0.7847717, 0.7868508, 
    0.7908277, 0.7867613, 0.7870871, 0.7833108, 0.7845109, 0.7758598, 
    0.780416, 0.7680395, 0.7639683, 0.7538216, 0.7486283, 0.7441791, 
    0.7424913, 0.7420118, 0.7418161,
  1.192281, 1.192544, 1.192521, 1.192529, 1.192554, 1.192517, 1.192362, 
    1.192547, 1.192458, 1.192319, 1.191841, 1.192524, 1.229236, 1.235678, 
    1.219249, 1.230246, 1.216988, 1.219573, 1.211734, 1.213998, 1.20377, 
    1.210684, 1.198349, 1.205434, 1.204335, 1.21091, 1.19246, 1.191976, 
    1.192475, 1.192435, 1.192454, 1.192554, 1.192515, 1.192246, 1.192314, 
    1.192502, 1.192414, 1.192527, 1.192075, 1.192092, 1.233319, 1.237281, 
    1.222261, 1.226601, 1.213904, 1.217142, 1.214057, 1.214996, 1.214044, 
    1.218781, 1.21676, 1.220899, 1.236543, 1.232022, 1.192347, 1.192548, 
    1.192376, 1.192111, 1.192156, 1.192234, 1.192503, 1.192546, 1.192437, 
    1.192293, 1.192094, 1.234595, 1.230571, 1.221376, 1.223055, 1.220206, 
    1.217463, 1.212805, 1.213577, 1.211509, 1.220282, 1.214476, 1.224008, 
    1.221427, 1.192029, 1.192505, 1.192554, 1.192526, 1.192188, 1.192462, 
    1.192375, 1.192536, 1.192553, 1.192553, 1.192288, 1.192468, 1.230331, 
    1.237903, 1.217784, 1.222711, 1.216592, 1.219729, 1.214337, 1.219193, 
    1.210736, 1.208866, 1.210145, 1.205207, 1.21946, 1.214056, 1.192552, 
    1.192554, 1.192554, 1.192483, 1.192473, 1.192244, 1.192455, 1.19251, 
    1.192552, 1.19251, 1.192423, 1.192064, 1.236179, 1.228228, 1.222394, 
    1.218426, 1.220865, 1.218712, 1.221117, 1.222239, 1.209568, 1.216741, 
    1.205922, 1.20653, 1.211459, 1.206461, 1.192554, 1.192543, 1.192394, 
    1.192525, 1.192211, 1.192428, 1.192505, 1.192465, 1.192381, 1.192279, 
    1.192005, 1.23708, 1.229795, 1.223323, 1.217303, 1.217748, 1.217591, 
    1.216232, 1.219588, 1.215678, 1.215017, 1.216742, 1.206611, 1.209536, 
    1.206542, 1.20845, 1.192548, 1.192551, 1.192555, 1.192538, 1.192554, 
    1.192318, 1.192163, 1.233147, 1.23716, 1.230751, 1.236515, 1.235501, 
    1.230538, 1.236207, 1.223683, 1.232225, 1.216179, 1.224901, 1.215625, 
    1.217329, 1.214503, 1.211952, 1.208716, 1.202664, 1.204075, 1.198953, 
    1.192479, 1.19234, 1.192355, 1.192138, 1.191925, 1.235677, 1.227958, 
    1.230883, 1.225495, 1.224402, 1.23258, 1.227583, 1.192206, 1.191974, 
    1.192119, 1.192471, 1.23021, 1.191802, 1.222297, 1.227383, 1.212317, 
    1.219894, 1.204849, 1.198211, 1.191852, 1.184271, 1.192233, 1.192363, 
    1.192107, 1.237496, 1.233064, 1.227075, 1.226456, 1.22532, 1.222358, 
    1.219848, 1.224959, 1.219215, 1.191911, 1.229408, 1.192403, 1.192018, 
    1.237776, 1.191802, 1.231215, 1.229275, 1.221269, 1.225432, 1.199861, 
    1.21141, 1.178395, 1.18793, 1.1924, 1.192234, 1.234778, 1.19177, 
    1.226671, 1.22355, 1.220991, 1.21769, 1.217332, 1.215358, 1.218586, 
    1.215487, 1.227062, 1.221939, 1.235812, 1.232489, 1.234022, 1.235695, 
    1.230503, 1.224879, 1.224759, 1.222934, 1.217736, 1.22662, 1.19834, 
    1.216079, 1.191982, 1.235981, 1.235269, 1.2372, 1.223864, 1.228759, 
    1.215407, 1.219069, 1.213048, 1.216053, 1.216493, 1.220309, 1.222663, 
    1.228536, 1.233239, 1.236921, 1.236068, 1.232011, 1.224532, 1.217299, 
    1.218897, 1.21351, 1.227585, 1.221755, 1.22402, 1.218081, 1.23096, 
    1.220021, 1.233698, 1.232522, 1.228855, 1.221355, 1.219674, 1.217867, 
    1.218983, 1.22434, 1.22521, 1.228945, 1.229969, 1.232778, 1.235085, 
    1.232978, 1.230749, 1.224338, 1.218452, 1.211916, 1.210297, 1.20246, 
    1.208852, 1.198239, 1.20728, 1.191481, 1.219378, 1.207545, 1.228688, 
    1.226473, 1.222429, 1.212966, 1.218109, 1.212087, 1.225244, 1.23187, 
    1.233563, 1.236698, 1.233491, 1.233753, 1.230657, 1.231655, 1.224123, 
    1.228191, 1.216504, 1.212136, 1.199493, 1.191512, 1.183204, 1.179475, 
    1.178333, 1.177854,
  0.5002306, 0.4900042, 0.49199, 0.4837597, 0.488323, 0.4829374, 0.4981552, 
    0.4895985, 0.4950586, 0.4993093, 0.4678519, 0.4833932, 0.4518529, 
    0.4616959, 0.4370518, 0.4533813, 0.4337747, 0.4375222, 0.4262669, 
    0.4294848, 0.4151588, 0.4247836, 0.4077797, 0.4174533, 0.415936, 
    0.4251018, 0.4802597, 0.4697816, 0.4808815, 0.4793847, 0.4800565, 
    0.4882283, 0.4923539, 0.5010141, 0.4994404, 0.4930809, 0.4787119, 
    0.4835826, 0.4713252, 0.4716014, 0.4580641, 0.4641818, 0.4414575, 
    0.4478934, 0.4293504, 0.4339978, 0.4295683, 0.4309105, 0.4295508, 
    0.4363712, 0.4334461, 0.4394585, 0.4630347, 0.4560805, 0.4768235, 
    0.4893971, 0.4977793, 0.5037391, 0.502896, 0.501289, 0.4930437, 
    0.4853113, 0.4794314, 0.4755046, 0.4716412, 0.4600243, 0.4538731, 
    0.4401579, 0.4426276, 0.4384462, 0.4344608, 0.4277862, 0.4288833, 
    0.4259481, 0.4385571, 0.4301678, 0.4440355, 0.4402331, 0.4705881, 
    0.482268, 0.4872436, 0.4916081, 0.5022478, 0.4948964, 0.4977924, 
    0.4909076, 0.4865399, 0.4886995, 0.4753973, 0.4805616, 0.453509, 
    0.4651503, 0.4349252, 0.4421206, 0.4332045, 0.4377495, 0.4299679, 
    0.4369699, 0.4248571, 0.4222293, 0.4240246, 0.4171391, 0.4373587, 
    0.4295679, 0.4887598, 0.4884075, 0.486767, 0.4939846, 0.4944269, 
    0.5010571, 0.4951572, 0.4926477, 0.4862872, 0.4825305, 0.478964, 
    0.471138, 0.4624713, 0.4503334, 0.4416534, 0.4358545, 0.4394086, 
    0.4362705, 0.4397787, 0.4414252, 0.4232133, 0.4334186, 0.4181279, 
    0.4189708, 0.4258782, 0.4188758, 0.4881602, 0.490188, 0.4972372, 
    0.4917193, 0.5017799, 0.4961443, 0.4929079, 0.4804528, 0.4777241, 
    0.475195, 0.4702078, 0.4638683, 0.452698, 0.443023, 0.4342293, 0.4348724, 
    0.434646, 0.4326859, 0.437544, 0.4318895, 0.4309417, 0.4334202, 
    0.4190837, 0.4231684, 0.4189887, 0.4216472, 0.4895288, 0.4861183, 
    0.4879607, 0.484497, 0.4869365, 0.4761032, 0.4728631, 0.4578009, 
    0.4639937, 0.4541462, 0.4629919, 0.461422, 0.4538241, 0.4625133, 
    0.4435546, 0.4563898, 0.4326098, 0.4453607, 0.4318133, 0.4342673, 
    0.4302063, 0.426576, 0.4220195, 0.4136409, 0.4155777, 0.4085945, 
    0.4810415, 0.4766308, 0.4770196, 0.4724111, 0.4690076, 0.4616939, 
    0.4499284, 0.4543461, 0.4462433, 0.44462, 0.4569329, 0.4493644, 
    0.4736834, 0.469731, 0.472084, 0.4806929, 0.4533264, 0.4673133, 
    0.4415101, 0.4490649, 0.4270931, 0.43799, 0.4166447, 0.407594, 0.3991242, 
    0.3892808, 0.4742273, 0.4772209, 0.4718637, 0.4645162, 0.4576724, 
    0.4486032, 0.4476776, 0.4459831, 0.4416008, 0.4379228, 0.4454469, 
    0.4370019, 0.4688138, 0.4521122, 0.4783528, 0.4704094, 0.4649521, 
    0.4673182, 0.4548517, 0.4519111, 0.4400007, 0.44615, 0.4098227, 
    0.4258091, 0.3818324, 0.3939979, 0.4782674, 0.4742379, 0.4603064, 
    0.4669015, 0.4479994, 0.443358, 0.4395928, 0.4347886, 0.4342712, 
    0.4314309, 0.4360872, 0.4316149, 0.4485839, 0.4409839, 0.4619018, 
    0.4567927, 0.4591419, 0.4617209, 0.4537701, 0.4453281, 0.4451492, 
    0.4424491, 0.434857, 0.4479229, 0.4077681, 0.4324659, 0.4698507, 
    0.4621646, 0.4610628, 0.4640554, 0.4438228, 0.4511333, 0.4315002, 
    0.4367884, 0.4281315, 0.4324284, 0.4330614, 0.4385958, 0.4420488, 
    0.4507973, 0.4579409, 0.4636213, 0.4622994, 0.4560637, 0.444813, 
    0.4342238, 0.4365386, 0.4287881, 0.4493683, 0.4407133, 0.444054, 
    0.4353546, 0.4544633, 0.438177, 0.4586447, 0.456843, 0.4512786, 
    0.4401268, 0.437669, 0.435046, 0.4366644, 0.4445283, 0.44582, 0.451414, 
    0.4529604, 0.4572352, 0.4607797, 0.4575408, 0.4541438, 0.4445255, 
    0.4358934, 0.4265242, 0.4242387, 0.4133615, 0.4222096, 0.4076313, 
    0.4200155, 0.3986368, 0.4372387, 0.4203833, 0.4510261, 0.4477035, 
    0.4417051, 0.4280151, 0.4353954, 0.4267674, 0.4458707, 0.4558483, 
    0.4584382, 0.4632753, 0.4583277, 0.4587298, 0.454004, 0.4555217, 
    0.4442069, 0.4502777, 0.433077, 0.4268357, 0.4093246, 0.3986777, 
    0.3879162, 0.3831898, 0.3817545, 0.3811548,
  0.04899357, 0.04712923, 0.0474883, 0.04600939, 0.04682634, 0.04586296, 
    0.04861216, 0.04705605, 0.04804596, 0.04882406, 0.0432199, 0.04594409, 
    0.04049848, 0.04215674, 0.03806951, 0.04075371, 0.03754215, 0.03814552, 
    0.03634823, 0.03685753, 0.03461802, 0.03611469, 0.03349244, 0.03497186, 
    0.03473766, 0.03616472, 0.04538786, 0.04355346, 0.04549796, 0.04523317, 
    0.04535191, 0.04680932, 0.04755424, 0.04913798, 0.04884817, 0.04768615, 
    0.04511441, 0.04597783, 0.04382122, 0.04386923, 0.04154088, 0.042581, 
    0.03878443, 0.03984112, 0.03683619, 0.03757794, 0.0368708, 0.03708434, 
    0.03686802, 0.03795968, 0.03748948, 0.03845919, 0.04238496, 0.04120649, 
    0.04478194, 0.04701974, 0.04854323, 0.04964194, 0.04948571, 0.04918868, 
    0.0476794, 0.04628632, 0.0452414, 0.04455051, 0.04387613, 0.04187271, 
    0.04083603, 0.03857284, 0.03897546, 0.03829505, 0.03765225, 0.03658824, 
    0.03676207, 0.03629798, 0.03831301, 0.0369661, 0.03920594, 0.03858506, 
    0.04369326, 0.04574395, 0.04663243, 0.04741913, 0.04936578, 0.04801639, 
    0.04854564, 0.0472924, 0.04650624, 0.04689409, 0.04453171, 0.04544129, 
    0.04077508, 0.04274688, 0.03772687, 0.03889262, 0.03745079, 0.03818227, 
    0.03693431, 0.03805629, 0.03612626, 0.03571434, 0.03599549, 0.03492332, 
    0.03811909, 0.03687074, 0.04690496, 0.04684155, 0.04654693, 0.0478504, 
    0.04793088, 0.0491459, 0.04806394, 0.04760753, 0.04646096, 0.0457906, 
    0.04515888, 0.0437887, 0.04228884, 0.04024556, 0.03881637, 0.0378764, 
    0.0384511, 0.03794343, 0.0385112, 0.03877917, 0.03586829, 0.03748509, 
    0.03507626, 0.03520691, 0.03628697, 0.03519218, 0.04679707, 0.04716241, 
    0.04844395, 0.04743927, 0.04927934, 0.04824408, 0.04765475, 0.04542203, 
    0.04494033, 0.04449627, 0.04362729, 0.04252737, 0.0406395, 0.03904011, 
    0.03761509, 0.03771838, 0.03768199, 0.03736778, 0.03814904, 0.0372405, 
    0.03708932, 0.03748535, 0.03522443, 0.03586126, 0.03520969, 0.03562342, 
    0.04704348, 0.04643071, 0.04676121, 0.04614087, 0.04657733, 0.04465546, 
    0.04408885, 0.04149643, 0.04254882, 0.04088176, 0.04237765, 0.04211013, 
    0.04082782, 0.042296, 0.03912714, 0.04125855, 0.03735561, 0.03942354, 
    0.03722833, 0.03762118, 0.03697222, 0.036397, 0.03568155, 0.03438493, 
    0.03468248, 0.03361579, 0.0455263, 0.0447481, 0.0448164, 0.0440101, 
    0.04341951, 0.04215639, 0.04017828, 0.04091526, 0.0395688, 0.03930184, 
    0.04135002, 0.04008468, 0.04423194, 0.04354468, 0.04395317, 0.04546455, 
    0.04074454, 0.04312705, 0.038793, 0.04003502, 0.03647865, 0.03822119, 
    0.03484695, 0.03346437, 0.03219633, 0.0307539, 0.04432696, 0.04485179, 
    0.04391484, 0.04263823, 0.04147475, 0.03995854, 0.03980545, 0.03952594, 
    0.0388078, 0.03821031, 0.03943771, 0.03806145, 0.043386, 0.04054173, 
    0.04505109, 0.04366225, 0.0427129, 0.04312788, 0.04100005, 0.04050818, 
    0.03854728, 0.03955342, 0.03380217, 0.03627608, 0.02968469, 0.03144095, 
    0.04503603, 0.04432882, 0.04192057, 0.04305611, 0.03985863, 0.03909494, 
    0.03848102, 0.03770492, 0.03762181, 0.03716731, 0.03791389, 0.03719667, 
    0.03995535, 0.03870725, 0.04219179, 0.04132639, 0.04172317, 0.04216101, 
    0.04081878, 0.03941817, 0.03938876, 0.03894628, 0.0377159, 0.03984599, 
    0.03349069, 0.03733261, 0.04356542, 0.04223656, 0.04204905, 0.04255937, 
    0.03917108, 0.04037859, 0.03717837, 0.03802698, 0.03664291, 0.03732662, 
    0.03742787, 0.03831928, 0.0388809, 0.04032269, 0.04152007, 0.04248514, 
    0.04225953, 0.04120367, 0.03933353, 0.0376142, 0.03798668, 0.03674696, 
    0.04008533, 0.03866319, 0.03920899, 0.03779593, 0.04093491, 0.03825146, 
    0.04163902, 0.04133487, 0.0404028, 0.03856777, 0.03816926, 0.0377463, 
    0.03800697, 0.03928679, 0.03949909, 0.04042534, 0.04068334, 0.04140099, 
    0.04200094, 0.04145253, 0.04088137, 0.03928632, 0.03788266, 0.03638883, 
    0.0360291, 0.03434212, 0.03571125, 0.03347, 0.0353692, 0.03212411, 
    0.0380997, 0.03542642, 0.04036076, 0.03980972, 0.03882482, 0.03662447, 
    0.0378025, 0.03642721, 0.03950743, 0.04116744, 0.0416041, 0.04242604, 
    0.04158543, 0.04165341, 0.04085794, 0.04111254, 0.03923405, 0.04023629, 
    0.03743037, 0.036438, 0.03372652, 0.03213017, 0.03055659, 0.02987812, 
    0.02967361, 0.02958838,
  0.00131427, 0.001238153, 0.001252693, 0.001193181, 0.001225934, 
    0.001187343, 0.001298572, 0.001235197, 0.001275388, 0.001307286, 
    0.001083652, 0.001190576, 0.0009803121, 0.001042861, 0.0008911084, 
    0.0009898534, 0.0008721279, 0.0008938554, 0.0008296767, 0.0008476969, 
    0.0007694578, 0.0008214579, 0.0007316489, 0.0007816464, 0.0007735715, 
    0.0008232164, 0.001168467, 0.001096559, 0.001172832, 0.001162343, 
    0.001167042, 0.001225248, 0.001255369, 0.001320231, 0.001308279, 
    0.001260729, 0.001157649, 0.001191922, 0.001106958, 0.001108826, 
    0.001019477, 0.001059074, 0.0009170615, 0.0009558845, 0.000846939, 
    0.0008734115, 0.0008481679, 0.0008557644, 0.0008480692, 0.0008871437, 
    0.00087024, 0.000905223, 0.001051572, 0.001006857, 0.001144543, 
    0.001233731, 0.001295742, 0.001341102, 0.00133462, 0.001322325, 
    0.001260454, 0.00120425, 0.001162669, 0.00113545, 0.001109094, 
    0.001032054, 0.000992937, 0.0009093537, 0.0009240392, 0.0008992681, 
    0.0008760789, 0.0008381523, 0.000844309, 0.0008279059, 0.0008999192, 
    0.0008515554, 0.0009324818, 0.0009097983, 0.001101984, 0.001182604, 
    0.001218132, 0.001249887, 0.001329652, 0.001274181, 0.001295841, 
    0.001244753, 0.001213064, 0.001228663, 0.001134712, 0.001170584, 
    0.0009906536, 0.001065437, 0.0008787603, 0.000921011, 0.0008688537, 
    0.0008951848, 0.0008504249, 0.0008906306, 0.0008218644, 0.0008074343, 
    0.0008172741, 0.0007799702, 0.0008928999, 0.000848166, 0.001229101, 
    0.001226546, 0.001214698, 0.001267413, 0.001270693, 0.001320558, 
    0.001276122, 0.001257534, 0.001211248, 0.001184461, 0.001159406, 
    0.001105693, 0.0010479, 0.0009708887, 0.0009182268, 0.0008841418, 
    0.0009049291, 0.0008865579, 0.0009071126, 0.0009168694, 0.0008128173, 
    0.0008700824, 0.0007852548, 0.0007897792, 0.000827518, 0.0007892685, 
    0.001224755, 0.001239494, 0.00129167, 0.001250704, 0.001326074, 
    0.001283485, 0.001259452, 0.001169821, 0.00115078, 0.001133322, 
    0.001099423, 0.00105702, 0.0009855799, 0.0009264046, 0.0008747447, 
    0.0008784551, 0.0008771472, 0.000865883, 0.0008939829, 0.0008613341, 
    0.0008559416, 0.0008700917, 0.0007903865, 0.0008125713, 0.0007898756, 
    0.000804261, 0.001234689, 0.001210035, 0.001223311, 0.001198432, 
    0.001215919, 0.00113957, 0.001117385, 0.001017796, 0.001057842, 
    0.0009946519, 0.001051292, 0.001041085, 0.0009926296, 0.001048173, 
    0.0009295924, 0.001008818, 0.0008654474, 0.0009404769, 0.0008608997, 
    0.0008749633, 0.0008517732, 0.0008313966, 0.0008062895, 0.0007614648, 
    0.0007716733, 0.0007352938, 0.001173956, 0.001143212, 0.001145899, 
    0.001114313, 0.001091369, 0.001042848, 0.0009683874, 0.0009959085, 
    0.0009458269, 0.0009360024, 0.001012267, 0.0009649109, 0.001122974, 
    0.001096219, 0.001112094, 0.001171506, 0.0009895097, 0.001080068, 
    0.000917374, 0.000963068, 0.0008342788, 0.0008965931, 0.0007773361, 
    0.0007306987, 0.0006882285, 0.0006410086, 0.00112669, 0.001147292, 
    0.001110601, 0.001061268, 0.001016977, 0.0009602325, 0.0009545651, 
    0.0009442474, 0.0009179139, 0.0008961994, 0.0009409984, 0.0008908173, 
    0.001090073, 0.0009819268, 0.001155149, 0.00110078, 0.001064132, 
    0.0010801, 0.0009990917, 0.0009806742, 0.000908424, 0.00094526, 
    0.000741607, 0.0008271347, 0.0006067723, 0.0006633534, 0.001154555, 
    0.001126763, 0.001033872, 0.001077333, 0.0009565327, 0.0009284126, 
    0.0009060156, 0.0008779712, 0.0008749858, 0.0008587221, 0.0008854929, 
    0.0008597694, 0.0009601143, 0.0009142474, 0.001044197, 0.001011376, 
    0.00102638, 0.001043023, 0.0009922907, 0.0009402794, 0.0009391975, 
    0.000922972, 0.000878366, 0.0009560649, 0.0007315895, 0.000864625, 
    0.001097023, 0.001045905, 0.001038759, 0.001058246, 0.0009312034, 
    0.0009758415, 0.0008591166, 0.0008895724, 0.000840087, 0.0008644107, 
    0.0008680332, 0.0009001466, 0.0009205827, 0.0009737593, 0.00101869, 
    0.001055403, 0.001046781, 0.00100675, 0.0009371669, 0.0008747129, 
    0.0008881178, 0.0008437734, 0.0009649351, 0.0009126421, 0.0009325935, 
    0.0008812441, 0.0009966461, 0.000897689, 0.001023191, 0.001011695, 
    0.0009767435, 0.0009091693, 0.000894714, 0.0008794587, 0.0008888501, 
    0.0009354498, 0.000943258, 0.0009775839, 0.0009872197, 0.001014191, 
    0.001036928, 0.001016137, 0.000994637, 0.0009354325, 0.0008843673, 
    0.0008311083, 0.0008184531, 0.00076, 0.0008073265, 0.0007308893, 
    0.0007954112, 0.0006858364, 0.000892199, 0.0007974001, 0.000975177, 
    0.0009547229, 0.0009185351, 0.0008394341, 0.0008814806, 0.0008324627, 
    0.0009435654, 0.001005386, 0.001021869, 0.001053143, 0.001021162, 
    0.001023736, 0.0009937588, 0.00100332, 0.0009335132, 0.0009705442, 
    0.0008681227, 0.0008328431, 0.0007390421, 0.000686037, 0.000634641, 
    0.0006129171, 0.000606421, 0.0006037209,
  8.639036e-06, 7.877293e-06, 8.021053e-06, 7.437973e-06, 7.757118e-06, 
    7.38154e-06, 8.480111e-06, 7.848163e-06, 8.247116e-06, 8.56821e-06, 
    6.403206e-06, 7.41278e-06, 5.47571e-06, 6.031217e-06, 4.716436e-06, 
    5.559251e-06, 4.560141e-06, 4.739214e-06, 4.217587e-06, 4.361798e-06, 
    3.748965e-06, 4.15241e-06, 3.143209e-06, 3.842126e-06, 3.78031e-06, 
    4.166324e-06, 7.200055e-06, 6.522464e-06, 7.241892e-06, 7.141493e-06, 
    7.18642e-06, 7.750391e-06, 8.047609e-06, 8.699624e-06, 8.578267e-06, 
    8.10087e-06, 7.096713e-06, 7.425792e-06, 6.619076e-06, 6.636481e-06, 
    5.821392e-06, 6.178177e-06, 4.933193e-06, 5.263839e-06, 4.355697e-06, 
    4.570652e-06, 4.365591e-06, 4.426938e-06, 4.364797e-06, 4.683632e-06, 
    4.5447e-06, 4.833887e-06, 6.110024e-06, 5.709207e-06, 6.97217e-06, 
    7.833734e-06, 8.451562e-06, 8.91284e-06, 8.846449e-06, 8.720951e-06, 
    8.09814e-06, 7.545339e-06, 7.144605e-06, 6.886191e-06, 6.638986e-06, 
    5.93393e-06, 5.586345e-06, 4.868455e-06, 4.99206e-06, 4.78421e-06, 
    4.592519e-06, 4.285192e-06, 4.33455e-06, 4.203512e-06, 4.789632e-06, 
    4.392909e-06, 5.063618e-06, 4.872181e-06, 6.572807e-06, 7.335846e-06, 
    7.680704e-06, 7.993249e-06, 8.795663e-06, 8.235046e-06, 8.452559e-06, 
    7.942444e-06, 7.631198e-06, 7.783909e-06, 6.879232e-06, 7.220342e-06, 
    5.566279e-06, 6.236173e-06, 4.61454e-06, 4.966483e-06, 4.533374e-06, 
    4.75025e-06, 4.383786e-06, 4.712479e-06, 4.155625e-06, 4.04208e-06, 
    4.119378e-06, 3.829262e-06, 4.731286e-06, 4.365576e-06, 7.78821e-06, 
    7.763128e-06, 7.647144e-06, 8.167453e-06, 8.200187e-06, 8.702957e-06, 
    8.254461e-06, 8.069102e-06, 7.613479e-06, 7.35374e-06, 7.113463e-06, 
    6.6073e-06, 6.076766e-06, 5.393632e-06, 4.943007e-06, 4.658849e-06, 
    4.831432e-06, 4.678792e-06, 4.84969e-06, 4.931576e-06, 4.084299e-06, 
    4.543412e-06, 3.869873e-06, 3.904771e-06, 4.200431e-06, 3.900826e-06, 
    7.745557e-06, 7.890515e-06, 8.410528e-06, 8.00134e-06, 8.759151e-06, 
    8.328248e-06, 8.088173e-06, 7.213024e-06, 7.031354e-06, 6.866123e-06, 
    6.549024e-06, 6.159492e-06, 5.521781e-06, 5.012073e-06, 4.581576e-06, 
    4.612031e-06, 4.601288e-06, 4.509136e-06, 4.740272e-06, 4.472115e-06, 
    4.428373e-06, 4.543489e-06, 3.909465e-06, 4.082366e-06, 3.905516e-06, 
    4.017268e-06, 7.843168e-06, 7.601654e-06, 7.731407e-06, 7.488843e-06, 
    7.659069e-06, 6.925111e-06, 6.716425e-06, 5.80641e-06, 6.166963e-06, 
    5.601431e-06, 6.107492e-06, 6.01519e-06, 5.583641e-06, 6.079239e-06, 
    5.039086e-06, 5.726592e-06, 4.505587e-06, 5.131712e-06, 4.468586e-06, 
    4.583369e-06, 4.394667e-06, 4.231273e-06, 4.033122e-06, 3.68835e-06, 
    3.765834e-06, 3.492572e-06, 7.252682e-06, 6.959562e-06, 6.985024e-06, 
    6.687697e-06, 6.474428e-06, 6.031099e-06, 5.371918e-06, 5.612495e-06, 
    5.177457e-06, 5.093563e-06, 5.757209e-06, 5.341789e-06, 6.768795e-06, 
    6.519311e-06, 6.666973e-06, 7.22918e-06, 5.556235e-06, 6.370226e-06, 
    4.935825e-06, 5.325842e-06, 4.254245e-06, 4.761953e-06, 3.809081e-06, 
    3.137962e-06, 2.90466e-06, 2.648231e-06, 6.803694e-06, 6.998239e-06, 
    6.65304e-06, 6.198154e-06, 5.799109e-06, 5.301337e-06, 5.252479e-06, 
    5.163936e-06, 4.940371e-06, 4.758681e-06, 5.136165e-06, 4.714025e-06, 
    6.462441e-06, 5.489817e-06, 7.072903e-06, 6.561621e-06, 6.224267e-06, 
    6.370522e-06, 5.640556e-06, 5.478873e-06, 4.860668e-06, 5.172603e-06, 
    3.539418e-06, 4.197388e-06, 2.464405e-06, 2.769171e-06, 7.067245e-06, 
    6.804378e-06, 5.950262e-06, 6.345094e-06, 5.269423e-06, 5.029083e-06, 
    4.840514e-06, 4.608056e-06, 4.583553e-06, 4.450907e-06, 4.669997e-06, 
    4.459406e-06, 5.300317e-06, 4.909522e-06, 6.043284e-06, 5.749292e-06, 
    5.883066e-06, 6.032686e-06, 5.580662e-06, 5.130026e-06, 5.120794e-06, 
    4.983041e-06, 4.611299e-06, 5.265393e-06, 3.142881e-06, 4.498887e-06, 
    6.526763e-06, 6.058715e-06, 5.994226e-06, 6.170636e-06, 5.052758e-06, 
    5.436718e-06, 4.454109e-06, 4.703717e-06, 4.300679e-06, 4.497142e-06, 
    4.526675e-06, 4.791527e-06, 4.962869e-06, 5.41859e-06, 5.814376e-06, 
    6.1448e-06, 6.066642e-06, 5.708264e-06, 5.103482e-06, 4.581316e-06, 
    4.691684e-06, 4.330248e-06, 5.341999e-06, 4.896037e-06, 5.064567e-06, 
    4.634972e-06, 5.618994e-06, 4.771066e-06, 5.854551e-06, 5.752133e-06, 
    5.444577e-06, 4.866911e-06, 4.746341e-06, 4.620281e-06, 4.697742e-06, 
    5.088858e-06, 5.155474e-06, 5.451903e-06, 5.536148e-06, 5.77431e-06, 
    5.977742e-06, 5.791632e-06, 5.601301e-06, 5.088711e-06, 4.660709e-06, 
    4.228978e-06, 4.128677e-06, 3.677283e-06, 4.041236e-06, 3.139014e-06, 
    3.948378e-06, 2.891593e-06, 4.725474e-06, 3.963821e-06, 5.430931e-06, 
    5.253836e-06, 4.945604e-06, 4.295451e-06, 4.636919e-06, 4.239765e-06, 
    5.158102e-06, 5.696184e-06, 5.842741e-06, 6.124273e-06, 5.83643e-06, 
    5.859424e-06, 5.593573e-06, 5.677907e-06, 5.072383e-06, 5.390639e-06, 
    4.527405e-06, 4.242796e-06, 3.520356e-06, 2.892688e-06, 2.613904e-06, 
    2.497263e-06, 2.462529e-06, 2.448112e-06,
  7.925084e-09, 6.760619e-09, 6.97744e-09, 6.107188e-09, 6.580481e-09, 
    6.024294e-09, 7.679049e-09, 6.71686e-09, 7.321225e-09, 7.815244e-09, 
    4.629064e-09, 6.070151e-09, 3.391637e-09, 4.121665e-09, 2.456743e-09, 
    3.499141e-09, 2.274772e-09, 2.483586e-09, 1.890341e-09, 2.049667e-09, 
    1.400645e-09, 1.819596e-09, 1.122215e-09, 1.494336e-09, 1.431953e-09, 
    1.834631e-09, 5.759393e-09, 4.79461e-09, 5.820228e-09, 5.674473e-09, 
    5.739595e-09, 6.570428e-09, 7.017646e-09, 8.019289e-09, 7.830821e-09, 
    7.098431e-09, 5.609728e-09, 6.089274e-09, 4.929698e-09, 4.954125e-09, 
    3.84182e-09, 4.320449e-09, 2.715378e-09, 3.122892e-09, 2.042851e-09, 
    2.286885e-09, 2.053908e-09, 2.122852e-09, 2.053019e-09, 2.418227e-09, 
    2.257009e-09, 2.59601e-09, 4.227985e-09, 3.694197e-09, 5.430525e-09, 
    6.695209e-09, 7.635018e-09, 8.352556e-09, 8.248493e-09, 8.052501e-09, 
    7.094284e-09, 6.265569e-09, 5.67898e-09, 5.307571e-09, 4.957643e-09, 
    3.991319e-09, 3.534187e-09, 2.637396e-09, 2.786816e-09, 2.536848e-09, 
    2.312146e-09, 1.964561e-09, 2.019274e-09, 1.874996e-09, 2.543287e-09, 
    2.084527e-09, 2.874318e-09, 2.641868e-09, 4.864894e-09, 5.957354e-09, 
    6.466476e-09, 6.935394e-09, 8.169068e-09, 7.302783e-09, 7.636554e-09, 
    6.858705e-09, 6.392844e-09, 6.620551e-09, 5.297647e-09, 5.788875e-09, 
    3.508223e-09, 4.399507e-09, 2.337661e-09, 2.755716e-09, 2.244004e-09, 
    2.496621e-09, 2.074287e-09, 2.452089e-09, 1.823067e-09, 1.701705e-09, 
    1.784051e-09, 1.481286e-09, 2.474235e-09, 2.053891e-09, 6.62699e-09, 
    6.589465e-09, 6.416542e-09, 7.199689e-09, 7.249577e-09, 8.024477e-09, 
    7.332451e-09, 7.050224e-09, 6.366532e-09, 5.983548e-09, 5.633927e-09, 
    4.913186e-09, 4.183037e-09, 3.286853e-09, 2.727253e-09, 2.389241e-09, 
    2.593077e-09, 2.412559e-09, 2.614907e-09, 2.713422e-09, 1.746535e-09, 
    2.255528e-09, 1.522609e-09, 1.558403e-09, 1.871642e-09, 1.554343e-09, 
    6.563206e-09, 6.780501e-09, 7.571822e-09, 6.947622e-09, 8.112059e-09, 
    7.445428e-09, 7.079154e-09, 5.778236e-09, 5.515522e-09, 5.278965e-09, 
    4.831661e-09, 4.295052e-09, 3.450818e-09, 2.811215e-09, 2.299495e-09, 
    2.33475e-09, 2.322297e-09, 2.216247e-09, 2.484835e-09, 2.174041e-09, 
    2.124473e-09, 2.255616e-09, 1.563237e-09, 1.744475e-09, 1.55917e-09, 
    1.675525e-09, 6.709363e-09, 6.348987e-09, 6.542075e-09, 6.182119e-09, 
    6.434275e-09, 5.36315e-09, 5.066677e-09, 3.822023e-09, 4.305202e-09, 
    3.553739e-09, 4.224559e-09, 4.100122e-09, 3.530686e-09, 4.186374e-09, 
    2.84424e-09, 3.71698e-09, 2.21219e-09, 2.958247e-09, 2.170029e-09, 
    2.301566e-09, 2.086503e-09, 1.905298e-09, 1.692239e-09, 1.340733e-09, 
    1.417466e-09, 1.153174e-09, 5.835941e-09, 5.412454e-09, 5.44896e-09, 
    5.026166e-09, 4.727767e-09, 4.121506e-09, 3.259272e-09, 3.568096e-09, 
    3.014986e-09, 2.911148e-09, 3.757187e-09, 3.221103e-09, 5.140719e-09, 
    4.790216e-09, 4.996987e-09, 5.801728e-09, 3.495245e-09, 4.583522e-09, 
    2.718561e-09, 3.200947e-09, 1.930481e-09, 2.510464e-09, 1.460884e-09, 
    1.115764e-09, 8.456971e-10, 5.885503e-10, 5.190195e-09, 5.467928e-09, 
    4.977391e-09, 4.347643e-09, 3.812385e-09, 3.170039e-09, 3.108644e-09, 
    2.998187e-09, 2.724062e-09, 2.506591e-09, 2.963758e-09, 2.453907e-09, 
    4.711122e-09, 3.409731e-09, 5.575368e-09, 4.849257e-09, 4.383249e-09, 
    4.583931e-09, 3.604571e-09, 3.395692e-09, 2.628057e-09, 3.008952e-09, 
    1.1972e-09, 1.86833e-09, 4.315431e-10, 7.044576e-10, 5.56721e-09, 
    5.191165e-09, 4.013129e-09, 4.548889e-09, 3.129901e-09, 2.831998e-09, 
    2.60393e-09, 2.33014e-09, 2.301779e-09, 2.149968e-09, 2.402268e-09, 
    2.159605e-09, 3.168753e-09, 2.686793e-09, 4.137902e-09, 3.74678e-09, 
    3.923578e-09, 4.12364e-09, 3.526829e-09, 2.956162e-09, 2.944747e-09, 
    2.775839e-09, 2.333901e-09, 3.124842e-09, 1.121811e-09, 2.204539e-09, 
    4.800603e-09, 4.158689e-09, 4.071985e-09, 4.310196e-09, 2.860993e-09, 
    3.341754e-09, 2.153596e-09, 2.44179e-09, 1.981681e-09, 2.202548e-09, 
    2.236322e-09, 2.545538e-09, 2.751328e-09, 3.318626e-09, 3.832547e-09, 
    4.275107e-09, 4.169377e-09, 3.692962e-09, 2.923375e-09, 2.299194e-09, 
    2.427666e-09, 2.014488e-09, 3.221368e-09, 2.670546e-09, 2.875484e-09, 
    2.361407e-09, 3.576534e-09, 2.521258e-09, 3.885725e-09, 3.750514e-09, 
    3.351793e-09, 2.635543e-09, 2.492002e-09, 2.344327e-09, 2.434773e-09, 
    2.905354e-09, 2.987685e-09, 3.361158e-09, 3.469327e-09, 3.779692e-09, 
    4.049894e-09, 3.802521e-09, 3.55357e-09, 2.905173e-09, 2.391413e-09, 
    1.902787e-09, 1.794036e-09, 1.329886e-09, 1.700812e-09, 1.117056e-09, 
    1.603491e-09, 8.315635e-10, 2.467385e-09, 1.619554e-09, 3.334366e-09, 
    3.110346e-09, 2.730397e-09, 1.975896e-09, 2.363673e-09, 1.914596e-09, 
    2.990946e-09, 3.677153e-09, 3.870073e-09, 4.247277e-09, 3.861717e-09, 
    3.892187e-09, 3.543551e-09, 3.653266e-09, 2.885086e-09, 3.283048e-09, 
    2.237159e-09, 1.917918e-09, 1.17922e-09, 8.327443e-10, 5.574495e-10, 
    4.578662e-10, 4.300631e-10, 4.187762e-10,
  4.3211e-13, 4.275388e-13, 4.283906e-13, 4.249701e-13, 4.268309e-13, 
    4.24644e-13, 4.311448e-13, 4.273669e-13, 4.297405e-13, 4.316792e-13, 
    4.191484e-13, 4.248244e-13, 4.142612e-13, 4.171461e-13, 4.105594e-13, 
    4.146863e-13, 4.098377e-13, 4.106659e-13, 4.083116e-13, 4.089443e-13, 
    4.063643e-13, 4.080305e-13, 4.052605e-13, 4.067371e-13, 4.064889e-13, 
    4.080902e-13, 4.236017e-13, 4.198012e-13, 4.238411e-13, 4.232674e-13, 
    4.235237e-13, 4.267914e-13, 4.285485e-13, 4.324795e-13, 4.317403e-13, 
    4.288657e-13, 4.230126e-13, 4.248996e-13, 4.203338e-13, 4.204301e-13, 
    4.160408e-13, 4.179308e-13, 4.115845e-13, 4.13198e-13, 4.089173e-13, 
    4.098858e-13, 4.089612e-13, 4.092349e-13, 4.089576e-13, 4.104067e-13, 
    4.097673e-13, 4.111115e-13, 4.175658e-13, 4.154574e-13, 4.22307e-13, 
    4.272818e-13, 4.309721e-13, 4.337861e-13, 4.333782e-13, 4.326097e-13, 
    4.288494e-13, 4.255929e-13, 4.232852e-13, 4.218227e-13, 4.204439e-13, 
    4.166314e-13, 4.148249e-13, 4.112755e-13, 4.118675e-13, 4.10877e-13, 
    4.09986e-13, 4.086064e-13, 4.088237e-13, 4.082506e-13, 4.109025e-13, 
    4.090827e-13, 4.12214e-13, 4.112932e-13, 4.200783e-13, 4.243806e-13, 
    4.263828e-13, 4.282254e-13, 4.330668e-13, 4.296681e-13, 4.309781e-13, 
    4.279241e-13, 4.260934e-13, 4.269884e-13, 4.217836e-13, 4.237177e-13, 
    4.147222e-13, 4.182428e-13, 4.100872e-13, 4.117443e-13, 4.097157e-13, 
    4.107175e-13, 4.090421e-13, 4.10541e-13, 4.080443e-13, 4.075619e-13, 
    4.078892e-13, 4.066852e-13, 4.106288e-13, 4.089611e-13, 4.270137e-13, 
    4.268662e-13, 4.261865e-13, 4.292633e-13, 4.294592e-13, 4.324998e-13, 
    4.297846e-13, 4.286764e-13, 4.259899e-13, 4.244837e-13, 4.231078e-13, 
    4.202687e-13, 4.173884e-13, 4.138467e-13, 4.116315e-13, 4.102918e-13, 
    4.110999e-13, 4.103842e-13, 4.111864e-13, 4.115768e-13, 4.077401e-13, 
    4.097614e-13, 4.068496e-13, 4.06992e-13, 4.082373e-13, 4.069759e-13, 
    4.26763e-13, 4.276169e-13, 4.307241e-13, 4.282734e-13, 4.328433e-13, 
    4.30228e-13, 4.2879e-13, 4.236758e-13, 4.226417e-13, 4.217101e-13, 
    4.199473e-13, 4.178306e-13, 4.144952e-13, 4.119641e-13, 4.099358e-13, 
    4.100757e-13, 4.100263e-13, 4.096055e-13, 4.106708e-13, 4.094381e-13, 
    4.092413e-13, 4.097617e-13, 4.070113e-13, 4.077319e-13, 4.069951e-13, 
    4.074578e-13, 4.273374e-13, 4.259209e-13, 4.2668e-13, 4.252647e-13, 
    4.262562e-13, 4.220416e-13, 4.208736e-13, 4.159626e-13, 4.178706e-13, 
    4.149022e-13, 4.175523e-13, 4.17061e-13, 4.148111e-13, 4.174016e-13, 
    4.120949e-13, 4.155475e-13, 4.095894e-13, 4.125463e-13, 4.094221e-13, 
    4.09944e-13, 4.090906e-13, 4.08371e-13, 4.075243e-13, 4.061258e-13, 
    4.064312e-13, 4.053786e-13, 4.239029e-13, 4.222358e-13, 4.223796e-13, 
    4.20714e-13, 4.195377e-13, 4.171455e-13, 4.137376e-13, 4.14959e-13, 
    4.127709e-13, 4.123598e-13, 4.157064e-13, 4.135865e-13, 4.211654e-13, 
    4.197839e-13, 4.20599e-13, 4.237683e-13, 4.146709e-13, 4.189688e-13, 
    4.115971e-13, 4.135068e-13, 4.08471e-13, 4.107724e-13, 4.06604e-13, 
    4.052348e-13, 4.041564e-13, 4.031282e-13, 4.213603e-13, 4.224543e-13, 
    4.205218e-13, 4.180381e-13, 4.159245e-13, 4.133845e-13, 4.131416e-13, 
    4.127044e-13, 4.116189e-13, 4.107571e-13, 4.125681e-13, 4.105482e-13, 
    4.19472e-13, 4.143328e-13, 4.228773e-13, 4.200167e-13, 4.181786e-13, 
    4.189704e-13, 4.151032e-13, 4.142772e-13, 4.112385e-13, 4.12747e-13, 
    4.055541e-13, 4.082241e-13, 4.024996e-13, 4.035918e-13, 4.228452e-13, 
    4.213642e-13, 4.167175e-13, 4.188322e-13, 4.132257e-13, 4.120464e-13, 
    4.111429e-13, 4.100574e-13, 4.099449e-13, 4.093425e-13, 4.103434e-13, 
    4.093808e-13, 4.133794e-13, 4.114712e-13, 4.172102e-13, 4.156653e-13, 
    4.163638e-13, 4.171539e-13, 4.147958e-13, 4.125381e-13, 4.124929e-13, 
    4.11824e-13, 4.100723e-13, 4.132057e-13, 4.052589e-13, 4.095591e-13, 
    4.198249e-13, 4.172923e-13, 4.169499e-13, 4.178903e-13, 4.121612e-13, 
    4.140639e-13, 4.093569e-13, 4.105002e-13, 4.086744e-13, 4.095512e-13, 
    4.096852e-13, 4.109115e-13, 4.117269e-13, 4.139724e-13, 4.160041e-13, 
    4.177518e-13, 4.173345e-13, 4.154526e-13, 4.124083e-13, 4.099346e-13, 
    4.104442e-13, 4.088047e-13, 4.135876e-13, 4.114069e-13, 4.122186e-13, 
    4.101814e-13, 4.149923e-13, 4.108152e-13, 4.162142e-13, 4.1568e-13, 
    4.141036e-13, 4.112682e-13, 4.106992e-13, 4.101136e-13, 4.104723e-13, 
    4.123369e-13, 4.126629e-13, 4.141406e-13, 4.145684e-13, 4.157953e-13, 
    4.168627e-13, 4.158855e-13, 4.149015e-13, 4.123362e-13, 4.103004e-13, 
    4.08361e-13, 4.079289e-13, 4.060826e-13, 4.075584e-13, 4.0524e-13, 
    4.071714e-13, 4.041e-13, 4.106016e-13, 4.072353e-13, 4.140347e-13, 
    4.131483e-13, 4.11644e-13, 4.086514e-13, 4.101904e-13, 4.084079e-13, 
    4.126758e-13, 4.153901e-13, 4.161524e-13, 4.17642e-13, 4.161194e-13, 
    4.162398e-13, 4.148619e-13, 4.152957e-13, 4.122567e-13, 4.138316e-13, 
    4.096885e-13, 4.084211e-13, 4.054824e-13, 4.041047e-13, 4.030037e-13, 
    4.02605e-13, 4.024937e-13, 4.024484e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  9.300609e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300608e-07, 9.300609e-07, 9.300608e-07, 9.300608e-07, 9.300609e-07, 
    9.300607e-07, 9.300608e-07, 9.300606e-07, 9.300607e-07, 9.300605e-07, 
    9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300604e-07, 9.300605e-07, 
    9.300604e-07, 9.300604e-07, 9.300603e-07, 9.300604e-07, 9.300604e-07, 
    9.300604e-07, 9.300608e-07, 9.300607e-07, 9.300608e-07, 9.300608e-07, 
    9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300609e-07, 9.300609e-07, 
    9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300607e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300605e-07, 9.300606e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300607e-07, 9.300606e-07, 9.300608e-07, 
    9.300608e-07, 9.300609e-07, 9.300609e-07, 9.300609e-07, 9.300609e-07, 
    9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300607e-07, 9.300607e-07, 
    9.300607e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300604e-07, 9.300605e-07, 9.300604e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300607e-07, 9.300608e-07, 
    9.300608e-07, 9.300608e-07, 9.300609e-07, 9.300608e-07, 9.300609e-07, 
    9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300607e-07, 9.300608e-07, 
    9.300606e-07, 9.300607e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300604e-07, 9.300604e-07, 
    9.300604e-07, 9.300604e-07, 9.300605e-07, 9.300605e-07, 9.300608e-07, 
    9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300609e-07, 
    9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300604e-07, 
    9.300605e-07, 9.300604e-07, 9.300604e-07, 9.300604e-07, 9.300604e-07, 
    9.300608e-07, 9.300608e-07, 9.300609e-07, 9.300608e-07, 9.300609e-07, 
    9.300609e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300604e-07, 9.300604e-07, 9.300604e-07, 
    9.300604e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300608e-07, 9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300607e-07, 
    9.300606e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300607e-07, 
    9.300605e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300604e-07, 9.300604e-07, 9.300604e-07, 
    9.300604e-07, 9.300603e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300606e-07, 
    9.300605e-07, 9.300605e-07, 9.300606e-07, 9.300606e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300608e-07, 9.300606e-07, 9.300607e-07, 
    9.300605e-07, 9.300606e-07, 9.300604e-07, 9.300605e-07, 9.300604e-07, 
    9.300603e-07, 9.300603e-07, 9.300602e-07, 9.300607e-07, 9.300608e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300606e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300607e-07, 9.300606e-07, 9.300608e-07, 9.300607e-07, 9.300607e-07, 
    9.300607e-07, 9.300606e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 
    9.300604e-07, 9.300604e-07, 9.300602e-07, 9.300603e-07, 9.300608e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300606e-07, 9.300605e-07, 9.300607e-07, 9.300606e-07, 
    9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300606e-07, 9.300603e-07, 9.300605e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300605e-07, 
    9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300604e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300606e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300606e-07, 9.300605e-07, 9.300607e-07, 9.300606e-07, 
    9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300606e-07, 9.300606e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 
    9.300604e-07, 9.300604e-07, 9.300604e-07, 9.300604e-07, 9.300603e-07, 
    9.300604e-07, 9.300603e-07, 9.300605e-07, 9.300604e-07, 9.300606e-07, 
    9.300606e-07, 9.300605e-07, 9.300604e-07, 9.300605e-07, 9.300604e-07, 
    9.300605e-07, 9.300606e-07, 9.300607e-07, 9.300607e-07, 9.300607e-07, 
    9.300607e-07, 9.300606e-07, 9.300606e-07, 9.300605e-07, 9.300606e-07, 
    9.300605e-07, 9.300604e-07, 9.300603e-07, 9.300603e-07, 9.300602e-07, 
    9.300602e-07, 9.300602e-07, 9.300602e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.333051e-16, 6.350136e-16, 6.346817e-16, 6.360584e-16, 6.35295e-16, 
    6.361961e-16, 6.336519e-16, 6.350812e-16, 6.34169e-16, 6.334594e-16, 
    6.38726e-16, 6.361198e-16, 6.414308e-16, 6.397716e-16, 6.439366e-16, 
    6.411724e-16, 6.444935e-16, 6.438574e-16, 6.457725e-16, 6.452241e-16, 
    6.476698e-16, 6.460255e-16, 6.48937e-16, 6.472776e-16, 6.475371e-16, 
    6.459711e-16, 6.366451e-16, 6.384016e-16, 6.365409e-16, 6.367915e-16, 
    6.366791e-16, 6.353106e-16, 6.346202e-16, 6.331749e-16, 6.334374e-16, 
    6.344991e-16, 6.369042e-16, 6.360885e-16, 6.381445e-16, 6.38098e-16, 
    6.403835e-16, 6.393534e-16, 6.431899e-16, 6.421008e-16, 6.45247e-16, 
    6.444562e-16, 6.452098e-16, 6.449813e-16, 6.452127e-16, 6.440528e-16, 
    6.445498e-16, 6.435289e-16, 6.395463e-16, 6.407177e-16, 6.372211e-16, 
    6.351141e-16, 6.337145e-16, 6.327202e-16, 6.328608e-16, 6.331287e-16, 
    6.345053e-16, 6.357991e-16, 6.367842e-16, 6.374427e-16, 6.380914e-16, 
    6.400519e-16, 6.410897e-16, 6.434098e-16, 6.429918e-16, 6.437003e-16, 
    6.443775e-16, 6.455133e-16, 6.453265e-16, 6.458265e-16, 6.436819e-16, 
    6.451074e-16, 6.427534e-16, 6.433975e-16, 6.38266e-16, 6.363087e-16, 
    6.354746e-16, 6.347454e-16, 6.329689e-16, 6.341959e-16, 6.337122e-16, 
    6.348629e-16, 6.355934e-16, 6.352322e-16, 6.374607e-16, 6.365946e-16, 
    6.411512e-16, 6.391901e-16, 6.442985e-16, 6.430776e-16, 6.445911e-16, 
    6.43819e-16, 6.451415e-16, 6.439514e-16, 6.460127e-16, 6.46461e-16, 
    6.461546e-16, 6.473318e-16, 6.438853e-16, 6.452096e-16, 6.35222e-16, 
    6.352809e-16, 6.355555e-16, 6.343481e-16, 6.342744e-16, 6.331676e-16, 
    6.341526e-16, 6.345717e-16, 6.356359e-16, 6.362647e-16, 6.368623e-16, 
    6.381756e-16, 6.396408e-16, 6.416878e-16, 6.431568e-16, 6.441408e-16, 
    6.435376e-16, 6.440701e-16, 6.434747e-16, 6.431957e-16, 6.46293e-16, 
    6.445544e-16, 6.471626e-16, 6.470184e-16, 6.458383e-16, 6.470347e-16, 
    6.353223e-16, 6.349833e-16, 6.338051e-16, 6.347272e-16, 6.330471e-16, 
    6.339875e-16, 6.345279e-16, 6.366123e-16, 6.370704e-16, 6.374945e-16, 
    6.383321e-16, 6.394062e-16, 6.412885e-16, 6.429245e-16, 6.44417e-16, 
    6.443077e-16, 6.443462e-16, 6.446792e-16, 6.438538e-16, 6.448147e-16, 
    6.449757e-16, 6.445544e-16, 6.469991e-16, 6.463011e-16, 6.470153e-16, 
    6.465609e-16, 6.350936e-16, 6.35664e-16, 6.353557e-16, 6.359352e-16, 
    6.355269e-16, 6.373415e-16, 6.378852e-16, 6.404272e-16, 6.393849e-16, 
    6.41044e-16, 6.395537e-16, 6.398177e-16, 6.410973e-16, 6.396343e-16, 
    6.42834e-16, 6.406649e-16, 6.446922e-16, 6.425279e-16, 6.448277e-16, 
    6.444105e-16, 6.451013e-16, 6.457195e-16, 6.464972e-16, 6.479307e-16, 
    6.475989e-16, 6.487973e-16, 6.365142e-16, 6.372533e-16, 6.371886e-16, 
    6.37962e-16, 6.385336e-16, 6.397722e-16, 6.417565e-16, 6.410108e-16, 
    6.4238e-16, 6.426543e-16, 6.405745e-16, 6.418517e-16, 6.37748e-16, 
    6.384114e-16, 6.380167e-16, 6.365724e-16, 6.411822e-16, 6.388178e-16, 
    6.43181e-16, 6.419026e-16, 6.456313e-16, 6.437775e-16, 6.474162e-16, 
    6.489683e-16, 6.504291e-16, 6.521326e-16, 6.376569e-16, 6.371548e-16, 
    6.38054e-16, 6.392966e-16, 6.404495e-16, 6.419806e-16, 6.421373e-16, 
    6.424238e-16, 6.431659e-16, 6.437896e-16, 6.425141e-16, 6.43946e-16, 
    6.385645e-16, 6.413874e-16, 6.369646e-16, 6.382973e-16, 6.392235e-16, 
    6.388176e-16, 6.409256e-16, 6.414219e-16, 6.434366e-16, 6.423958e-16, 
    6.48585e-16, 6.458495e-16, 6.534295e-16, 6.513149e-16, 6.369793e-16, 
    6.376553e-16, 6.400054e-16, 6.388877e-16, 6.420829e-16, 6.428679e-16, 
    6.435063e-16, 6.443216e-16, 6.444098e-16, 6.448926e-16, 6.441013e-16, 
    6.448615e-16, 6.419838e-16, 6.432703e-16, 6.397374e-16, 6.405978e-16, 
    6.402022e-16, 6.397678e-16, 6.41108e-16, 6.425338e-16, 6.425648e-16, 
    6.430217e-16, 6.443075e-16, 6.420958e-16, 6.489367e-16, 6.447144e-16, 
    6.383922e-16, 6.396921e-16, 6.398784e-16, 6.393749e-16, 6.427892e-16, 
    6.41553e-16, 6.448809e-16, 6.439822e-16, 6.454546e-16, 6.44723e-16, 
    6.446154e-16, 6.436754e-16, 6.430898e-16, 6.416097e-16, 6.404042e-16, 
    6.39448e-16, 6.396704e-16, 6.407207e-16, 6.426211e-16, 6.444175e-16, 
    6.440241e-16, 6.453428e-16, 6.418514e-16, 6.433159e-16, 6.427497e-16, 
    6.442256e-16, 6.409908e-16, 6.437441e-16, 6.40286e-16, 6.405896e-16, 
    6.415285e-16, 6.434148e-16, 6.438327e-16, 6.442778e-16, 6.440033e-16, 
    6.426694e-16, 6.424514e-16, 6.415058e-16, 6.412444e-16, 6.405236e-16, 
    6.399263e-16, 6.404718e-16, 6.410445e-16, 6.426702e-16, 6.441338e-16, 
    6.457282e-16, 6.461184e-16, 6.479773e-16, 6.464635e-16, 6.489601e-16, 
    6.468366e-16, 6.505112e-16, 6.439044e-16, 6.467752e-16, 6.415714e-16, 
    6.42133e-16, 6.431474e-16, 6.454735e-16, 6.442187e-16, 6.456863e-16, 
    6.424428e-16, 6.407566e-16, 6.403207e-16, 6.39506e-16, 6.403393e-16, 
    6.402716e-16, 6.410686e-16, 6.408126e-16, 6.427242e-16, 6.416978e-16, 
    6.446125e-16, 6.456748e-16, 6.486715e-16, 6.505054e-16, 6.523707e-16, 
    6.531932e-16, 6.534435e-16, 6.53548e-16 ;

 CWDC_TO_LITR2C =
  4.813119e-16, 4.826103e-16, 4.823581e-16, 4.834043e-16, 4.828242e-16, 
    4.835091e-16, 4.815754e-16, 4.826617e-16, 4.819685e-16, 4.814291e-16, 
    4.854317e-16, 4.83451e-16, 4.874874e-16, 4.862264e-16, 4.893918e-16, 
    4.87291e-16, 4.898151e-16, 4.893316e-16, 4.90787e-16, 4.903703e-16, 
    4.922291e-16, 4.909794e-16, 4.931921e-16, 4.91931e-16, 4.921282e-16, 
    4.90938e-16, 4.838503e-16, 4.851852e-16, 4.837711e-16, 4.839615e-16, 
    4.838761e-16, 4.82836e-16, 4.823114e-16, 4.812129e-16, 4.814124e-16, 
    4.822194e-16, 4.840472e-16, 4.834273e-16, 4.849898e-16, 4.849545e-16, 
    4.866914e-16, 4.859086e-16, 4.888243e-16, 4.879966e-16, 4.903877e-16, 
    4.897867e-16, 4.903594e-16, 4.901859e-16, 4.903617e-16, 4.894801e-16, 
    4.898579e-16, 4.89082e-16, 4.860552e-16, 4.869455e-16, 4.84288e-16, 
    4.826868e-16, 4.81623e-16, 4.808674e-16, 4.809742e-16, 4.811778e-16, 
    4.822241e-16, 4.832073e-16, 4.83956e-16, 4.844565e-16, 4.849494e-16, 
    4.864394e-16, 4.872282e-16, 4.889915e-16, 4.886737e-16, 4.892122e-16, 
    4.897269e-16, 4.905901e-16, 4.904481e-16, 4.908282e-16, 4.891983e-16, 
    4.902816e-16, 4.884926e-16, 4.889822e-16, 4.850821e-16, 4.835946e-16, 
    4.829607e-16, 4.824065e-16, 4.810563e-16, 4.819889e-16, 4.816213e-16, 
    4.824958e-16, 4.83051e-16, 4.827765e-16, 4.844701e-16, 4.838119e-16, 
    4.872749e-16, 4.857845e-16, 4.896669e-16, 4.88739e-16, 4.898892e-16, 
    4.893025e-16, 4.903076e-16, 4.89403e-16, 4.909697e-16, 4.913104e-16, 
    4.910775e-16, 4.919722e-16, 4.893529e-16, 4.903593e-16, 4.827687e-16, 
    4.828135e-16, 4.830222e-16, 4.821046e-16, 4.820485e-16, 4.812074e-16, 
    4.819559e-16, 4.822745e-16, 4.830833e-16, 4.835612e-16, 4.840154e-16, 
    4.850135e-16, 4.86127e-16, 4.876827e-16, 4.887992e-16, 4.89547e-16, 
    4.890886e-16, 4.894933e-16, 4.890408e-16, 4.888287e-16, 4.911827e-16, 
    4.898613e-16, 4.918436e-16, 4.91734e-16, 4.908371e-16, 4.917464e-16, 
    4.828449e-16, 4.825873e-16, 4.816919e-16, 4.823927e-16, 4.811158e-16, 
    4.818305e-16, 4.822412e-16, 4.838254e-16, 4.841735e-16, 4.844958e-16, 
    4.851324e-16, 4.859487e-16, 4.873793e-16, 4.886226e-16, 4.897569e-16, 
    4.896739e-16, 4.897031e-16, 4.899562e-16, 4.893289e-16, 4.900592e-16, 
    4.901816e-16, 4.898613e-16, 4.917193e-16, 4.911888e-16, 4.917316e-16, 
    4.913863e-16, 4.826711e-16, 4.831047e-16, 4.828703e-16, 4.833108e-16, 
    4.830004e-16, 4.843796e-16, 4.847927e-16, 4.867247e-16, 4.859325e-16, 
    4.871934e-16, 4.860608e-16, 4.862614e-16, 4.872339e-16, 4.861221e-16, 
    4.885538e-16, 4.869053e-16, 4.89966e-16, 4.883212e-16, 4.90069e-16, 
    4.89752e-16, 4.90277e-16, 4.907468e-16, 4.913379e-16, 4.924273e-16, 
    4.921752e-16, 4.930859e-16, 4.837508e-16, 4.843125e-16, 4.842633e-16, 
    4.848511e-16, 4.852855e-16, 4.862269e-16, 4.87735e-16, 4.871681e-16, 
    4.882088e-16, 4.884172e-16, 4.868366e-16, 4.878072e-16, 4.846885e-16, 
    4.851926e-16, 4.848927e-16, 4.83795e-16, 4.872985e-16, 4.855016e-16, 
    4.888175e-16, 4.87846e-16, 4.906798e-16, 4.89271e-16, 4.920363e-16, 
    4.932159e-16, 4.943261e-16, 4.956208e-16, 4.846193e-16, 4.842377e-16, 
    4.84921e-16, 4.858654e-16, 4.867417e-16, 4.879052e-16, 4.880243e-16, 
    4.882421e-16, 4.88806e-16, 4.892801e-16, 4.883107e-16, 4.89399e-16, 
    4.853091e-16, 4.874544e-16, 4.840931e-16, 4.85106e-16, 4.858099e-16, 
    4.855014e-16, 4.871034e-16, 4.874806e-16, 4.890118e-16, 4.882208e-16, 
    4.929246e-16, 4.908457e-16, 4.966064e-16, 4.949993e-16, 4.841043e-16, 
    4.84618e-16, 4.864041e-16, 4.855547e-16, 4.87983e-16, 4.885796e-16, 
    4.890648e-16, 4.896844e-16, 4.897514e-16, 4.901184e-16, 4.89517e-16, 
    4.900947e-16, 4.879077e-16, 4.888854e-16, 4.862004e-16, 4.868544e-16, 
    4.865537e-16, 4.862235e-16, 4.872421e-16, 4.883257e-16, 4.883492e-16, 
    4.886965e-16, 4.896737e-16, 4.879928e-16, 4.931919e-16, 4.899829e-16, 
    4.85178e-16, 4.86166e-16, 4.863076e-16, 4.859249e-16, 4.885198e-16, 
    4.875803e-16, 4.901095e-16, 4.894265e-16, 4.905455e-16, 4.899895e-16, 
    4.899077e-16, 4.891933e-16, 4.887482e-16, 4.876233e-16, 4.867072e-16, 
    4.859804e-16, 4.861495e-16, 4.869477e-16, 4.883921e-16, 4.897573e-16, 
    4.894583e-16, 4.904605e-16, 4.878071e-16, 4.889201e-16, 4.884898e-16, 
    4.896115e-16, 4.87153e-16, 4.892455e-16, 4.866174e-16, 4.868481e-16, 
    4.875616e-16, 4.889952e-16, 4.893128e-16, 4.896511e-16, 4.894425e-16, 
    4.884287e-16, 4.88263e-16, 4.875444e-16, 4.873457e-16, 4.867979e-16, 
    4.86344e-16, 4.867586e-16, 4.871938e-16, 4.884294e-16, 4.895417e-16, 
    4.907535e-16, 4.910499e-16, 4.924628e-16, 4.913122e-16, 4.932097e-16, 
    4.915958e-16, 4.943885e-16, 4.893673e-16, 4.915492e-16, 4.875943e-16, 
    4.880211e-16, 4.88792e-16, 4.905598e-16, 4.896062e-16, 4.907215e-16, 
    4.882566e-16, 4.86975e-16, 4.866437e-16, 4.860246e-16, 4.866579e-16, 
    4.866064e-16, 4.872121e-16, 4.870175e-16, 4.884703e-16, 4.876903e-16, 
    4.899055e-16, 4.907129e-16, 4.929904e-16, 4.943841e-16, 4.958017e-16, 
    4.964268e-16, 4.96617e-16, 4.966965e-16 ;

 CWDC_TO_LITR3C =
  1.519932e-16, 1.524033e-16, 1.523236e-16, 1.52654e-16, 1.524708e-16, 
    1.526871e-16, 1.520765e-16, 1.524195e-16, 1.522006e-16, 1.520302e-16, 
    1.532942e-16, 1.526687e-16, 1.539434e-16, 1.535452e-16, 1.545448e-16, 
    1.538814e-16, 1.546784e-16, 1.545258e-16, 1.549854e-16, 1.548538e-16, 
    1.554408e-16, 1.550461e-16, 1.557449e-16, 1.553466e-16, 1.554089e-16, 
    1.550331e-16, 1.527948e-16, 1.532164e-16, 1.527698e-16, 1.5283e-16, 
    1.52803e-16, 1.524745e-16, 1.523088e-16, 1.51962e-16, 1.52025e-16, 
    1.522798e-16, 1.52857e-16, 1.526612e-16, 1.531547e-16, 1.531435e-16, 
    1.53692e-16, 1.534448e-16, 1.543656e-16, 1.541042e-16, 1.548593e-16, 
    1.546695e-16, 1.548503e-16, 1.547955e-16, 1.548511e-16, 1.545727e-16, 
    1.54692e-16, 1.544469e-16, 1.534911e-16, 1.537723e-16, 1.529331e-16, 
    1.524274e-16, 1.520915e-16, 1.518529e-16, 1.518866e-16, 1.519509e-16, 
    1.522813e-16, 1.525918e-16, 1.528282e-16, 1.529862e-16, 1.531419e-16, 
    1.536125e-16, 1.538615e-16, 1.544184e-16, 1.54318e-16, 1.544881e-16, 
    1.546506e-16, 1.549232e-16, 1.548783e-16, 1.549984e-16, 1.544837e-16, 
    1.548258e-16, 1.542608e-16, 1.544154e-16, 1.531838e-16, 1.527141e-16, 
    1.525139e-16, 1.523389e-16, 1.519125e-16, 1.52207e-16, 1.520909e-16, 
    1.523671e-16, 1.525424e-16, 1.524557e-16, 1.529906e-16, 1.527827e-16, 
    1.538763e-16, 1.534056e-16, 1.546316e-16, 1.543386e-16, 1.547019e-16, 
    1.545166e-16, 1.54834e-16, 1.545483e-16, 1.550431e-16, 1.551506e-16, 
    1.550771e-16, 1.553596e-16, 1.545325e-16, 1.548503e-16, 1.524533e-16, 
    1.524674e-16, 1.525333e-16, 1.522435e-16, 1.522258e-16, 1.519602e-16, 
    1.521966e-16, 1.522972e-16, 1.525526e-16, 1.527035e-16, 1.52847e-16, 
    1.531622e-16, 1.535138e-16, 1.540051e-16, 1.543576e-16, 1.545938e-16, 
    1.54449e-16, 1.545768e-16, 1.544339e-16, 1.54367e-16, 1.551103e-16, 
    1.54693e-16, 1.55319e-16, 1.552844e-16, 1.550012e-16, 1.552883e-16, 
    1.524774e-16, 1.52396e-16, 1.521132e-16, 1.523345e-16, 1.519313e-16, 
    1.52157e-16, 1.522867e-16, 1.52787e-16, 1.528969e-16, 1.529987e-16, 
    1.531997e-16, 1.534575e-16, 1.539092e-16, 1.543019e-16, 1.546601e-16, 
    1.546338e-16, 1.546431e-16, 1.54723e-16, 1.545249e-16, 1.547555e-16, 
    1.547942e-16, 1.54693e-16, 1.552798e-16, 1.551123e-16, 1.552837e-16, 
    1.551746e-16, 1.524224e-16, 1.525594e-16, 1.524854e-16, 1.526245e-16, 
    1.525264e-16, 1.52962e-16, 1.530925e-16, 1.537025e-16, 1.534524e-16, 
    1.538506e-16, 1.534929e-16, 1.535562e-16, 1.538633e-16, 1.535122e-16, 
    1.542801e-16, 1.537596e-16, 1.547261e-16, 1.542067e-16, 1.547586e-16, 
    1.546585e-16, 1.548243e-16, 1.549727e-16, 1.551593e-16, 1.555034e-16, 
    1.554237e-16, 1.557114e-16, 1.527634e-16, 1.529408e-16, 1.529253e-16, 
    1.531109e-16, 1.532481e-16, 1.535453e-16, 1.540216e-16, 1.538426e-16, 
    1.541712e-16, 1.54237e-16, 1.537379e-16, 1.540444e-16, 1.530595e-16, 
    1.532187e-16, 1.53124e-16, 1.527774e-16, 1.538837e-16, 1.533163e-16, 
    1.543634e-16, 1.540566e-16, 1.549515e-16, 1.545066e-16, 1.553799e-16, 
    1.557524e-16, 1.56103e-16, 1.565118e-16, 1.530377e-16, 1.529172e-16, 
    1.53133e-16, 1.534312e-16, 1.537079e-16, 1.540753e-16, 1.54113e-16, 
    1.541817e-16, 1.543598e-16, 1.545095e-16, 1.542034e-16, 1.54547e-16, 
    1.532555e-16, 1.53933e-16, 1.528715e-16, 1.531914e-16, 1.534136e-16, 
    1.533162e-16, 1.538221e-16, 1.539413e-16, 1.544248e-16, 1.54175e-16, 
    1.556604e-16, 1.550039e-16, 1.568231e-16, 1.563156e-16, 1.52875e-16, 
    1.530373e-16, 1.536013e-16, 1.533331e-16, 1.540999e-16, 1.542883e-16, 
    1.544415e-16, 1.546372e-16, 1.546583e-16, 1.547742e-16, 1.545843e-16, 
    1.547668e-16, 1.540761e-16, 1.543849e-16, 1.53537e-16, 1.537435e-16, 
    1.536485e-16, 1.535443e-16, 1.538659e-16, 1.542081e-16, 1.542155e-16, 
    1.543252e-16, 1.546338e-16, 1.54103e-16, 1.557448e-16, 1.547314e-16, 
    1.532141e-16, 1.535261e-16, 1.535708e-16, 1.5345e-16, 1.542694e-16, 
    1.539727e-16, 1.547714e-16, 1.545557e-16, 1.549091e-16, 1.547335e-16, 
    1.547077e-16, 1.544821e-16, 1.543415e-16, 1.539863e-16, 1.53697e-16, 
    1.534675e-16, 1.535209e-16, 1.53773e-16, 1.542291e-16, 1.546602e-16, 
    1.545658e-16, 1.548823e-16, 1.540443e-16, 1.543958e-16, 1.542599e-16, 
    1.546141e-16, 1.538378e-16, 1.544986e-16, 1.536686e-16, 1.537415e-16, 
    1.539668e-16, 1.544195e-16, 1.545198e-16, 1.546267e-16, 1.545608e-16, 
    1.542407e-16, 1.541883e-16, 1.539614e-16, 1.538986e-16, 1.537257e-16, 
    1.535823e-16, 1.537133e-16, 1.538507e-16, 1.542408e-16, 1.545921e-16, 
    1.549748e-16, 1.550684e-16, 1.555146e-16, 1.551512e-16, 1.557504e-16, 
    1.552408e-16, 1.561227e-16, 1.54537e-16, 1.552261e-16, 1.539771e-16, 
    1.541119e-16, 1.543554e-16, 1.549136e-16, 1.546125e-16, 1.549647e-16, 
    1.541863e-16, 1.537816e-16, 1.53677e-16, 1.534814e-16, 1.536814e-16, 
    1.536652e-16, 1.538565e-16, 1.53795e-16, 1.542538e-16, 1.540075e-16, 
    1.54707e-16, 1.54962e-16, 1.556812e-16, 1.561213e-16, 1.56569e-16, 
    1.567664e-16, 1.568264e-16, 1.568515e-16 ;

 CWDC_vr =
  5.310744e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310744e-05, 5.310743e-05, 5.310744e-05, 5.310744e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310743e-05, 5.310741e-05, 
    5.310742e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310744e-05, 5.310744e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310742e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310742e-05, 5.310743e-05, 5.310742e-05, 5.310743e-05, 
    5.310743e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310742e-05, 5.310742e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310742e-05, 5.310743e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 
    5.310744e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310743e-05, 5.310743e-05, 5.310744e-05, 5.310743e-05, 5.310744e-05, 
    5.310744e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310743e-05, 
    5.310742e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310743e-05, 
    5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310743e-05, 
    5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.31074e-05, 5.31074e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 
    5.310743e-05, 5.310742e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310741e-05, 5.310741e-05, 5.31074e-05, 5.31074e-05, 5.310743e-05, 
    5.310743e-05, 5.310742e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310742e-05, 5.310742e-05, 5.310743e-05, 5.310742e-05, 
    5.310742e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 5.310741e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 
    5.310742e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310741e-05, 5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.31074e-05, 5.310741e-05, 5.310741e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310743e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.31074e-05, 5.31074e-05, 
    5.31074e-05, 5.31074e-05, 5.31074e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860121e-09, 1.860122e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860122e-09, 1.860121e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860122e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.86012e-09, 1.860121e-09, 1.860122e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860122e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.86012e-09, 1.860121e-09, 1.860122e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.86012e-09, 
    1.86012e-09, 1.86012e-09, 1.86012e-09 ;

 CWDN_TO_LITR2N =
  9.626239e-19, 9.652206e-19, 9.647161e-19, 9.668087e-19, 9.656485e-19, 
    9.670181e-19, 9.631509e-19, 9.653234e-19, 9.639369e-19, 9.628582e-19, 
    9.708635e-19, 9.669021e-19, 9.749747e-19, 9.724529e-19, 9.787836e-19, 
    9.74582e-19, 9.796301e-19, 9.786632e-19, 9.815741e-19, 9.807406e-19, 
    9.844581e-19, 9.819587e-19, 9.863842e-19, 9.83862e-19, 9.842564e-19, 
    9.818761e-19, 9.677005e-19, 9.703704e-19, 9.675421e-19, 9.67923e-19, 
    9.677523e-19, 9.656722e-19, 9.646227e-19, 9.624258e-19, 9.628249e-19, 
    9.644387e-19, 9.680943e-19, 9.668545e-19, 9.699796e-19, 9.699091e-19, 
    9.733829e-19, 9.718172e-19, 9.776486e-19, 9.759932e-19, 9.807754e-19, 
    9.795734e-19, 9.807189e-19, 9.803717e-19, 9.807233e-19, 9.789602e-19, 
    9.797158e-19, 9.78164e-19, 9.721103e-19, 9.738909e-19, 9.685761e-19, 
    9.653735e-19, 9.63246e-19, 9.617348e-19, 9.619485e-19, 9.623557e-19, 
    9.644481e-19, 9.664147e-19, 9.67912e-19, 9.689129e-19, 9.698988e-19, 
    9.728789e-19, 9.744563e-19, 9.77983e-19, 9.773475e-19, 9.784244e-19, 
    9.794538e-19, 9.811801e-19, 9.808962e-19, 9.816563e-19, 9.783965e-19, 
    9.805633e-19, 9.769852e-19, 9.779643e-19, 9.701643e-19, 9.671892e-19, 
    9.659213e-19, 9.64813e-19, 9.621127e-19, 9.639777e-19, 9.632426e-19, 
    9.649916e-19, 9.66102e-19, 9.655529e-19, 9.689402e-19, 9.676238e-19, 
    9.745498e-19, 9.71569e-19, 9.793338e-19, 9.77478e-19, 9.797785e-19, 
    9.78605e-19, 9.806152e-19, 9.788061e-19, 9.819394e-19, 9.826208e-19, 
    9.821551e-19, 9.839444e-19, 9.787057e-19, 9.807186e-19, 9.655374e-19, 
    9.65627e-19, 9.660444e-19, 9.642092e-19, 9.64097e-19, 9.624147e-19, 
    9.639119e-19, 9.645489e-19, 9.661665e-19, 9.671223e-19, 9.680308e-19, 
    9.700269e-19, 9.722539e-19, 9.753655e-19, 9.775982e-19, 9.790941e-19, 
    9.781772e-19, 9.789867e-19, 9.780816e-19, 9.776574e-19, 9.823653e-19, 
    9.797226e-19, 9.83687e-19, 9.834679e-19, 9.816743e-19, 9.834926e-19, 
    9.656899e-19, 9.651746e-19, 9.633838e-19, 9.647853e-19, 9.622315e-19, 
    9.63661e-19, 9.644824e-19, 9.676508e-19, 9.683469e-19, 9.689915e-19, 
    9.702648e-19, 9.718973e-19, 9.747585e-19, 9.772451e-19, 9.795138e-19, 
    9.793477e-19, 9.794061e-19, 9.799124e-19, 9.786579e-19, 9.801183e-19, 
    9.803631e-19, 9.797226e-19, 9.834386e-19, 9.823776e-19, 9.834633e-19, 
    9.827726e-19, 9.653422e-19, 9.662093e-19, 9.657407e-19, 9.666216e-19, 
    9.660009e-19, 9.687592e-19, 9.695855e-19, 9.734494e-19, 9.71865e-19, 
    9.743868e-19, 9.721216e-19, 9.72523e-19, 9.744679e-19, 9.722442e-19, 
    9.771076e-19, 9.738106e-19, 9.799321e-19, 9.766424e-19, 9.801381e-19, 
    9.79504e-19, 9.80554e-19, 9.814936e-19, 9.826758e-19, 9.848547e-19, 
    9.843504e-19, 9.861719e-19, 9.675016e-19, 9.686251e-19, 9.685267e-19, 
    9.697022e-19, 9.70571e-19, 9.724538e-19, 9.754699e-19, 9.743364e-19, 
    9.764175e-19, 9.768344e-19, 9.736733e-19, 9.756146e-19, 9.69377e-19, 
    9.703853e-19, 9.697854e-19, 9.6759e-19, 9.745969e-19, 9.710031e-19, 
    9.77635e-19, 9.75692e-19, 9.813596e-19, 9.785418e-19, 9.840727e-19, 
    9.864317e-19, 9.886522e-19, 9.912415e-19, 9.692385e-19, 9.684754e-19, 
    9.698421e-19, 9.717307e-19, 9.734833e-19, 9.758105e-19, 9.760487e-19, 
    9.764842e-19, 9.776121e-19, 9.785602e-19, 9.766214e-19, 9.787979e-19, 
    9.706181e-19, 9.749089e-19, 9.681863e-19, 9.702119e-19, 9.716197e-19, 
    9.710027e-19, 9.742069e-19, 9.749613e-19, 9.780236e-19, 9.764416e-19, 
    9.858493e-19, 9.816913e-19, 9.932128e-19, 9.899986e-19, 9.682085e-19, 
    9.692361e-19, 9.728082e-19, 9.711093e-19, 9.75966e-19, 9.771592e-19, 
    9.781296e-19, 9.793687e-19, 9.795028e-19, 9.802367e-19, 9.79034e-19, 
    9.801895e-19, 9.758154e-19, 9.777708e-19, 9.724008e-19, 9.737087e-19, 
    9.731073e-19, 9.724471e-19, 9.744842e-19, 9.766513e-19, 9.766985e-19, 
    9.773929e-19, 9.793474e-19, 9.759856e-19, 9.863838e-19, 9.799658e-19, 
    9.703561e-19, 9.723321e-19, 9.726151e-19, 9.718497e-19, 9.770396e-19, 
    9.751606e-19, 9.80219e-19, 9.78853e-19, 9.81091e-19, 9.799791e-19, 
    9.798154e-19, 9.783866e-19, 9.774965e-19, 9.752467e-19, 9.734144e-19, 
    9.719609e-19, 9.72299e-19, 9.738954e-19, 9.767841e-19, 9.795146e-19, 
    9.789167e-19, 9.80921e-19, 9.756141e-19, 9.778401e-19, 9.769795e-19, 
    9.792229e-19, 9.74306e-19, 9.784912e-19, 9.732347e-19, 9.736962e-19, 
    9.751233e-19, 9.779905e-19, 9.786257e-19, 9.793022e-19, 9.78885e-19, 
    9.768575e-19, 9.765261e-19, 9.750888e-19, 9.746914e-19, 9.735958e-19, 
    9.72688e-19, 9.735172e-19, 9.743876e-19, 9.768587e-19, 9.790834e-19, 
    9.815069e-19, 9.821e-19, 9.849256e-19, 9.826245e-19, 9.864194e-19, 
    9.831916e-19, 9.88777e-19, 9.787347e-19, 9.830984e-19, 9.751885e-19, 
    9.760421e-19, 9.77584e-19, 9.811196e-19, 9.792124e-19, 9.814432e-19, 
    9.765132e-19, 9.739501e-19, 9.732875e-19, 9.720491e-19, 9.733158e-19, 
    9.732128e-19, 9.744242e-19, 9.740351e-19, 9.769407e-19, 9.753807e-19, 
    9.79811e-19, 9.814257e-19, 9.859808e-19, 9.887682e-19, 9.916034e-19, 
    9.928536e-19, 9.93234e-19, 9.93393e-19 ;

 CWDN_TO_LITR3N =
  3.039865e-19, 3.048065e-19, 3.046472e-19, 3.05308e-19, 3.049416e-19, 
    3.053741e-19, 3.041529e-19, 3.04839e-19, 3.044011e-19, 3.040605e-19, 
    3.065885e-19, 3.053375e-19, 3.078868e-19, 3.070904e-19, 3.090896e-19, 
    3.077627e-19, 3.093569e-19, 3.090516e-19, 3.099708e-19, 3.097076e-19, 
    3.108815e-19, 3.100922e-19, 3.114897e-19, 3.106932e-19, 3.108178e-19, 
    3.100661e-19, 3.055897e-19, 3.064328e-19, 3.055396e-19, 3.056599e-19, 
    3.05606e-19, 3.049491e-19, 3.046177e-19, 3.039239e-19, 3.0405e-19, 
    3.045596e-19, 3.05714e-19, 3.053225e-19, 3.063093e-19, 3.062871e-19, 
    3.073841e-19, 3.068896e-19, 3.087312e-19, 3.082084e-19, 3.097185e-19, 
    3.09339e-19, 3.097007e-19, 3.095911e-19, 3.097021e-19, 3.091453e-19, 
    3.093839e-19, 3.088939e-19, 3.069822e-19, 3.075445e-19, 3.058661e-19, 
    3.048548e-19, 3.04183e-19, 3.037057e-19, 3.037732e-19, 3.039018e-19, 
    3.045626e-19, 3.051836e-19, 3.056564e-19, 3.059725e-19, 3.062839e-19, 
    3.072249e-19, 3.077231e-19, 3.088367e-19, 3.08636e-19, 3.089761e-19, 
    3.093012e-19, 3.098464e-19, 3.097567e-19, 3.099967e-19, 3.089673e-19, 
    3.096515e-19, 3.085216e-19, 3.088308e-19, 3.063676e-19, 3.054282e-19, 
    3.050278e-19, 3.046778e-19, 3.038251e-19, 3.04414e-19, 3.041819e-19, 
    3.047342e-19, 3.050848e-19, 3.049115e-19, 3.059811e-19, 3.055654e-19, 
    3.077526e-19, 3.068113e-19, 3.092633e-19, 3.086773e-19, 3.094037e-19, 
    3.090332e-19, 3.096679e-19, 3.090967e-19, 3.100861e-19, 3.103013e-19, 
    3.101542e-19, 3.107193e-19, 3.090649e-19, 3.097006e-19, 3.049066e-19, 
    3.049348e-19, 3.050666e-19, 3.044871e-19, 3.044517e-19, 3.039205e-19, 
    3.043932e-19, 3.045944e-19, 3.051052e-19, 3.054071e-19, 3.056939e-19, 
    3.063243e-19, 3.070276e-19, 3.080101e-19, 3.087153e-19, 3.091876e-19, 
    3.08898e-19, 3.091537e-19, 3.088679e-19, 3.087339e-19, 3.102206e-19, 
    3.093861e-19, 3.10638e-19, 3.105688e-19, 3.100024e-19, 3.105766e-19, 
    3.049547e-19, 3.04792e-19, 3.042265e-19, 3.046691e-19, 3.038626e-19, 
    3.04314e-19, 3.045734e-19, 3.055739e-19, 3.057938e-19, 3.059973e-19, 
    3.063994e-19, 3.069149e-19, 3.078185e-19, 3.086037e-19, 3.093202e-19, 
    3.092677e-19, 3.092862e-19, 3.09446e-19, 3.090499e-19, 3.095111e-19, 
    3.095883e-19, 3.093861e-19, 3.105596e-19, 3.102245e-19, 3.105674e-19, 
    3.103492e-19, 3.048449e-19, 3.051187e-19, 3.049708e-19, 3.052489e-19, 
    3.050529e-19, 3.059239e-19, 3.061849e-19, 3.074051e-19, 3.069048e-19, 
    3.077011e-19, 3.069858e-19, 3.071125e-19, 3.077267e-19, 3.070245e-19, 
    3.085603e-19, 3.075191e-19, 3.094522e-19, 3.084134e-19, 3.095173e-19, 
    3.093171e-19, 3.096486e-19, 3.099454e-19, 3.103187e-19, 3.110068e-19, 
    3.108475e-19, 3.114227e-19, 3.055268e-19, 3.058816e-19, 3.058505e-19, 
    3.062217e-19, 3.064961e-19, 3.070907e-19, 3.080431e-19, 3.076852e-19, 
    3.083424e-19, 3.08474e-19, 3.074758e-19, 3.080888e-19, 3.06119e-19, 
    3.064375e-19, 3.06248e-19, 3.055547e-19, 3.077674e-19, 3.066326e-19, 
    3.087269e-19, 3.081132e-19, 3.09903e-19, 3.090132e-19, 3.107598e-19, 
    3.115048e-19, 3.12206e-19, 3.130237e-19, 3.060753e-19, 3.058343e-19, 
    3.062659e-19, 3.068623e-19, 3.074158e-19, 3.081507e-19, 3.082259e-19, 
    3.083634e-19, 3.087196e-19, 3.09019e-19, 3.084068e-19, 3.090941e-19, 
    3.06511e-19, 3.078659e-19, 3.05743e-19, 3.063827e-19, 3.068273e-19, 
    3.066324e-19, 3.076443e-19, 3.078825e-19, 3.088496e-19, 3.0835e-19, 
    3.113208e-19, 3.100078e-19, 3.136462e-19, 3.126311e-19, 3.0575e-19, 
    3.060746e-19, 3.072026e-19, 3.066661e-19, 3.081998e-19, 3.085766e-19, 
    3.08883e-19, 3.092744e-19, 3.093167e-19, 3.095485e-19, 3.091686e-19, 
    3.095335e-19, 3.081522e-19, 3.087697e-19, 3.070739e-19, 3.07487e-19, 
    3.072971e-19, 3.070885e-19, 3.077318e-19, 3.084162e-19, 3.084311e-19, 
    3.086504e-19, 3.092676e-19, 3.08206e-19, 3.114896e-19, 3.094629e-19, 
    3.064282e-19, 3.070522e-19, 3.071416e-19, 3.068999e-19, 3.085388e-19, 
    3.079455e-19, 3.095429e-19, 3.091115e-19, 3.098182e-19, 3.094671e-19, 
    3.094154e-19, 3.089642e-19, 3.086831e-19, 3.079726e-19, 3.07394e-19, 
    3.06935e-19, 3.070418e-19, 3.075459e-19, 3.084581e-19, 3.093204e-19, 
    3.091316e-19, 3.097645e-19, 3.080887e-19, 3.087916e-19, 3.085199e-19, 
    3.092283e-19, 3.076756e-19, 3.089972e-19, 3.073373e-19, 3.07483e-19, 
    3.079337e-19, 3.088391e-19, 3.090397e-19, 3.092534e-19, 3.091216e-19, 
    3.084813e-19, 3.083767e-19, 3.079228e-19, 3.077973e-19, 3.074513e-19, 
    3.071646e-19, 3.074265e-19, 3.077014e-19, 3.084817e-19, 3.091842e-19, 
    3.099495e-19, 3.101368e-19, 3.110291e-19, 3.103025e-19, 3.115008e-19, 
    3.104816e-19, 3.122454e-19, 3.090741e-19, 3.104521e-19, 3.079542e-19, 
    3.082238e-19, 3.087107e-19, 3.098272e-19, 3.09225e-19, 3.099294e-19, 
    3.083726e-19, 3.075632e-19, 3.073539e-19, 3.069629e-19, 3.073629e-19, 
    3.073304e-19, 3.077129e-19, 3.0759e-19, 3.085076e-19, 3.080149e-19, 
    3.09414e-19, 3.099239e-19, 3.113623e-19, 3.122426e-19, 3.131379e-19, 
    3.135327e-19, 3.136529e-19, 3.137031e-19 ;

 CWDN_vr =
  1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062149e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062149e-07, 1.062148e-07, 1.062149e-07, 1.062149e-07, 1.062148e-07, 
    1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 
    1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504 ;

 DEADSTEMN =
  6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05 ;

 DENIT =
  1.095659e-14, 1.099812e-14, 1.099e-14, 1.102352e-14, 1.10049e-14, 
    1.102682e-14, 1.096491e-14, 1.099965e-14, 1.097744e-14, 1.096016e-14, 
    1.108844e-14, 1.102487e-14, 1.115442e-14, 1.111384e-14, 1.121569e-14, 
    1.114807e-14, 1.12293e-14, 1.121367e-14, 1.126058e-14, 1.124711e-14, 
    1.130714e-14, 1.126674e-14, 1.133822e-14, 1.129745e-14, 1.130381e-14, 
    1.126532e-14, 1.103777e-14, 1.108067e-14, 1.10352e-14, 1.104132e-14, 
    1.103855e-14, 1.100521e-14, 1.098843e-14, 1.095324e-14, 1.095959e-14, 
    1.098542e-14, 1.104393e-14, 1.102402e-14, 1.107408e-14, 1.107296e-14, 
    1.11287e-14, 1.110355e-14, 1.119731e-14, 1.117062e-14, 1.124765e-14, 
    1.122825e-14, 1.124671e-14, 1.124108e-14, 1.124673e-14, 1.121832e-14, 
    1.123045e-14, 1.120545e-14, 1.110848e-14, 1.113707e-14, 1.105174e-14, 
    1.100046e-14, 1.096636e-14, 1.09422e-14, 1.094558e-14, 1.095209e-14, 
    1.098554e-14, 1.101696e-14, 1.104094e-14, 1.105695e-14, 1.107274e-14, 
    1.112065e-14, 1.114595e-14, 1.120267e-14, 1.11924e-14, 1.120974e-14, 
    1.12263e-14, 1.125411e-14, 1.124952e-14, 1.126176e-14, 1.120917e-14, 
    1.124411e-14, 1.11864e-14, 1.120218e-14, 1.107728e-14, 1.102947e-14, 
    1.10092e-14, 1.09914e-14, 1.094819e-14, 1.097802e-14, 1.096624e-14, 
    1.099417e-14, 1.101194e-14, 1.100312e-14, 1.105737e-14, 1.103625e-14, 
    1.114742e-14, 1.109952e-14, 1.122439e-14, 1.119447e-14, 1.12315e-14, 
    1.121259e-14, 1.124496e-14, 1.12158e-14, 1.126628e-14, 1.12773e-14, 
    1.126973e-14, 1.129861e-14, 1.121407e-14, 1.124653e-14, 1.100298e-14, 
    1.100442e-14, 1.101107e-14, 1.098169e-14, 1.097989e-14, 1.095295e-14, 
    1.097687e-14, 1.098707e-14, 1.101292e-14, 1.10282e-14, 1.104273e-14, 
    1.107475e-14, 1.111049e-14, 1.116047e-14, 1.119638e-14, 1.122044e-14, 
    1.120566e-14, 1.121868e-14, 1.120409e-14, 1.119723e-14, 1.127312e-14, 
    1.12305e-14, 1.129441e-14, 1.129087e-14, 1.126191e-14, 1.129122e-14, 
    1.100539e-14, 1.09971e-14, 1.096846e-14, 1.099084e-14, 1.094999e-14, 
    1.097285e-14, 1.098598e-14, 1.103667e-14, 1.104778e-14, 1.105813e-14, 
    1.107852e-14, 1.11047e-14, 1.115068e-14, 1.119067e-14, 1.122719e-14, 
    1.122448e-14, 1.122542e-14, 1.123355e-14, 1.121333e-14, 1.123684e-14, 
    1.124077e-14, 1.123044e-14, 1.129034e-14, 1.127322e-14, 1.129072e-14, 
    1.127954e-14, 1.099977e-14, 1.101362e-14, 1.10061e-14, 1.102021e-14, 
    1.101024e-14, 1.105445e-14, 1.106768e-14, 1.112969e-14, 1.110419e-14, 
    1.114472e-14, 1.110826e-14, 1.111472e-14, 1.114601e-14, 1.111018e-14, 
    1.118842e-14, 1.113536e-14, 1.123385e-14, 1.118088e-14, 1.123713e-14, 
    1.122688e-14, 1.124378e-14, 1.125895e-14, 1.127798e-14, 1.131319e-14, 
    1.1305e-14, 1.133444e-14, 1.10343e-14, 1.105229e-14, 1.105069e-14, 
    1.106951e-14, 1.108344e-14, 1.111366e-14, 1.116213e-14, 1.114386e-14, 
    1.117731e-14, 1.118404e-14, 1.113314e-14, 1.116438e-14, 1.106416e-14, 
    1.108033e-14, 1.107067e-14, 1.103545e-14, 1.114792e-14, 1.109017e-14, 
    1.119676e-14, 1.116545e-14, 1.125673e-14, 1.121133e-14, 1.13005e-14, 
    1.133867e-14, 1.137452e-14, 1.141648e-14, 1.10621e-14, 1.104983e-14, 
    1.107172e-14, 1.110207e-14, 1.113015e-14, 1.116758e-14, 1.117138e-14, 
    1.117836e-14, 1.119649e-14, 1.121177e-14, 1.118055e-14, 1.121555e-14, 
    1.108408e-14, 1.115292e-14, 1.104497e-14, 1.107748e-14, 1.110001e-14, 
    1.10901e-14, 1.114153e-14, 1.115364e-14, 1.120293e-14, 1.117743e-14, 
    1.13292e-14, 1.126203e-14, 1.144838e-14, 1.139629e-14, 1.104553e-14, 
    1.106197e-14, 1.111931e-14, 1.109202e-14, 1.117002e-14, 1.118924e-14, 
    1.120482e-14, 1.12248e-14, 1.122691e-14, 1.123875e-14, 1.121931e-14, 
    1.123794e-14, 1.116746e-14, 1.119894e-14, 1.111254e-14, 1.113353e-14, 
    1.112385e-14, 1.111321e-14, 1.114593e-14, 1.118083e-14, 1.118154e-14, 
    1.11927e-14, 1.122428e-14, 1.116999e-14, 1.133784e-14, 1.123416e-14, 
    1.107992e-14, 1.111165e-14, 1.111614e-14, 1.110385e-14, 1.118726e-14, 
    1.115702e-14, 1.123846e-14, 1.121641e-14, 1.125246e-14, 1.123454e-14, 
    1.123186e-14, 1.120884e-14, 1.119447e-14, 1.115827e-14, 1.112877e-14, 
    1.110541e-14, 1.11108e-14, 1.113647e-14, 1.118291e-14, 1.122688e-14, 
    1.121723e-14, 1.124949e-14, 1.116398e-14, 1.119984e-14, 1.118594e-14, 
    1.122206e-14, 1.11433e-14, 1.121075e-14, 1.112605e-14, 1.113344e-14, 
    1.115637e-14, 1.120256e-14, 1.121271e-14, 1.122363e-14, 1.121685e-14, 
    1.118422e-14, 1.117885e-14, 1.115569e-14, 1.114928e-14, 1.113166e-14, 
    1.111703e-14, 1.113037e-14, 1.114433e-14, 1.118409e-14, 1.12199e-14, 
    1.125894e-14, 1.126849e-14, 1.131416e-14, 1.127697e-14, 1.133833e-14, 
    1.128617e-14, 1.13764e-14, 1.121458e-14, 1.128498e-14, 1.115741e-14, 
    1.117112e-14, 1.119597e-14, 1.125293e-14, 1.122212e-14, 1.125812e-14, 
    1.117862e-14, 1.11374e-14, 1.112669e-14, 1.110681e-14, 1.112711e-14, 
    1.112546e-14, 1.11449e-14, 1.113862e-14, 1.118535e-14, 1.116024e-14, 
    1.123156e-14, 1.125761e-14, 1.133115e-14, 1.137623e-14, 1.142212e-14, 
    1.144236e-14, 1.144852e-14, 1.145108e-14 ;

 DISPVEGC =
  0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638 ;

 DISPVEGN =
  0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959 ;

 DSTDEP =
  2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  6.265611, 6.281866, 6.278709, 6.291808, 6.284558, 6.293118, 6.268916, 
    6.282502, 6.273832, 6.26709, 6.317191, 6.292393, 6.343135, 6.327245, 
    6.368863, 6.340642, 6.374258, 6.368121, 6.386682, 6.381361, 6.405095, 
    6.389139, 6.417484, 6.401298, 6.403816, 6.388608, 6.297404, 6.314094, 
    6.29641, 6.298789, 6.297728, 6.284698, 6.278101, 6.26439, 6.266882, 
    6.276964, 6.29986, 6.29211, 6.311711, 6.311269, 6.333107, 6.323251, 
    6.361673, 6.349604, 6.381584, 6.373917, 6.381218, 6.379007, 6.381247, 
    6.370008, 6.37482, 6.36495, 6.32509, 6.336307, 6.302886, 6.282793, 
    6.269506, 6.260073, 6.261406, 6.263942, 6.277022, 6.289359, 6.298735, 
    6.305011, 6.311204, 6.329888, 6.33986, 6.363783, 6.359766, 6.366591, 
    6.373156, 6.384159, 6.38235, 6.387197, 6.366429, 6.380215, 6.357474, 
    6.363681, 6.312795, 6.294204, 6.286236, 6.279312, 6.262429, 6.274078, 
    6.269481, 6.280444, 6.287403, 6.283966, 6.305183, 6.296926, 6.340452, 
    6.321678, 6.372391, 6.360592, 6.375226, 6.367758, 6.38055, 6.369037, 
    6.389009, 6.393355, 6.390383, 6.401843, 6.368396, 6.381208, 6.283864, 
    6.284425, 6.287047, 6.275526, 6.274827, 6.264317, 6.273676, 6.277659, 
    6.287813, 6.293785, 6.299474, 6.312002, 6.325984, 6.345616, 6.361355, 
    6.37087, 6.36504, 6.370186, 6.364429, 6.361739, 6.39172, 6.374858, 
    6.400193, 6.398791, 6.387308, 6.39895, 6.28482, 6.281592, 6.27037, 
    6.279151, 6.263175, 6.2721, 6.277231, 6.297079, 6.301461, 6.305498, 
    6.313498, 6.323755, 6.341783, 6.359107, 6.373543, 6.372486, 6.372857, 
    6.376076, 6.368091, 6.377389, 6.378941, 6.374868, 6.398603, 6.391815, 
    6.398762, 6.394343, 6.282644, 6.288075, 6.285141, 6.290648, 6.286765, 
    6.304023, 6.309205, 6.333508, 6.323547, 6.339433, 6.325166, 6.327686, 
    6.339911, 6.325943, 6.358218, 6.335775, 6.376202, 6.353668, 6.377515, 
    6.37348, 6.380172, 6.38616, 6.39372, 6.407664, 6.404436, 6.416132, 
    6.296162, 6.303191, 6.302589, 6.309965, 6.315416, 6.327261, 6.346286, 
    6.339132, 6.352293, 6.35651, 6.334949, 6.347193, 6.307912, 6.31423, 
    6.310483, 6.296706, 6.340755, 6.318112, 6.361587, 6.347693, 6.385303, 
    6.367332, 6.402656, 6.417765, 6.432111, 6.448807, 6.307049, 6.302268, 
    6.310848, 6.322688, 6.333742, 6.348441, 6.349956, 6.352709, 6.36145, 
    6.367473, 6.353561, 6.368986, 6.315658, 6.342732, 6.300444, 6.313138, 
    6.321997, 6.318128, 6.338319, 6.343081, 6.364046, 6.352445, 6.414015, 
    6.387398, 6.461617, 6.440776, 6.300593, 6.307041, 6.329478, 6.3188, 
    6.349432, 6.358568, 6.364738, 6.372606, 6.37347, 6.37814, 6.370487, 
    6.377845, 6.348471, 6.362453, 6.326931, 6.335165, 6.331382, 6.327222, 
    6.340068, 6.355327, 6.35565, 6.360044, 6.372386, 6.349557, 6.4174, 
    6.376336, 6.314074, 6.326466, 6.328273, 6.323462, 6.357808, 6.344333, 
    6.37803, 6.369335, 6.383596, 6.376503, 6.375459, 6.366369, 6.36071, 
    6.344872, 6.333306, 6.324163, 6.32629, 6.336339, 6.356173, 6.373535, 
    6.369722, 6.382512, 6.347205, 6.362882, 6.357416, 6.371686, 6.338935, 
    6.366953, 6.332185, 6.335094, 6.344097, 6.36382, 6.367889, 6.372183, 
    6.36954, 6.356643, 6.352971, 6.343886, 6.341365, 6.334463, 6.32874, 
    6.333961, 6.339443, 6.356661, 6.370788, 6.386241, 6.390039, 6.408074, 
    6.393346, 6.417623, 6.396911, 6.432839, 6.368534, 6.396369, 6.344517, 
    6.349916, 6.361244, 6.383744, 6.371618, 6.385817, 6.352891, 6.33667, 
    6.332516, 6.324713, 6.332695, 6.332047, 6.339691, 6.337235, 6.357182, 
    6.345731, 6.375424, 6.385712, 6.414893, 6.432829, 6.451191, 6.459296, 
    6.461768, 6.4628 ;

 EFLX_LH_TOT_R =
  6.265611, 6.281866, 6.278709, 6.291808, 6.284558, 6.293118, 6.268916, 
    6.282502, 6.273832, 6.26709, 6.317191, 6.292393, 6.343135, 6.327245, 
    6.368863, 6.340642, 6.374258, 6.368121, 6.386682, 6.381361, 6.405095, 
    6.389139, 6.417484, 6.401298, 6.403816, 6.388608, 6.297404, 6.314094, 
    6.29641, 6.298789, 6.297728, 6.284698, 6.278101, 6.26439, 6.266882, 
    6.276964, 6.29986, 6.29211, 6.311711, 6.311269, 6.333107, 6.323251, 
    6.361673, 6.349604, 6.381584, 6.373917, 6.381218, 6.379007, 6.381247, 
    6.370008, 6.37482, 6.36495, 6.32509, 6.336307, 6.302886, 6.282793, 
    6.269506, 6.260073, 6.261406, 6.263942, 6.277022, 6.289359, 6.298735, 
    6.305011, 6.311204, 6.329888, 6.33986, 6.363783, 6.359766, 6.366591, 
    6.373156, 6.384159, 6.38235, 6.387197, 6.366429, 6.380215, 6.357474, 
    6.363681, 6.312795, 6.294204, 6.286236, 6.279312, 6.262429, 6.274078, 
    6.269481, 6.280444, 6.287403, 6.283966, 6.305183, 6.296926, 6.340452, 
    6.321678, 6.372391, 6.360592, 6.375226, 6.367758, 6.38055, 6.369037, 
    6.389009, 6.393355, 6.390383, 6.401843, 6.368396, 6.381208, 6.283864, 
    6.284425, 6.287047, 6.275526, 6.274827, 6.264317, 6.273676, 6.277659, 
    6.287813, 6.293785, 6.299474, 6.312002, 6.325984, 6.345616, 6.361355, 
    6.37087, 6.36504, 6.370186, 6.364429, 6.361739, 6.39172, 6.374858, 
    6.400193, 6.398791, 6.387308, 6.39895, 6.28482, 6.281592, 6.27037, 
    6.279151, 6.263175, 6.2721, 6.277231, 6.297079, 6.301461, 6.305498, 
    6.313498, 6.323755, 6.341783, 6.359107, 6.373543, 6.372486, 6.372857, 
    6.376076, 6.368091, 6.377389, 6.378941, 6.374868, 6.398603, 6.391815, 
    6.398762, 6.394343, 6.282644, 6.288075, 6.285141, 6.290648, 6.286765, 
    6.304023, 6.309205, 6.333508, 6.323547, 6.339433, 6.325166, 6.327686, 
    6.339911, 6.325943, 6.358218, 6.335775, 6.376202, 6.353668, 6.377515, 
    6.37348, 6.380172, 6.38616, 6.39372, 6.407664, 6.404436, 6.416132, 
    6.296162, 6.303191, 6.302589, 6.309965, 6.315416, 6.327261, 6.346286, 
    6.339132, 6.352293, 6.35651, 6.334949, 6.347193, 6.307912, 6.31423, 
    6.310483, 6.296706, 6.340755, 6.318112, 6.361587, 6.347693, 6.385303, 
    6.367332, 6.402656, 6.417765, 6.432111, 6.448807, 6.307049, 6.302268, 
    6.310848, 6.322688, 6.333742, 6.348441, 6.349956, 6.352709, 6.36145, 
    6.367473, 6.353561, 6.368986, 6.315658, 6.342732, 6.300444, 6.313138, 
    6.321997, 6.318128, 6.338319, 6.343081, 6.364046, 6.352445, 6.414015, 
    6.387398, 6.461617, 6.440776, 6.300593, 6.307041, 6.329478, 6.3188, 
    6.349432, 6.358568, 6.364738, 6.372606, 6.37347, 6.37814, 6.370487, 
    6.377845, 6.348471, 6.362453, 6.326931, 6.335165, 6.331382, 6.327222, 
    6.340068, 6.355327, 6.35565, 6.360044, 6.372386, 6.349557, 6.4174, 
    6.376336, 6.314074, 6.326466, 6.328273, 6.323462, 6.357808, 6.344333, 
    6.37803, 6.369335, 6.383596, 6.376503, 6.375459, 6.366369, 6.36071, 
    6.344872, 6.333306, 6.324163, 6.32629, 6.336339, 6.356173, 6.373535, 
    6.369722, 6.382512, 6.347205, 6.362882, 6.357416, 6.371686, 6.338935, 
    6.366953, 6.332185, 6.335094, 6.344097, 6.36382, 6.367889, 6.372183, 
    6.36954, 6.356643, 6.352971, 6.343886, 6.341365, 6.334463, 6.32874, 
    6.333961, 6.339443, 6.356661, 6.370788, 6.386241, 6.390039, 6.408074, 
    6.393346, 6.417623, 6.396911, 6.432839, 6.368534, 6.396369, 6.344517, 
    6.349916, 6.361244, 6.383744, 6.371618, 6.385817, 6.352891, 6.33667, 
    6.332516, 6.324713, 6.332695, 6.332047, 6.339691, 6.337235, 6.357182, 
    6.345731, 6.375424, 6.385712, 6.414893, 6.432829, 6.451191, 6.459296, 
    6.461768, 6.4628 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122 ;

 ER =
  6.359163e-08, 6.387121e-08, 6.381686e-08, 6.404235e-08, 6.391726e-08, 
    6.406492e-08, 6.364831e-08, 6.388231e-08, 6.373293e-08, 6.36168e-08, 
    6.447997e-08, 6.405241e-08, 6.492405e-08, 6.465138e-08, 6.533632e-08, 
    6.488163e-08, 6.542801e-08, 6.53232e-08, 6.563863e-08, 6.554826e-08, 
    6.595173e-08, 6.568033e-08, 6.616087e-08, 6.588692e-08, 6.592978e-08, 
    6.567138e-08, 6.413845e-08, 6.442674e-08, 6.412137e-08, 6.416248e-08, 
    6.414403e-08, 6.391985e-08, 6.380688e-08, 6.357025e-08, 6.361321e-08, 
    6.3787e-08, 6.418097e-08, 6.404723e-08, 6.438426e-08, 6.437665e-08, 
    6.475187e-08, 6.458269e-08, 6.521333e-08, 6.503409e-08, 6.555204e-08, 
    6.542178e-08, 6.554592e-08, 6.550827e-08, 6.554641e-08, 6.535537e-08, 
    6.543722e-08, 6.526912e-08, 6.461438e-08, 6.480681e-08, 6.423289e-08, 
    6.38878e-08, 6.365858e-08, 6.349591e-08, 6.351891e-08, 6.356274e-08, 
    6.378801e-08, 6.399981e-08, 6.416121e-08, 6.426918e-08, 6.437556e-08, 
    6.469757e-08, 6.486799e-08, 6.524958e-08, 6.518071e-08, 6.529738e-08, 
    6.540882e-08, 6.559594e-08, 6.556514e-08, 6.564758e-08, 6.529429e-08, 
    6.552909e-08, 6.514148e-08, 6.52475e-08, 6.44045e-08, 6.40833e-08, 
    6.394681e-08, 6.38273e-08, 6.353659e-08, 6.373735e-08, 6.365821e-08, 
    6.384649e-08, 6.396612e-08, 6.390695e-08, 6.427213e-08, 6.413016e-08, 
    6.487809e-08, 6.455593e-08, 6.539582e-08, 6.519484e-08, 6.544399e-08, 
    6.531685e-08, 6.55347e-08, 6.533864e-08, 6.567826e-08, 6.575221e-08, 
    6.570168e-08, 6.58958e-08, 6.532778e-08, 6.554592e-08, 6.39053e-08, 
    6.391495e-08, 6.39599e-08, 6.376228e-08, 6.375019e-08, 6.356908e-08, 
    6.373023e-08, 6.379886e-08, 6.397305e-08, 6.40761e-08, 6.417405e-08, 
    6.438941e-08, 6.462994e-08, 6.496626e-08, 6.520787e-08, 6.536983e-08, 
    6.527052e-08, 6.53582e-08, 6.526018e-08, 6.521424e-08, 6.572451e-08, 
    6.543799e-08, 6.586788e-08, 6.584409e-08, 6.564954e-08, 6.584677e-08, 
    6.392172e-08, 6.386619e-08, 6.367338e-08, 6.382427e-08, 6.354936e-08, 
    6.370324e-08, 6.379173e-08, 6.413313e-08, 6.420814e-08, 6.427769e-08, 
    6.441505e-08, 6.459135e-08, 6.49006e-08, 6.516968e-08, 6.54153e-08, 
    6.539731e-08, 6.540364e-08, 6.545852e-08, 6.53226e-08, 6.548083e-08, 
    6.550739e-08, 6.543795e-08, 6.58409e-08, 6.572579e-08, 6.584358e-08, 
    6.576862e-08, 6.388424e-08, 6.397768e-08, 6.392719e-08, 6.402214e-08, 
    6.395525e-08, 6.425269e-08, 6.434187e-08, 6.475913e-08, 6.458788e-08, 
    6.486043e-08, 6.461556e-08, 6.465896e-08, 6.486933e-08, 6.462879e-08, 
    6.515485e-08, 6.479821e-08, 6.546065e-08, 6.510453e-08, 6.548296e-08, 
    6.541424e-08, 6.552803e-08, 6.562993e-08, 6.575814e-08, 6.59947e-08, 
    6.593991e-08, 6.613774e-08, 6.411698e-08, 6.423819e-08, 6.422751e-08, 
    6.435434e-08, 6.444814e-08, 6.465145e-08, 6.497752e-08, 6.485489e-08, 
    6.508e-08, 6.512519e-08, 6.47832e-08, 6.499319e-08, 6.431929e-08, 
    6.442818e-08, 6.436335e-08, 6.412655e-08, 6.488316e-08, 6.449487e-08, 
    6.521186e-08, 6.500152e-08, 6.56154e-08, 6.531011e-08, 6.590976e-08, 
    6.616612e-08, 6.640736e-08, 6.668932e-08, 6.430432e-08, 6.422197e-08, 
    6.436942e-08, 6.457343e-08, 6.476271e-08, 6.501435e-08, 6.504009e-08, 
    6.508724e-08, 6.520934e-08, 6.531201e-08, 6.510215e-08, 6.533775e-08, 
    6.445345e-08, 6.491686e-08, 6.419084e-08, 6.440948e-08, 6.456141e-08, 
    6.449476e-08, 6.484088e-08, 6.492246e-08, 6.525397e-08, 6.50826e-08, 
    6.610285e-08, 6.565147e-08, 6.690398e-08, 6.655396e-08, 6.41932e-08, 
    6.430404e-08, 6.46898e-08, 6.450625e-08, 6.503114e-08, 6.516034e-08, 
    6.526538e-08, 6.539964e-08, 6.541413e-08, 6.549368e-08, 6.536332e-08, 
    6.548853e-08, 6.501489e-08, 6.522654e-08, 6.46457e-08, 6.478708e-08, 
    6.472204e-08, 6.46507e-08, 6.487087e-08, 6.510545e-08, 6.511046e-08, 
    6.518567e-08, 6.539766e-08, 6.503327e-08, 6.616113e-08, 6.546461e-08, 
    6.44249e-08, 6.463841e-08, 6.466889e-08, 6.458619e-08, 6.514739e-08, 
    6.494405e-08, 6.549174e-08, 6.534372e-08, 6.558625e-08, 6.546573e-08, 
    6.5448e-08, 6.529321e-08, 6.519684e-08, 6.495338e-08, 6.475528e-08, 
    6.459818e-08, 6.463471e-08, 6.480727e-08, 6.51198e-08, 6.541545e-08, 
    6.535068e-08, 6.556781e-08, 6.499309e-08, 6.523408e-08, 6.514095e-08, 
    6.538381e-08, 6.485164e-08, 6.530484e-08, 6.47358e-08, 6.47857e-08, 
    6.494002e-08, 6.525044e-08, 6.53191e-08, 6.539243e-08, 6.534718e-08, 
    6.512773e-08, 6.509178e-08, 6.493626e-08, 6.489333e-08, 6.477483e-08, 
    6.467673e-08, 6.476636e-08, 6.486049e-08, 6.512782e-08, 6.536873e-08, 
    6.563138e-08, 6.569566e-08, 6.600256e-08, 6.575274e-08, 6.616501e-08, 
    6.581453e-08, 6.642122e-08, 6.533109e-08, 6.58042e-08, 6.494704e-08, 
    6.503938e-08, 6.520641e-08, 6.558949e-08, 6.538266e-08, 6.562454e-08, 
    6.509037e-08, 6.481324e-08, 6.474151e-08, 6.460773e-08, 6.474458e-08, 
    6.473344e-08, 6.486439e-08, 6.482231e-08, 6.51367e-08, 6.496782e-08, 
    6.544756e-08, 6.562262e-08, 6.611701e-08, 6.642009e-08, 6.672858e-08, 
    6.686479e-08, 6.690624e-08, 6.692357e-08 ;

 ERRH2O =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRH2OSNO =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRSEB =
  -1.476203e-14, -7.60264e-15, -4.508943e-15, -7.046479e-15, -9.455054e-15, 
    -5.95794e-15, -1.302894e-14, -1.280743e-14, -2.101688e-15, -2.45333e-15, 
    -1.077052e-14, -2.287377e-16, -1.569488e-14, -7.869937e-15, -2.04615e-14, 
    -9.59848e-16, -2.817901e-15, -1.059036e-14, -1.32837e-14, -1.170554e-14, 
    -1.519579e-14, -5.142135e-15, -1.294947e-14, -2.930562e-15, 
    -1.060642e-14, -1.118337e-14, -1.052144e-14, -1.982162e-14, 
    -1.253492e-14, -1.397486e-14, -9.813404e-15, -7.933848e-15, 
    -1.543418e-14, -8.606963e-15, -4.315236e-15, -4.312975e-15, 
    -1.042418e-14, -8.426359e-15, -9.669485e-15, -1.208619e-14, 
    -1.108093e-14, -1.700479e-14, -1.636519e-14, -9.9513e-15, -3.94989e-15, 
    -1.354375e-14, -9.220583e-15, -1.315678e-14, -9.252801e-15, 
    -9.592762e-15, -1.268669e-14, -6.629385e-15, -1.587693e-14, 
    -8.755405e-15, -1.445176e-14, -3.370445e-15, -1.605973e-14, -1.34778e-14, 
    -6.467685e-15, -8.549436e-15, -1.574129e-14, -1.669194e-14, 
    -9.282188e-15, -7.749831e-15, -5.778552e-15, -1.066358e-14, 
    -9.466417e-15, -1.169341e-14, -9.929201e-15, -2.47065e-14, -8.374489e-15, 
    -1.049117e-14, -3.964066e-15, -5.047961e-15, -6.368025e-15, 
    -6.500414e-15, -8.807652e-15, -1.264199e-14, -1.443026e-14, 
    -2.364615e-15, -1.362244e-14, -6.187751e-15, -1.130188e-14, 
    -5.761319e-15, 5.308633e-15, -1.322296e-14, -6.90569e-15, -6.828631e-15, 
    -2.58046e-15, -1.596893e-14, 2.666836e-16, -1.324927e-14, -4.040089e-15, 
    -2.662325e-15, -1.056436e-14, -2.342362e-15, -2.412495e-16, 
    -1.452481e-14, -1.45556e-14, -1.281945e-14, -6.541895e-15, -1.455385e-14, 
    -1.71244e-14, -1.169352e-14, -8.223158e-15, -1.814805e-14, -7.022676e-15, 
    -4.066442e-15, -5.895013e-15, -2.412766e-15, -1.522253e-14, 
    -7.877457e-15, -6.5227e-15, -1.01298e-14, -1.944756e-14, -7.056676e-15, 
    -1.525767e-14, -2.954596e-15, -1.278989e-14, -5.51168e-15, -1.138837e-14, 
    -7.474904e-15, -1.553483e-15, -1.512685e-14, -1.302716e-14, 
    -8.206519e-15, -3.495341e-15, -1.16083e-14, -1.349472e-14, -1.047129e-14, 
    -3.429051e-15, -1.100651e-14, -8.66716e-15, -1.546287e-14, -2.780052e-15, 
    -6.686934e-15, -1.383873e-14, -4.313127e-15, -7.883708e-15, 
    -4.364647e-15, -2.328804e-15, -3.181617e-15, -1.581227e-14, 
    -9.481181e-15, -2.500058e-15, -9.55685e-15, -7.668315e-15, -5.753648e-15, 
    -8.369442e-15, -7.410407e-15, -2.648701e-15, -4.551011e-15, -1.95549e-14, 
    -6.495759e-15, -6.071027e-15, -4.282038e-15, -1.530475e-14, 
    -1.301373e-14, -4.270038e-15, -5.267672e-15, -1.498496e-14, 6.078484e-16, 
    -1.008893e-14, -8.976331e-15, -3.485216e-15, -2.197358e-14, 
    -9.835979e-15, -1.398294e-14, -4.7994e-15, -2.84633e-15, -3.879795e-15, 
    -9.663793e-15, -1.164176e-14, -4.796612e-15, -1.08445e-14, -1.021733e-14, 
    -1.789525e-14, -9.511677e-15, -4.97499e-15, -1.639865e-14, -9.759618e-15, 
    -1.277784e-14, -8.298883e-15, 4.663925e-15, -1.282956e-14, -8.566645e-15, 
    -1.138672e-14, -2.031125e-14, -1.092832e-14, -5.149656e-15, 
    -7.944152e-15, -8.394101e-15, -1.232341e-14, -3.723341e-15, 
    -1.072339e-15, -5.687067e-16, -9.6556e-15, -1.518992e-14, -6.445346e-15, 
    -1.216626e-14, -8.986129e-15, -1.16162e-14, -1.62073e-14, -1.446825e-14, 
    -1.374157e-14, -1.622786e-14, -1.29448e-14, -1.027706e-14, -1.295729e-14, 
    -1.224584e-14, -1.249781e-14, -1.042851e-14, -1.920957e-15, 
    -9.853677e-15, -6.737431e-15, -1.320809e-14, -1.571768e-14, -5.53656e-15, 
    -1.11142e-14, -1.529545e-14, -1.476977e-14, 9.659312e-16, -1.193016e-14, 
    -1.370455e-14, -8.56509e-15, -1.039778e-14, -1.447408e-14, -5.126342e-15, 
    -3.956087e-16, -5.019558e-15, -5.566155e-15, -8.359704e-15, 
    -2.554776e-15, -2.03837e-14, -3.240762e-15, -5.838757e-15, -8.012697e-15, 
    -1.451451e-14, -1.512276e-14, -1.914856e-14, -1.038014e-14, -1.1314e-14, 
    -1.283761e-14, -4.635811e-15, -8.746527e-15, -1.007215e-14, 
    -1.272753e-14, -1.424952e-14, -1.0505e-14, -1.466772e-15, -1.188315e-14, 
    -1.172464e-14, -1.691998e-14, -1.236655e-14, -9.772671e-15, -5.86797e-15, 
    -1.190921e-14, -2.349252e-15, 2.521281e-15, -7.899152e-15, -4.603405e-15, 
    -1.953087e-14, -8.165722e-15, -1.348104e-14, -1.653103e-14, 
    -1.487592e-14, -1.649581e-14, -1.231488e-14, -6.902886e-15, 
    -1.041371e-14, -7.635102e-15, -1.010894e-14, -2.248865e-15, 
    -1.637269e-14, -8.40505e-15, -8.83018e-15, -1.038409e-14, -1.26429e-14, 
    -6.68294e-15, -1.051764e-14, -1.691491e-14, -7.681307e-15, -7.13001e-15, 
    -1.185778e-14, -9.179095e-15, -3.51248e-15, -1.115295e-14, -7.029189e-15, 
    -1.326793e-14, -1.309435e-14, -6.280539e-15, -8.386431e-15, 
    -7.350658e-15, -5.110151e-15, -1.444781e-14, -1.51312e-14, -1.388162e-14, 
    -1.496585e-15, -5.544231e-15, -1.319142e-14, -1.181213e-14, 
    -9.771641e-15, -1.317383e-14, -3.379814e-15, -6.543355e-15, 
    -1.018473e-14, -1.958283e-14, -5.890755e-15, -8.883766e-15, 1.497526e-15, 
    -8.126374e-15, -1.29636e-14, -1.803747e-15, -1.100874e-14, -6.350786e-15, 
    1.647544e-15, -1.668759e-14, -7.382958e-15, -1.07461e-14, -5.564539e-15, 
    -9.106556e-15, -8.36322e-15, -6.197511e-15, -8.909165e-15, -2.620719e-14, 
    -7.677567e-15, 1.139544e-15, -1.173185e-14, 1.743273e-15, -2.074917e-14, 
    -1.418557e-14, -4.986783e-15, -8.432015e-15, -1.147529e-14, -6.29539e-15, 
    -1.585613e-14, -7.69955e-15, -1.021103e-14 ;

 ERRSOI =
  -71.2503, -71.34345, -71.32575, -71.40002, -71.35948, -71.40762, -71.26998, 
    -71.34644, -71.29809, -71.25979, -71.54214, -71.40353, -71.69436, 
    -71.60431, -71.8334, -71.67923, -71.86488, -71.8308, -71.93796, 
    -71.90735, -72.0408, -71.95211, -72.1132, -72.0206, -72.03437, -71.94888, 
    -71.43314, -71.52427, -71.42734, -71.44042, -71.43497, -71.35968, 
    -71.32061, -71.24444, -71.25859, -71.31523, -71.44634, -71.40299, 
    -71.5159, -71.51339, -71.63821, -71.58185, -71.7937, -71.73373, 
    -71.90866, -71.86433, -71.90626, -71.89378, -71.90642, -71.84154, 
    -71.86922, -71.81277, -71.59206, -71.6562, -71.46423, -71.34647, -71.273, 
    -71.21956, -71.2271, -71.24113, -71.31552, -71.38718, -71.44131, 
    -71.47727, -71.513, -71.61656, -71.67552, -71.80493, -71.78312, 
    -71.82127, -71.86001, -71.92299, -71.91285, -71.94025, -71.82141, 
    -71.89978, -71.77034, -71.8055, -71.51647, -71.41497, -71.36655, 
    -71.32893, -71.23278, -71.29882, -71.27263, -71.33627, -71.37586, 
    -71.35654, -71.47827, -71.43066, -71.67902, -71.5719, -71.85551, 
    -71.78773, -71.87199, -71.82928, -71.90197, -71.83656, -71.95095, 
    -71.97518, -71.95848, -72.0248, -71.83276, -71.90565, -71.3557, 
    -71.35881, -71.37406, -71.30698, -71.30325, -71.24374, -71.29725, 
    -71.31953, -71.37865, -71.41249, -71.44511, -71.517, -71.59639, 
    -71.70951, -71.79205, -71.84713, -71.81375, -71.84317, -71.81005, 
    -71.79482, -71.96569, -71.8691, -72.01524, -72.00735, -71.94064, 
    -72.00826, -71.36111, -71.34299, -71.27814, -71.3289, -71.23735, 
    -71.28778, -71.31635, -71.4303, -71.45686, -71.47957, -71.52591, 
    -71.5847, -71.68764, -71.77856, -71.86253, -71.8565, -71.85856, 
    -71.87669, -71.83092, -71.88427, -71.89263, -71.86983, -72.00626, 
    -71.96732, -72.00719, -71.98197, -71.34904, -71.37982, -71.36308, 
    -71.39422, -71.37178, -71.46984, -71.49925, -71.63907, -71.58318, 
    -71.67388, -71.59289, -71.60687, -71.67419, -71.59766, -71.77234, 
    -71.65144, -71.87742, -71.75383, -71.88501, -71.86215, -71.90063, 
    -71.93443, -71.97816, -72.05716, -72.0391, -72.10629, -71.42633, 
    -71.46577, -71.46346, -71.50561, -71.53653, -71.60515, -71.71404, 
    -71.67343, -71.74931, -71.76425, -71.64959, -71.71877, -71.49308, 
    -71.52823, -71.50817, -71.42875, -71.68117, -71.5507, -71.79319, 
    -71.7224, -71.92945, -71.82516, -72.02889, -72.11324, -72.19831, 
    -72.29153, -71.48859, -71.46164, -71.51096, -71.57713, -71.64198, 
    -71.72649, -71.7358, -71.7513, -71.79307, -71.82755, -71.75507, 
    -71.83632, -71.53402, -71.69306, -71.45036, -71.52171, -71.57375, 
    -71.5521, -71.66909, -71.6963, -71.80673, -71.75023, -72.09137, 
    -71.93991, -72.36665, -72.24611, -71.45194, -71.48905, -71.61676, 
    -71.55613, -71.73277, -71.77595, -71.81203, -71.85627, -71.86192, 
    -71.88832, -71.84493, -71.88706, -71.72666, -71.79849, -71.60355, 
    -71.65018, -71.62914, -71.60517, -71.67901, -71.75602, -71.75956, 
    -71.78392, -71.8493, -71.73351, -72.10746, -71.87281, -71.52943, 
    -71.5985, -71.61066, -71.58349, -71.77156, -71.703, -71.88795, -71.83829, 
    -71.92017, -71.8793, -71.8732, -71.82122, -71.78838, -71.70576, 
    -71.63932, -71.58766, -71.59981, -71.65662, -71.76116, -71.86159, 
    -71.83929, -71.91397, -71.71986, -71.8002, -71.76854, -71.85149, 
    -71.67192, -71.81906, -71.63377, -71.65038, -71.70165, -71.80438, 
    -71.82994, -71.85384, -71.83949, -71.76417, -71.75259, -71.70087, 
    -71.68567, -71.6469, -71.61394, -71.64359, -71.67433, -71.76499, 
    -71.84572, -71.93463, -71.95715, -72.05659, -71.973, -72.10838, 
    -71.98929, -72.19766, -71.83038, -71.98967, -71.70463, -71.73568, 
    -71.78996, -71.91867, -71.85113, -71.93105, -71.7523, -71.65763, 
    -71.63554, -71.59045, -71.63657, -71.6329, -71.67696, -71.6629, 
    -71.76803, -71.71155, -71.87253, -71.93089, -72.09855, -72.20051, 
    -72.30766, -72.35403, -72.36834, -72.3742 ;

 ERRSOL =
  4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18 ;

 ESAI =
  0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  -1.949492, -1.948384, -1.948594, -1.94771, -1.948192, -1.947619, -1.949257, 
    -1.948349, -1.948923, -1.949378, -1.946017, -1.947668, -1.944213, 
    -1.945278, -1.942567, -1.944392, -1.942192, -1.942597, -1.941318, 
    -1.941684, -1.940089, -1.941149, -1.939219, -1.94033, -1.940166, 
    -1.941188, -1.947314, -1.946229, -1.947384, -1.947228, -1.947292, 
    -1.94819, -1.948657, -1.94956, -1.949392, -1.94872, -1.947157, -1.947674, 
    -1.946325, -1.946355, -1.944877, -1.945544, -1.943039, -1.943744, 
    -1.941668, -1.942197, -1.941697, -1.941846, -1.941695, -1.942469, 
    -1.942139, -1.942812, -1.945423, -1.944664, -1.946943, -1.948349, 
    -1.949222, -1.949856, -1.949766, -1.9496, -1.948716, -1.947862, 
    -1.947216, -1.946787, -1.946359, -1.945135, -1.944436, -1.942906, 
    -1.943164, -1.942711, -1.942249, -1.941498, -1.941619, -1.941292, 
    -1.942709, -1.941775, -1.943316, -1.942898, -1.946321, -1.947531, 
    -1.94811, -1.948557, -1.949699, -1.948915, -1.949226, -1.948469, 
    -1.947997, -1.948227, -1.946775, -1.947344, -1.944394, -1.945662, 
    -1.942303, -1.94311, -1.942106, -1.942615, -1.941749, -1.942528, 
    -1.941163, -1.940874, -1.941073, -1.940279, -1.942574, -1.941705, 
    -1.948237, -1.9482, -1.948018, -1.948818, -1.948862, -1.949569, 
    -1.948933, -1.948668, -1.947963, -1.94756, -1.947171, -1.946312, 
    -1.945373, -1.944033, -1.943058, -1.942402, -1.9428, -1.94245, -1.942844, 
    -1.943025, -1.940988, -1.942141, -1.940394, -1.940488, -1.941287, 
    -1.940477, -1.948173, -1.948388, -1.94916, -1.948556, -1.949645, 
    -1.949046, -1.948707, -1.947349, -1.947031, -1.94676, -1.946206, 
    -1.94551, -1.944291, -1.943219, -1.942219, -1.942291, -1.942266, 
    -1.94205, -1.942596, -1.94196, -1.94186, -1.942132, -1.940501, -1.940967, 
    -1.94049, -1.940792, -1.948316, -1.94795, -1.948149, -1.947779, 
    -1.948046, -1.946877, -1.946525, -1.944868, -1.945528, -1.944455, 
    -1.945413, -1.945248, -1.944453, -1.945356, -1.943294, -1.944722, 
    -1.942042, -1.943508, -1.941951, -1.942223, -1.941764, -1.941361, 
    -1.940838, -1.939891, -1.940108, -1.939301, -1.947395, -1.946925, 
    -1.946952, -1.946448, -1.94608, -1.945268, -1.943978, -1.944459, 
    -1.943559, -1.943389, -1.944741, -1.943923, -1.946598, -1.94618, 
    -1.946417, -1.947367, -1.944368, -1.945913, -1.943045, -1.943879, 
    -1.94142, -1.942665, -1.94023, -1.939219, -1.938193, -1.937068, 
    -1.946652, -1.946973, -1.946384, -1.945601, -1.944832, -1.943831, 
    -1.94372, -1.943536, -1.943046, -1.942636, -1.943492, -1.942531, 
    -1.946113, -1.944227, -1.947109, -1.946257, -1.94564, -1.945896, 
    -1.94451, -1.944188, -1.942884, -1.943548, -1.939482, -1.941297, 
    -1.936157, -1.937617, -1.947089, -1.946646, -1.945131, -1.945848, 
    -1.943756, -1.94325, -1.94282, -1.942294, -1.942226, -1.941912, 
    -1.942428, -1.941926, -1.943829, -1.942981, -1.945287, -1.944735, 
    -1.944984, -1.945268, -1.944393, -1.943488, -1.943444, -1.943155, 
    -1.942381, -1.943747, -1.939291, -1.9421, -1.946164, -1.945348, 
    -1.945203, -1.945524, -1.943302, -1.944109, -1.941916, -1.942508, 
    -1.941531, -1.942019, -1.942092, -1.942711, -1.943102, -1.944077, 
    -1.944864, -1.945475, -1.945331, -1.944659, -1.943426, -1.942231, 
    -1.942497, -1.941605, -1.943909, -1.942962, -1.943338, -1.942351, 
    -1.944477, -1.942741, -1.944929, -1.944732, -1.944125, -1.942913, 
    -1.942607, -1.942323, -1.942493, -1.94339, -1.943521, -1.944134, 
    -1.944314, -1.944773, -1.945164, -1.944813, -1.944449, -1.94338, 
    -1.94242, -1.941359, -1.941089, -1.9399, -1.940902, -1.93928, -1.940709, 
    -1.938204, -1.942604, -1.940703, -1.944089, -1.943721, -1.943084, 
    -1.941551, -1.942355, -1.941402, -1.943524, -1.944647, -1.944908, 
    -1.945442, -1.944896, -1.944939, -1.944417, -1.944584, -1.943344, 
    -1.944007, -1.9421, -1.941404, -1.939394, -1.938167, -1.936871, -1.93631, 
    -1.936136, -1.936065 ;

 FCH4 =
  1.670047e-13, 1.654605e-13, 1.65762e-13, 1.64507e-13, 1.652045e-13, 
    1.643808e-13, 1.66693e-13, 1.653989e-13, 1.662264e-13, 1.668664e-13, 
    1.620408e-13, 1.644507e-13, 1.585915e-13, 1.6001e-13, 1.563955e-13, 
    1.58814e-13, 1.558989e-13, 1.564663e-13, 1.547469e-13, 1.55243e-13, 
    1.530064e-13, 1.545169e-13, 1.518254e-13, 1.533694e-13, 1.531295e-13, 
    1.545664e-13, 1.639688e-13, 1.623429e-13, 1.640646e-13, 1.63834e-13, 
    1.639375e-13, 1.651902e-13, 1.658174e-13, 1.67122e-13, 1.66886e-13, 
    1.659274e-13, 1.637301e-13, 1.644797e-13, 1.625834e-13, 1.626265e-13, 
    1.594904e-13, 1.60363e-13, 1.57057e-13, 1.580113e-13, 1.552224e-13, 
    1.559327e-13, 1.552559e-13, 1.554617e-13, 1.552532e-13, 1.562925e-13, 
    1.558488e-13, 1.567576e-13, 1.602004e-13, 1.592047e-13, 1.634381e-13, 
    1.653684e-13, 1.666365e-13, 1.675294e-13, 1.674036e-13, 1.671632e-13, 
    1.659218e-13, 1.647445e-13, 1.63841e-13, 1.632336e-13, 1.626327e-13, 
    1.597717e-13, 1.588854e-13, 1.568626e-13, 1.572315e-13, 1.566056e-13, 
    1.56003e-13, 1.549816e-13, 1.551506e-13, 1.546976e-13, 1.566221e-13, 
    1.55348e-13, 1.574409e-13, 1.568738e-13, 1.62469e-13, 1.642778e-13, 
    1.650402e-13, 1.657041e-13, 1.673067e-13, 1.662019e-13, 1.666385e-13, 
    1.655977e-13, 1.649324e-13, 1.652618e-13, 1.632169e-13, 1.640153e-13, 
    1.588325e-13, 1.605001e-13, 1.560735e-13, 1.571559e-13, 1.55812e-13, 
    1.565005e-13, 1.553173e-13, 1.563829e-13, 1.545284e-13, 1.541193e-13, 
    1.543991e-13, 1.533196e-13, 1.564416e-13, 1.552559e-13, 1.652711e-13, 
    1.652174e-13, 1.649671e-13, 1.660641e-13, 1.66131e-13, 1.671285e-13, 
    1.662412e-13, 1.658617e-13, 1.648938e-13, 1.643182e-13, 1.637689e-13, 
    1.625543e-13, 1.601204e-13, 1.583695e-13, 1.570862e-13, 1.562143e-13, 
    1.5675e-13, 1.562772e-13, 1.568056e-13, 1.570521e-13, 1.542728e-13, 
    1.558447e-13, 1.534757e-13, 1.536084e-13, 1.546868e-13, 1.535935e-13, 
    1.651797e-13, 1.654884e-13, 1.665549e-13, 1.657209e-13, 1.672367e-13, 
    1.663902e-13, 1.659012e-13, 1.639987e-13, 1.635773e-13, 1.631856e-13, 
    1.62409e-13, 1.603186e-13, 1.587145e-13, 1.572905e-13, 1.559678e-13, 
    1.560655e-13, 1.560311e-13, 1.55733e-13, 1.564696e-13, 1.556114e-13, 
    1.554665e-13, 1.558448e-13, 1.536262e-13, 1.542657e-13, 1.536112e-13, 
    1.540282e-13, 1.653881e-13, 1.64868e-13, 1.651493e-13, 1.646199e-13, 
    1.64993e-13, 1.633266e-13, 1.628233e-13, 1.594527e-13, 1.603364e-13, 
    1.589249e-13, 1.601942e-13, 1.599709e-13, 1.588784e-13, 1.601262e-13, 
    1.573697e-13, 1.592496e-13, 1.557214e-13, 1.576378e-13, 1.555998e-13, 
    1.559736e-13, 1.553537e-13, 1.547948e-13, 1.540864e-13, 1.527649e-13, 
    1.530726e-13, 1.519567e-13, 1.640892e-13, 1.634083e-13, 1.634683e-13, 
    1.627527e-13, 1.622213e-13, 1.600096e-13, 1.583101e-13, 1.589537e-13, 
    1.577679e-13, 1.575277e-13, 1.593275e-13, 1.582275e-13, 1.629508e-13, 
    1.623347e-13, 1.627018e-13, 1.640356e-13, 1.588059e-13, 1.61956e-13, 
    1.570648e-13, 1.581835e-13, 1.548747e-13, 1.565369e-13, 1.532415e-13, 
    1.517957e-13, 1.504155e-13, 1.487801e-13, 1.630353e-13, 1.634995e-13, 
    1.626674e-13, 1.604105e-13, 1.594341e-13, 1.581157e-13, 1.579795e-13, 
    1.577295e-13, 1.570783e-13, 1.565266e-13, 1.576503e-13, 1.563877e-13, 
    1.621914e-13, 1.586292e-13, 1.636746e-13, 1.624407e-13, 1.604721e-13, 
    1.619566e-13, 1.590269e-13, 1.585998e-13, 1.56839e-13, 1.577541e-13, 
    1.521545e-13, 1.546763e-13, 1.475192e-13, 1.495682e-13, 1.636613e-13, 
    1.630369e-13, 1.598118e-13, 1.618912e-13, 1.580269e-13, 1.573403e-13, 
    1.567777e-13, 1.560529e-13, 1.559742e-13, 1.555414e-13, 1.562495e-13, 
    1.555694e-13, 1.581129e-13, 1.569861e-13, 1.600392e-13, 1.593074e-13, 
    1.596449e-13, 1.600134e-13, 1.588702e-13, 1.576328e-13, 1.576061e-13, 
    1.57205e-13, 1.560639e-13, 1.580156e-13, 1.518242e-13, 1.557001e-13, 
    1.623531e-13, 1.600768e-13, 1.599197e-13, 1.60345e-13, 1.574094e-13, 
    1.584863e-13, 1.555519e-13, 1.563555e-13, 1.550348e-13, 1.556937e-13, 
    1.557902e-13, 1.566279e-13, 1.571452e-13, 1.584373e-13, 1.594727e-13, 
    1.602835e-13, 1.600958e-13, 1.592023e-13, 1.575564e-13, 1.559671e-13, 
    1.563179e-13, 1.551359e-13, 1.58228e-13, 1.569457e-13, 1.574438e-13, 
    1.561386e-13, 1.589708e-13, 1.565656e-13, 1.595736e-13, 1.593146e-13, 
    1.585075e-13, 1.56858e-13, 1.564884e-13, 1.560919e-13, 1.563368e-13, 
    1.575142e-13, 1.577054e-13, 1.585272e-13, 1.587526e-13, 1.593711e-13, 
    1.598792e-13, 1.594151e-13, 1.589245e-13, 1.575137e-13, 1.562203e-13, 
    1.547868e-13, 1.544323e-13, 1.527207e-13, 1.541165e-13, 1.518022e-13, 
    1.537735e-13, 1.503359e-13, 1.564239e-13, 1.538308e-13, 1.584706e-13, 
    1.579833e-13, 1.570941e-13, 1.550172e-13, 1.561448e-13, 1.548245e-13, 
    1.577129e-13, 1.591713e-13, 1.59544e-13, 1.602345e-13, 1.595282e-13, 
    1.595858e-13, 1.589041e-13, 1.591239e-13, 1.574664e-13, 1.583612e-13, 
    1.557926e-13, 1.54835e-13, 1.520742e-13, 1.503423e-13, 1.485503e-13, 
    1.477504e-13, 1.475059e-13, 1.474035e-13 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  8.215103, 8.23025, 8.227304, 8.239517, 8.232751, 8.240738, 8.218173, 
    8.23085, 8.222755, 8.216468, 8.263208, 8.240061, 8.287348, 8.272523, 
    8.31143, 8.285034, 8.31645, 8.310719, 8.328, 8.323045, 8.345184, 
    8.330288, 8.356703, 8.341627, 8.343981, 8.329796, 8.244718, 8.260323, 
    8.243793, 8.246017, 8.24502, 8.232889, 8.226757, 8.21395, 8.216274, 
    8.225683, 8.247017, 8.239784, 8.258036, 8.257624, 8.277985, 8.268795, 
    8.304711, 8.293348, 8.323252, 8.316114, 8.322915, 8.320853, 8.322942, 
    8.312478, 8.316959, 8.307761, 8.270514, 8.280972, 8.249829, 8.231142, 
    8.218728, 8.209929, 8.211172, 8.213542, 8.225739, 8.237221, 8.245952, 
    8.251798, 8.257564, 8.275023, 8.284295, 8.306689, 8.302931, 8.309302, 
    8.315405, 8.325657, 8.323969, 8.328488, 8.309138, 8.32199, 8.30079, 
    8.30658, 8.259116, 8.241735, 8.234345, 8.227869, 8.212128, 8.222994, 
    8.218707, 8.228912, 8.2354, 8.232193, 8.251958, 8.24427, 8.284846, 
    8.26734, 8.314693, 8.303702, 8.317332, 8.310373, 8.322298, 8.311565, 
    8.330173, 8.334229, 8.331456, 8.342121, 8.31097, 8.322913, 8.232101, 
    8.232625, 8.235065, 8.224343, 8.22369, 8.213885, 8.22261, 8.226327, 
    8.235776, 8.241345, 8.246645, 8.258314, 8.271356, 8.289649, 8.304414, 
    8.313272, 8.307839, 8.312635, 8.307274, 8.304764, 8.332707, 8.316999, 
    8.340586, 8.339279, 8.328594, 8.339427, 8.232993, 8.229981, 8.21953, 
    8.227708, 8.212819, 8.221147, 8.225938, 8.244428, 8.248491, 8.252257, 
    8.259704, 8.269265, 8.286075, 8.302325, 8.315762, 8.314776, 8.315123, 
    8.318127, 8.310686, 8.319349, 8.320802, 8.317, 8.339105, 8.332782, 
    8.339252, 8.335135, 8.230961, 8.236025, 8.23329, 8.238427, 8.234811, 
    8.250899, 8.25573, 8.278376, 8.269075, 8.283887, 8.270579, 8.272935, 
    8.284363, 8.271299, 8.301511, 8.280498, 8.318244, 8.297175, 8.319466, 
    8.315703, 8.321936, 8.327521, 8.334558, 8.347555, 8.344543, 8.355433, 
    8.243557, 8.250115, 8.24954, 8.256413, 8.261497, 8.27253, 8.290264, 
    8.28359, 8.295852, 8.299898, 8.279691, 8.291116, 8.254511, 8.260409, 
    8.2569, 8.244072, 8.285124, 8.264026, 8.304631, 8.291573, 8.326724, 
    8.309998, 8.342886, 8.356984, 8.370303, 8.385876, 8.253701, 8.249241, 
    8.257232, 8.268289, 8.278574, 8.292272, 8.293676, 8.296245, 8.304496, 
    8.310108, 8.297053, 8.311517, 8.261771, 8.28696, 8.247553, 8.259395, 
    8.267637, 8.264024, 8.282829, 8.287269, 8.30693, 8.295994, 8.353498, 
    8.328694, 8.397775, 8.378393, 8.247683, 8.253687, 8.27461, 8.264648, 
    8.293188, 8.301818, 8.307558, 8.3149, 8.315697, 8.320051, 8.312916, 
    8.319772, 8.2923, 8.305435, 8.272218, 8.2799, 8.276366, 8.27249, 
    8.284461, 8.298814, 8.299094, 8.303199, 8.314768, 8.293303, 8.35669, 
    8.318436, 8.260238, 8.271814, 8.273476, 8.268986, 8.30111, 8.288442, 
    8.319946, 8.311843, 8.325128, 8.318521, 8.317551, 8.30908, 8.303812, 
    8.288949, 8.27817, 8.269637, 8.271621, 8.280997, 8.299599, 8.315765, 
    8.312219, 8.324117, 8.291114, 8.305843, 8.300755, 8.314036, 8.283412, 
    8.309693, 8.277114, 8.279826, 8.288222, 8.306733, 8.310496, 8.314507, 
    8.312033, 8.300034, 8.296492, 8.28802, 8.28568, 8.279236, 8.273904, 
    8.278774, 8.283892, 8.300041, 8.313208, 8.3276, 8.331128, 8.347974, 
    8.334248, 8.356902, 8.337621, 8.371043, 8.311138, 8.33707, 8.288607, 
    8.293637, 8.304328, 8.325294, 8.313973, 8.327219, 8.296415, 8.281318, 
    8.277425, 8.270155, 8.277591, 8.276986, 8.284108, 8.281819, 8.300526, 
    8.289739, 8.317524, 8.327115, 8.354287, 8.370996, 8.388062, 8.395606, 
    8.397904, 8.398865 ;

 FGR =
  -325.1869, -325.9453, -325.7983, -326.409, -326.0709, -326.4702, -325.3414, 
    -325.9747, -325.5709, -325.2563, -327.5912, -326.4364, -328.7964, 
    -328.0598, -329.9227, -328.6807, -330.1715, -329.889, -330.7437, 
    -330.499, -331.5886, -330.8567, -332.1565, -331.4148, -331.5301, 
    -330.8323, -326.6706, -327.4471, -326.6241, -326.735, -326.6857, 
    -326.0773, -325.7694, -325.1302, -325.2466, -325.7167, -326.7849, 
    -326.4235, -327.3378, -327.3172, -328.332, -327.8745, -329.5914, 
    -329.0965, -330.5092, -330.1562, -330.4923, -330.3906, -330.4936, 
    -329.976, -330.1977, -329.7427, -327.9598, -328.4803, -326.9262, 
    -325.9878, -325.3689, -324.9284, -324.9907, -325.109, -325.7194, 
    -326.295, -326.7328, -327.0255, -327.3142, -328.1817, -328.6447, 
    -329.6886, -329.5035, -329.8182, -330.1211, -330.6276, -330.5445, 
    -330.7672, -329.811, -330.446, -329.3977, -329.6842, -327.3865, 
    -326.5213, -326.1483, -325.8263, -325.0384, -325.5822, -325.3676, 
    -325.8793, -326.2036, -326.0435, -327.0335, -326.6484, -328.6721, 
    -327.8011, -330.0858, -329.5416, -330.2165, -329.8724, -330.4615, 
    -329.9313, -330.8506, -331.0502, -330.9137, -331.44, -329.9018, 
    -330.4917, -326.0387, -326.0648, -326.187, -325.6497, -325.6171, 
    -325.1267, -325.5637, -325.7492, -326.2228, -326.5017, -326.7672, 
    -327.3511, -328.0011, -328.9115, -329.5768, -330.0158, -329.747, 
    -329.9843, -329.7188, -329.5947, -330.975, -330.1994, -331.3643, -331.3, 
    -330.7723, -331.3073, -326.0832, -325.9329, -325.4093, -325.8191, 
    -325.0734, -325.49, -325.7291, -326.6551, -326.86, -327.0481, -327.4209, 
    -327.8979, -328.7341, -329.4728, -330.139, -330.0903, -330.1074, 
    -330.2556, -329.8876, -330.3161, -330.3874, -330.2, -331.2914, -330.9796, 
    -331.2986, -331.0958, -325.9819, -326.235, -326.0981, -326.3551, 
    -326.1736, -326.9789, -327.2203, -328.3501, -327.8882, -328.6251, 
    -327.9635, -328.0804, -328.6466, -327.9996, -329.4315, -328.4552, 
    -330.2614, -329.2836, -330.3219, -330.1361, -330.4443, -330.7196, 
    -331.0671, -331.7067, -331.5589, -332.0948, -326.6127, -326.9403, 
    -326.9126, -327.2563, -327.51, -328.0608, -328.9427, -328.6115, 
    -329.2209, -329.3531, -328.4177, -328.9846, -327.1605, -327.4544, 
    -327.2803, -326.6379, -328.6863, -327.6351, -329.5875, -329.008, 
    -330.6802, -329.8523, -331.4772, -332.169, -332.8255, -333.5866, 
    -327.1204, -326.8977, -327.2975, -327.8479, -328.3615, -329.0425, 
    -329.1128, -329.24, -329.5813, -329.8592, -329.2792, -329.929, -327.5202, 
    -328.778, -326.8124, -327.4035, -327.8159, -327.6362, -328.5739, 
    -328.7945, -329.7008, -329.228, -331.9973, -330.7762, -334.17, -333.2206, 
    -326.8195, -327.1202, -328.1634, -327.6675, -329.0886, -329.4481, 
    -329.7331, -330.0956, -330.1356, -330.3506, -329.9982, -330.3371, 
    -329.0439, -329.6276, -328.0456, -328.4275, -328.2522, -328.0591, 
    -328.6549, -329.2981, -329.3134, -329.5161, -330.0841, -329.0943, 
    -332.1515, -330.2663, -327.4478, -328.0233, -328.1077, -327.8844, 
    -329.413, -328.8524, -330.3456, -329.9451, -330.6018, -330.2753, 
    -330.2272, -329.8083, -329.5471, -328.8773, -328.3412, -327.917, 
    -328.0158, -328.4818, -329.3372, -330.1384, -329.9626, -330.5519, 
    -328.9854, -329.6472, -329.3947, -330.0533, -328.6023, -329.8338, 
    -328.2895, -328.4243, -328.8415, -329.6901, -329.8784, -330.0761, 
    -329.9545, -329.359, -329.2521, -328.8318, -328.7148, -328.3951, 
    -328.1295, -328.3717, -328.6257, -329.36, -330.0118, -330.7233, 
    -330.8981, -331.7249, -331.0493, -332.1616, -331.2121, -332.8578, 
    -329.9073, -331.1879, -328.8611, -329.111, -329.5713, -330.608, 
    -330.0502, -330.7035, -329.2484, -328.4969, -328.3048, -327.9425, 
    -328.3131, -328.283, -328.6375, -328.5237, -329.3841, -328.9172, 
    -330.2255, -330.6988, -332.0379, -332.8579, -333.6956, -334.0645, 
    -334.177, -334.2239 ;

 FGR12 =
  -224.2574, -224.2202, -224.2273, -224.1978, -224.2139, -224.1947, 
    -224.2495, -224.219, -224.2383, -224.2536, -224.1419, -224.1964, 
    -224.0845, -224.1183, -224.0342, -224.0902, -224.0228, -224.0352, 
    -223.9965, -224.0075, -223.9602, -223.9915, -223.9349, -223.9673, 
    -223.9624, -223.9926, -224.1846, -224.1487, -224.1869, -224.1817, 
    -224.1838, -224.2138, -224.2292, -224.2598, -224.2541, -224.2314, 
    -224.1793, -224.1966, -224.152, -224.1529, -224.1055, -224.1268, 
    -224.0487, -224.0699, -224.007, -224.023, -224.0079, -224.0124, 
    -224.0078, -224.0313, -224.0212, -224.0417, -224.1229, -224.0987, 
    -224.1722, -224.219, -224.2483, -224.2698, -224.2667, -224.2611, 
    -224.2313, -224.2029, -224.1813, -224.167, -224.1531, -224.1137, 
    -224.0916, -224.0446, -224.0526, -224.0386, -224.0246, -224.0019, 
    -224.0055, -223.9957, -224.0386, -224.0102, -224.0573, -224.0444, 
    -224.1517, -224.1918, -224.211, -224.226, -224.2645, -224.2379, 
    -224.2484, -224.2231, -224.2074, -224.2151, -224.1667, -224.1856, 
    -224.0902, -224.1306, -224.0262, -224.0509, -224.0202, -224.0357, 
    -224.0094, -224.0331, -223.9919, -223.9833, -223.9892, -223.9657, 
    -224.0344, -224.0081, -224.2154, -224.2141, -224.2081, -224.2347, 
    -224.2362, -224.2601, -224.2386, -224.2297, -224.2063, -224.1928, 
    -224.1798, -224.1515, -224.1213, -224.0789, -224.0493, -224.0292, 
    -224.0414, -224.0306, -224.0427, -224.0483, -223.9866, -224.0213, 
    -223.9691, -223.9719, -223.9956, -223.9715, -224.2132, -224.2204, 
    -224.2462, -224.226, -224.2626, -224.2424, -224.231, -224.1857, 
    -224.1751, -224.1661, -224.1481, -224.1257, -224.0871, -224.0542, 
    -224.0236, -224.0258, -224.0251, -224.0185, -224.0351, -224.0158, 
    -224.0128, -224.021, -223.9723, -223.9861, -223.9719, -223.9809, 
    -224.218, -224.2059, -224.2125, -224.2001, -224.209, -224.1699, 
    -224.1584, -224.1052, -224.1263, -224.0921, -224.1226, -224.1173, 
    -224.0921, -224.1208, -224.0565, -224.1006, -224.0182, -224.0626, 
    -224.0155, -224.0238, -224.0099, -223.9978, -223.9822, -223.9544, 
    -223.9608, -223.9373, -224.1873, -224.1716, -224.1725, -224.1559, 
    -224.1441, -224.118, -224.0772, -224.0923, -224.0641, -224.0595, 
    -224.1013, -224.0755, -224.1608, -224.1472, -224.1549, -224.1863, 
    -224.0894, -224.1387, -224.0489, -224.0741, -223.9996, -224.0372, 
    -223.9643, -223.935, -223.9056, -223.8741, -224.1626, -224.1733, 
    -224.1539, -224.1286, -224.1041, -224.0726, -224.0692, -224.0634, 
    -224.0489, -224.0363, -224.0621, -224.0331, -224.1451, -224.085, 
    -224.1777, -224.1497, -224.1299, -224.1381, -224.0939, -224.0838, 
    -224.0439, -224.0638, -223.9426, -223.9959, -223.8489, -223.8894, 
    -224.1771, -224.1624, -224.1136, -224.1366, -224.0703, -224.0552, 
    -224.042, -224.0259, -224.0239, -224.0143, -224.03, -224.0148, -224.0725, 
    -224.0469, -224.1186, -224.101, -224.1089, -224.118, -224.0903, 
    -224.0625, -224.0612, -224.0523, -224.0285, -224.07, -223.937, -224.0201, 
    -224.1468, -224.1205, -224.1159, -224.1262, -224.0568, -224.0813, 
    -224.0145, -224.0324, -224.0029, -224.0176, -224.0198, -224.0386, 
    -224.0506, -224.0803, -224.1051, -224.1246, -224.12, -224.0986, 
    -224.0606, -224.024, -224.0321, -224.0051, -224.0751, -224.0463, 
    -224.0579, -224.0276, -224.0929, -224.0395, -224.1072, -224.101, 
    -224.0818, -224.0448, -224.0355, -224.0268, -224.032, -224.0595, 
    -224.063, -224.0821, -224.0878, -224.1023, -224.1147, -224.1035, 
    -224.092, -224.0592, -224.0298, -223.9977, -223.9897, -223.9547, 
    -223.9842, -223.9368, -223.9785, -223.906, -224.0354, -223.9782, 
    -224.0807, -224.0692, -224.0501, -224.0034, -224.0278, -223.999, 
    -224.063, -224.0983, -224.1065, -224.1236, -224.1061, -224.1075, 
    -224.091, -224.0963, -224.0581, -224.0782, -224.02, -223.9991, -223.94, 
    -223.9049, -223.8686, -223.8531, -223.8484, -223.8465 ;

 FGR_R =
  -325.1869, -325.9453, -325.7983, -326.409, -326.0709, -326.4702, -325.3414, 
    -325.9747, -325.5709, -325.2563, -327.5912, -326.4364, -328.7964, 
    -328.0598, -329.9227, -328.6807, -330.1715, -329.889, -330.7437, 
    -330.499, -331.5886, -330.8567, -332.1565, -331.4148, -331.5301, 
    -330.8323, -326.6706, -327.4471, -326.6241, -326.735, -326.6857, 
    -326.0773, -325.7694, -325.1302, -325.2466, -325.7167, -326.7849, 
    -326.4235, -327.3378, -327.3172, -328.332, -327.8745, -329.5914, 
    -329.0965, -330.5092, -330.1562, -330.4923, -330.3906, -330.4936, 
    -329.976, -330.1977, -329.7427, -327.9598, -328.4803, -326.9262, 
    -325.9878, -325.3689, -324.9284, -324.9907, -325.109, -325.7194, 
    -326.295, -326.7328, -327.0255, -327.3142, -328.1817, -328.6447, 
    -329.6886, -329.5035, -329.8182, -330.1211, -330.6276, -330.5445, 
    -330.7672, -329.811, -330.446, -329.3977, -329.6842, -327.3865, 
    -326.5213, -326.1483, -325.8263, -325.0384, -325.5822, -325.3676, 
    -325.8793, -326.2036, -326.0435, -327.0335, -326.6484, -328.6721, 
    -327.8011, -330.0858, -329.5416, -330.2165, -329.8724, -330.4615, 
    -329.9313, -330.8506, -331.0502, -330.9137, -331.44, -329.9018, 
    -330.4917, -326.0387, -326.0648, -326.187, -325.6497, -325.6171, 
    -325.1267, -325.5637, -325.7492, -326.2228, -326.5017, -326.7672, 
    -327.3511, -328.0011, -328.9115, -329.5768, -330.0158, -329.747, 
    -329.9843, -329.7188, -329.5947, -330.975, -330.1994, -331.3643, -331.3, 
    -330.7723, -331.3073, -326.0832, -325.9329, -325.4093, -325.8191, 
    -325.0734, -325.49, -325.7291, -326.6551, -326.86, -327.0481, -327.4209, 
    -327.8979, -328.7341, -329.4728, -330.139, -330.0903, -330.1074, 
    -330.2556, -329.8876, -330.3161, -330.3874, -330.2, -331.2914, -330.9796, 
    -331.2986, -331.0958, -325.9819, -326.235, -326.0981, -326.3551, 
    -326.1736, -326.9789, -327.2203, -328.3501, -327.8882, -328.6251, 
    -327.9635, -328.0804, -328.6466, -327.9996, -329.4315, -328.4552, 
    -330.2614, -329.2836, -330.3219, -330.1361, -330.4443, -330.7196, 
    -331.0671, -331.7067, -331.5589, -332.0948, -326.6127, -326.9403, 
    -326.9126, -327.2563, -327.51, -328.0608, -328.9427, -328.6115, 
    -329.2209, -329.3531, -328.4177, -328.9846, -327.1605, -327.4544, 
    -327.2803, -326.6379, -328.6863, -327.6351, -329.5875, -329.008, 
    -330.6802, -329.8523, -331.4772, -332.169, -332.8255, -333.5866, 
    -327.1204, -326.8977, -327.2975, -327.8479, -328.3615, -329.0425, 
    -329.1128, -329.24, -329.5813, -329.8592, -329.2792, -329.929, -327.5202, 
    -328.778, -326.8124, -327.4035, -327.8159, -327.6362, -328.5739, 
    -328.7945, -329.7008, -329.228, -331.9973, -330.7762, -334.17, -333.2206, 
    -326.8195, -327.1202, -328.1634, -327.6675, -329.0886, -329.4481, 
    -329.7331, -330.0956, -330.1356, -330.3506, -329.9982, -330.3371, 
    -329.0439, -329.6276, -328.0456, -328.4275, -328.2522, -328.0591, 
    -328.6549, -329.2981, -329.3134, -329.5161, -330.0841, -329.0943, 
    -332.1515, -330.2663, -327.4478, -328.0233, -328.1077, -327.8844, 
    -329.413, -328.8524, -330.3456, -329.9451, -330.6018, -330.2753, 
    -330.2272, -329.8083, -329.5471, -328.8773, -328.3412, -327.917, 
    -328.0158, -328.4818, -329.3372, -330.1384, -329.9626, -330.5519, 
    -328.9854, -329.6472, -329.3947, -330.0533, -328.6023, -329.8338, 
    -328.2895, -328.4243, -328.8415, -329.6901, -329.8784, -330.0761, 
    -329.9545, -329.359, -329.2521, -328.8318, -328.7148, -328.3951, 
    -328.1295, -328.3717, -328.6257, -329.36, -330.0118, -330.7233, 
    -330.8981, -331.7249, -331.0493, -332.1616, -331.2121, -332.8578, 
    -329.9073, -331.1879, -328.8611, -329.111, -329.5713, -330.608, 
    -330.0502, -330.7035, -329.2484, -328.4969, -328.3048, -327.9425, 
    -328.3131, -328.283, -328.6375, -328.5237, -329.3841, -328.9172, 
    -330.2255, -330.6988, -332.0379, -332.8579, -333.6956, -334.0645, 
    -334.177, -334.2239 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  74.72346, 74.77625, 74.76602, 74.80855, 74.785, 74.81282, 74.73421, 
    74.7783, 74.75019, 74.72829, 74.89099, 74.81046, 74.97538, 74.92381, 
    75.05312, 74.96728, 75.07053, 75.05077, 75.1106, 75.09346, 75.16971, 
    75.1185, 75.20944, 75.15755, 75.16562, 75.11679, 74.82678, 74.88091, 
    74.82355, 74.83128, 74.82784, 74.78544, 74.76401, 74.71951, 74.72761, 
    74.76035, 74.83475, 74.80957, 74.87328, 74.87184, 74.94286, 74.91084, 
    75.02993, 74.99641, 75.09418, 75.06947, 75.09299, 75.08588, 75.09309, 
    75.05685, 75.07237, 75.04053, 74.91681, 74.95325, 74.8446, 74.77921, 
    74.73613, 74.70546, 74.70979, 74.71803, 74.76053, 74.80061, 74.83112, 
    74.85152, 74.87164, 74.93233, 74.96475, 75.03674, 75.02378, 75.04581, 
    75.06702, 75.10246, 75.09665, 75.11224, 75.04531, 75.08975, 75.01637, 
    75.03643, 74.87667, 74.81638, 74.79038, 74.76797, 74.71312, 74.75098, 
    74.73604, 74.77166, 74.79424, 74.78309, 74.85208, 74.82524, 74.96667, 
    74.90569, 75.06454, 75.02644, 75.07369, 75.04961, 75.09084, 75.05373, 
    75.11808, 75.13203, 75.12249, 75.15932, 75.05166, 75.09296, 74.78275, 
    74.78457, 74.79308, 74.75568, 74.75341, 74.71926, 74.74969, 74.7626, 
    74.79558, 74.81501, 74.83352, 74.87421, 74.91969, 74.98345, 75.02891, 
    75.05965, 75.04083, 75.05743, 75.03886, 75.03017, 75.12678, 75.07249, 
    75.15402, 75.14953, 75.11259, 75.15003, 74.78585, 74.77539, 74.73894, 
    74.76747, 74.71555, 74.74456, 74.7612, 74.82571, 74.83999, 74.8531, 
    74.87909, 74.91247, 74.97102, 75.02163, 75.06827, 75.06486, 75.06606, 
    75.07643, 75.05067, 75.08066, 75.08565, 75.07254, 75.14892, 75.12711, 
    75.14943, 75.13524, 74.7788, 74.79642, 74.7869, 74.80479, 74.79214, 
    74.84827, 74.8651, 74.94413, 74.91179, 74.96339, 74.91706, 74.92525, 
    74.96488, 74.91959, 75.01873, 74.95148, 75.07684, 75.00951, 75.08107, 
    75.06807, 75.08964, 75.10891, 75.13323, 75.17798, 75.16763, 75.20513, 
    74.82275, 74.84558, 74.84366, 74.86761, 74.88532, 74.92388, 74.98564, 
    74.96244, 75.00513, 75.01324, 74.94887, 74.98857, 74.86092, 74.88142, 
    74.86928, 74.82451, 74.96767, 74.89407, 75.02966, 74.99021, 75.10615, 
    75.04819, 75.16192, 75.21031, 75.25624, 75.30946, 74.85813, 74.84261, 
    74.87048, 74.90897, 74.94493, 74.99263, 74.99756, 75.00647, 75.02923, 
    75.04868, 75.00921, 75.05357, 74.88602, 74.9741, 74.83667, 74.87787, 
    74.90673, 74.89415, 74.95981, 74.97526, 75.03759, 75.00562, 75.1983, 
    75.11285, 75.35026, 75.28387, 74.83717, 74.85812, 74.93106, 74.89634, 
    74.99586, 75.0199, 75.03986, 75.06523, 75.06803, 75.08308, 75.05841, 
    75.08213, 74.99273, 75.03246, 74.92281, 74.94955, 74.93728, 74.92376, 
    74.96548, 75.00938, 75.01047, 75.02466, 75.0644, 74.99626, 75.20908, 
    75.07716, 74.88097, 74.92124, 74.92716, 74.91153, 75.01744, 74.97931, 
    75.08273, 75.0547, 75.10066, 75.0778, 75.07444, 75.04512, 75.02682, 
    74.98106, 74.94351, 74.91381, 74.92073, 74.95335, 75.01213, 75.06822, 
    75.05592, 75.09717, 74.98863, 75.03383, 75.01616, 75.06227, 74.96179, 
    75.04688, 74.93989, 74.94933, 74.97855, 75.03683, 75.05003, 75.06387, 
    75.05535, 75.01366, 75.00731, 74.97787, 74.96967, 74.94729, 74.9287, 
    74.94565, 74.96342, 75.01373, 75.05936, 75.10916, 75.1214, 75.17924, 
    75.13197, 75.20979, 75.14334, 75.25848, 75.05204, 75.14166, 74.97992, 
    74.99743, 75.02852, 75.10109, 75.06206, 75.10777, 75.00706, 74.95441, 
    74.94096, 74.9156, 74.94154, 74.93944, 74.96426, 74.95629, 75.01542, 
    74.98386, 75.07432, 75.10744, 75.20115, 75.25851, 75.31709, 75.34289, 
    75.35075, 75.35403 ;

 FIRA_R =
  74.72346, 74.77625, 74.76602, 74.80855, 74.785, 74.81282, 74.73421, 
    74.7783, 74.75019, 74.72829, 74.89099, 74.81046, 74.97538, 74.92381, 
    75.05312, 74.96728, 75.07053, 75.05077, 75.1106, 75.09346, 75.16971, 
    75.1185, 75.20944, 75.15755, 75.16562, 75.11679, 74.82678, 74.88091, 
    74.82355, 74.83128, 74.82784, 74.78544, 74.76401, 74.71951, 74.72761, 
    74.76035, 74.83475, 74.80957, 74.87328, 74.87184, 74.94286, 74.91084, 
    75.02993, 74.99641, 75.09418, 75.06947, 75.09299, 75.08588, 75.09309, 
    75.05685, 75.07237, 75.04053, 74.91681, 74.95325, 74.8446, 74.77921, 
    74.73613, 74.70546, 74.70979, 74.71803, 74.76053, 74.80061, 74.83112, 
    74.85152, 74.87164, 74.93233, 74.96475, 75.03674, 75.02378, 75.04581, 
    75.06702, 75.10246, 75.09665, 75.11224, 75.04531, 75.08975, 75.01637, 
    75.03643, 74.87667, 74.81638, 74.79038, 74.76797, 74.71312, 74.75098, 
    74.73604, 74.77166, 74.79424, 74.78309, 74.85208, 74.82524, 74.96667, 
    74.90569, 75.06454, 75.02644, 75.07369, 75.04961, 75.09084, 75.05373, 
    75.11808, 75.13203, 75.12249, 75.15932, 75.05166, 75.09296, 74.78275, 
    74.78457, 74.79308, 74.75568, 74.75341, 74.71926, 74.74969, 74.7626, 
    74.79558, 74.81501, 74.83352, 74.87421, 74.91969, 74.98345, 75.02891, 
    75.05965, 75.04083, 75.05743, 75.03886, 75.03017, 75.12678, 75.07249, 
    75.15402, 75.14953, 75.11259, 75.15003, 74.78585, 74.77539, 74.73894, 
    74.76747, 74.71555, 74.74456, 74.7612, 74.82571, 74.83999, 74.8531, 
    74.87909, 74.91247, 74.97102, 75.02163, 75.06827, 75.06486, 75.06606, 
    75.07643, 75.05067, 75.08066, 75.08565, 75.07254, 75.14892, 75.12711, 
    75.14943, 75.13524, 74.7788, 74.79642, 74.7869, 74.80479, 74.79214, 
    74.84827, 74.8651, 74.94413, 74.91179, 74.96339, 74.91706, 74.92525, 
    74.96488, 74.91959, 75.01873, 74.95148, 75.07684, 75.00951, 75.08107, 
    75.06807, 75.08964, 75.10891, 75.13323, 75.17798, 75.16763, 75.20513, 
    74.82275, 74.84558, 74.84366, 74.86761, 74.88532, 74.92388, 74.98564, 
    74.96244, 75.00513, 75.01324, 74.94887, 74.98857, 74.86092, 74.88142, 
    74.86928, 74.82451, 74.96767, 74.89407, 75.02966, 74.99021, 75.10615, 
    75.04819, 75.16192, 75.21031, 75.25624, 75.30946, 74.85813, 74.84261, 
    74.87048, 74.90897, 74.94493, 74.99263, 74.99756, 75.00647, 75.02923, 
    75.04868, 75.00921, 75.05357, 74.88602, 74.9741, 74.83667, 74.87787, 
    74.90673, 74.89415, 74.95981, 74.97526, 75.03759, 75.00562, 75.1983, 
    75.11285, 75.35026, 75.28387, 74.83717, 74.85812, 74.93106, 74.89634, 
    74.99586, 75.0199, 75.03986, 75.06523, 75.06803, 75.08308, 75.05841, 
    75.08213, 74.99273, 75.03246, 74.92281, 74.94955, 74.93728, 74.92376, 
    74.96548, 75.00938, 75.01047, 75.02466, 75.0644, 74.99626, 75.20908, 
    75.07716, 74.88097, 74.92124, 74.92716, 74.91153, 75.01744, 74.97931, 
    75.08273, 75.0547, 75.10066, 75.0778, 75.07444, 75.04512, 75.02682, 
    74.98106, 74.94351, 74.91381, 74.92073, 74.95335, 75.01213, 75.06822, 
    75.05592, 75.09717, 74.98863, 75.03383, 75.01616, 75.06227, 74.96179, 
    75.04688, 74.93989, 74.94933, 74.97855, 75.03683, 75.05003, 75.06387, 
    75.05535, 75.01366, 75.00731, 74.97787, 74.96967, 74.94729, 74.9287, 
    74.94565, 74.96342, 75.01373, 75.05936, 75.10916, 75.1214, 75.17924, 
    75.13197, 75.20979, 75.14334, 75.25848, 75.05204, 75.14166, 74.97992, 
    74.99743, 75.02852, 75.10109, 75.06206, 75.10777, 75.00706, 74.95441, 
    74.94096, 74.9156, 74.94154, 74.93944, 74.96426, 74.95629, 75.01542, 
    74.98386, 75.07432, 75.10744, 75.20115, 75.25851, 75.31709, 75.34289, 
    75.35075, 75.35403 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  263.6844, 263.7372, 263.727, 263.7695, 263.7459, 263.7738, 263.6952, 
    263.7392, 263.7111, 263.6892, 263.8519, 263.7714, 263.9363, 263.8847, 
    264.0141, 263.9282, 264.0315, 264.0117, 264.0715, 264.0544, 264.1306, 
    264.0794, 264.1704, 264.1185, 264.1266, 264.0777, 263.7877, 263.8419, 
    263.7845, 263.7922, 263.7888, 263.7464, 263.7249, 263.6805, 263.6885, 
    263.7213, 263.7957, 263.7705, 263.8342, 263.8328, 263.9038, 263.8718, 
    263.9909, 263.9574, 264.0551, 264.0304, 264.0539, 264.0468, 264.054, 
    264.0178, 264.0333, 264.0015, 263.8777, 263.9142, 263.8055, 263.7401, 
    263.6971, 263.6664, 263.6707, 263.679, 263.7215, 263.7615, 263.7921, 
    263.8125, 263.8326, 263.8933, 263.9257, 263.9977, 263.9847, 264.0067, 
    264.028, 264.0634, 264.0576, 264.0732, 264.0063, 264.0507, 263.9773, 
    263.9974, 263.8376, 263.7773, 263.7513, 263.7289, 263.674, 263.7119, 
    263.697, 263.7326, 263.7552, 263.744, 263.813, 263.7862, 263.9276, 
    263.8666, 264.0255, 263.9874, 264.0346, 264.0106, 264.0518, 264.0147, 
    264.079, 264.093, 264.0834, 264.1203, 264.0126, 264.0539, 263.7437, 
    263.7455, 263.754, 263.7166, 263.7144, 263.6802, 263.7106, 263.7235, 
    263.7565, 263.7759, 263.7945, 263.8351, 263.8806, 263.9444, 263.9898, 
    264.0206, 264.0018, 264.0184, 263.9998, 263.9911, 264.0877, 264.0334, 
    264.115, 264.1105, 264.0735, 264.111, 263.7468, 263.7363, 263.6999, 
    263.7284, 263.6765, 263.7055, 263.7221, 263.7867, 263.8009, 263.814, 
    263.84, 263.8734, 263.9319, 263.9826, 264.0292, 264.0258, 264.027, 
    264.0374, 264.0116, 264.0416, 264.0466, 264.0335, 264.1099, 264.088, 
    264.1104, 264.0962, 263.7397, 263.7574, 263.7478, 263.7657, 263.7531, 
    263.8092, 263.826, 263.9051, 263.8727, 263.9243, 263.878, 263.8862, 
    263.9258, 263.8805, 263.9797, 263.9124, 264.0378, 263.9705, 264.042, 
    264.029, 264.0506, 264.0699, 264.0942, 264.1389, 264.1286, 264.1661, 
    263.7837, 263.8065, 263.8046, 263.8286, 263.8463, 263.8848, 263.9466, 
    263.9234, 263.9661, 263.9742, 263.9098, 263.9495, 263.8219, 263.8424, 
    263.8302, 263.7854, 263.9286, 263.855, 263.9906, 263.9511, 264.0671, 
    264.0091, 264.1229, 264.1713, 264.2172, 264.2704, 263.8191, 263.8036, 
    263.8314, 263.8699, 263.9059, 263.9536, 263.9585, 263.9674, 263.9902, 
    264.0096, 263.9702, 264.0145, 263.847, 263.935, 263.7976, 263.8388, 
    263.8677, 263.8551, 263.9207, 263.9362, 263.9985, 263.9666, 264.1592, 
    264.0738, 264.3112, 264.2448, 263.7981, 263.8191, 263.892, 263.8573, 
    263.9568, 263.9808, 264.0008, 264.0262, 264.029, 264.044, 264.0193, 
    264.0431, 263.9537, 263.9934, 263.8838, 263.9105, 263.8982, 263.8847, 
    263.9264, 263.9703, 263.9714, 263.9856, 264.0253, 263.9572, 264.17, 
    264.0381, 263.8419, 263.8822, 263.8881, 263.8725, 263.9784, 263.9402, 
    264.0437, 264.0156, 264.0616, 264.0388, 264.0354, 264.006, 263.9878, 
    263.942, 263.9044, 263.8748, 263.8817, 263.9143, 263.9731, 264.0292, 
    264.0168, 264.0581, 263.9496, 263.9948, 263.9771, 264.0232, 263.9227, 
    264.0078, 263.9008, 263.9103, 263.9395, 263.9978, 264.011, 264.0248, 
    264.0163, 263.9746, 263.9683, 263.9388, 263.9306, 263.9082, 263.8896, 
    263.9066, 263.9244, 263.9747, 264.0203, 264.0701, 264.0823, 264.1402, 
    264.0929, 264.1707, 264.1043, 264.2194, 264.013, 264.1026, 263.9409, 
    263.9584, 263.9895, 264.062, 264.023, 264.0687, 263.968, 263.9153, 
    263.9019, 263.8765, 263.9025, 263.9004, 263.9252, 263.9172, 263.9763, 
    263.9448, 264.0352, 264.0684, 264.1621, 264.2195, 264.278, 264.3038, 
    264.3117, 264.315 ;

 FLDS =
  188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSA_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658 ;

 FSDSND =
  0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004 ;

 FSDSNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSDSNI =
  0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284 ;

 FSDSVD =
  0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081 ;

 FSDSVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSDSVI =
  0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228 ;

 FSDSVILN =
  0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012 ;

 FSH =
  244.1978, 244.8872, 244.7535, 245.3086, 245.0014, 245.3643, 244.3383, 
    244.9139, 244.5469, 244.2609, 246.3831, 245.3335, 247.4779, 246.8088, 
    248.5007, 247.3728, 248.7267, 248.4701, 249.2464, 249.0241, 250.0138, 
    249.3491, 250.5295, 249.8559, 249.9607, 249.3269, 245.5464, 246.2521, 
    245.5042, 245.6049, 245.5601, 245.0071, 244.7273, 244.1463, 244.2521, 
    244.6794, 245.6503, 245.3219, 246.1528, 246.1341, 247.056, 246.6404, 
    248.1998, 247.7505, 249.0334, 248.7128, 249.0181, 248.9257, 249.0193, 
    248.5491, 248.7505, 248.3373, 246.7179, 247.1907, 245.7787, 244.9258, 
    244.3633, 243.9629, 244.0195, 244.127, 244.6819, 245.205, 245.603, 
    245.869, 246.1313, 246.9195, 247.3401, 248.2881, 248.12, 248.4058, 
    248.681, 249.141, 249.0655, 249.2678, 248.3993, 248.976, 248.0239, 
    248.2841, 246.1971, 245.4107, 245.0717, 244.779, 244.0629, 244.5571, 
    244.3621, 244.8272, 245.1219, 244.9764, 245.8763, 245.5262, 247.365, 
    246.5737, 248.6489, 248.1546, 248.7675, 248.455, 248.9901, 248.5085, 
    249.3436, 249.5248, 249.4008, 249.8788, 248.4817, 249.0176, 244.9721, 
    244.9958, 245.1068, 244.6185, 244.5889, 244.1431, 244.5403, 244.709, 
    245.1395, 245.3929, 245.6342, 246.1649, 246.7554, 247.5825, 248.1866, 
    248.5853, 248.3412, 248.5567, 248.3156, 248.2028, 249.4565, 248.752, 
    249.8101, 249.7517, 249.2724, 249.7583, 245.0125, 244.8759, 244.4, 
    244.7724, 244.0946, 244.4733, 244.6906, 245.5323, 245.7185, 245.8895, 
    246.2283, 246.6617, 247.4213, 248.0921, 248.6972, 248.653, 248.6685, 
    248.8031, 248.4689, 248.858, 248.9228, 248.7526, 249.7439, 249.4607, 
    249.7505, 249.5662, 244.9205, 245.1505, 245.0261, 245.2597, 245.0947, 
    245.8266, 246.0461, 247.0725, 246.6528, 247.3223, 246.7212, 246.8274, 
    247.3418, 246.7541, 248.0545, 247.1679, 248.8083, 247.9204, 248.8633, 
    248.6946, 248.9745, 249.2245, 249.5402, 250.1211, 249.9868, 250.4735, 
    245.4938, 245.7916, 245.7664, 246.0788, 246.3093, 246.8097, 247.6108, 
    247.3099, 247.8635, 247.9833, 247.1339, 247.6488, 245.9917, 246.2587, 
    246.1006, 245.5167, 247.3779, 246.4229, 248.1962, 247.6701, 249.1888, 
    248.4368, 249.9126, 250.5409, 251.1371, 251.8283, 245.9552, 245.7528, 
    246.1162, 246.6162, 247.0828, 247.7014, 247.7653, 247.8809, 248.1907, 
    248.443, 247.9164, 248.5064, 246.3185, 247.4612, 245.6753, 246.2125, 
    246.5872, 246.4239, 247.2758, 247.4762, 248.2992, 247.8699, 250.3849, 
    249.2759, 252.3581, 251.4959, 245.6818, 245.955, 246.9029, 246.4524, 
    247.7433, 248.0696, 248.3285, 248.6578, 248.6941, 248.8894, 248.5693, 
    248.8771, 247.7027, 248.2326, 246.7958, 247.1428, 246.9835, 246.8081, 
    247.3494, 247.9333, 247.9473, 248.1314, 248.6473, 247.7485, 250.525, 
    248.8128, 246.2527, 246.7756, 246.8523, 246.6494, 248.0378, 247.5287, 
    248.8848, 248.5211, 249.1175, 248.821, 248.7773, 248.3968, 248.1595, 
    247.5513, 247.0644, 246.679, 246.7688, 247.1921, 247.9689, 248.6967, 
    248.537, 249.0722, 247.6496, 248.2504, 248.0211, 248.6194, 247.3016, 
    248.42, 247.0174, 247.1399, 247.5188, 248.2895, 248.4605, 248.6401, 
    248.5296, 247.9887, 247.8918, 247.51, 247.4038, 247.1134, 246.8721, 
    247.0921, 247.3228, 247.9896, 248.5817, 249.2279, 249.3866, 250.1376, 
    249.524, 250.5342, 249.6718, 251.1664, 248.4867, 249.6499, 247.5366, 
    247.7636, 248.1816, 249.1232, 248.6166, 249.2099, 247.8885, 247.2059, 
    247.0313, 246.7022, 247.0388, 247.0115, 247.3336, 247.2302, 248.0115, 
    247.5877, 248.7757, 249.2056, 250.4219, 251.1665, 251.9273, 252.2623, 
    252.3644, 252.407 ;

 FSH_G =
  257.464, 258.1543, 258.0204, 258.5763, 258.2686, 258.632, 257.6047, 
    258.181, 257.8135, 257.5271, 259.6521, 258.6012, 260.7484, 260.0785, 
    261.7726, 260.6432, 261.9989, 261.7419, 262.5193, 262.2967, 263.2877, 
    262.6221, 263.8042, 263.1296, 263.2345, 262.5999, 258.8144, 259.521, 
    258.7721, 258.873, 258.8281, 258.2744, 257.9941, 257.4124, 257.5183, 
    257.9462, 258.9184, 258.5895, 259.4216, 259.4029, 260.326, 259.9099, 
    261.4713, 261.0214, 262.3061, 261.985, 262.2907, 262.1982, 262.2919, 
    261.8211, 262.0227, 261.6089, 259.9875, 260.4609, 259.047, 258.1929, 
    257.6296, 257.2287, 257.2854, 257.3931, 257.9487, 258.4725, 258.8711, 
    259.1374, 259.4001, 260.1893, 260.6104, 261.5597, 261.3914, 261.6776, 
    261.9531, 262.4137, 262.3381, 262.5407, 261.6711, 262.2485, 261.2952, 
    261.5557, 259.4659, 258.6785, 258.339, 258.046, 257.3288, 257.8238, 
    257.6285, 258.0942, 258.3893, 258.2436, 259.1447, 258.7942, 260.6354, 
    259.8431, 261.921, 261.426, 262.0398, 261.7269, 262.2626, 261.7805, 
    262.6166, 262.798, 262.6739, 263.1526, 261.7536, 262.2902, 258.2393, 
    258.263, 258.3742, 257.8852, 257.8556, 257.4092, 257.8069, 257.9758, 
    258.4069, 258.6607, 258.9023, 259.4337, 260.025, 260.8531, 261.458, 
    261.8573, 261.6129, 261.8286, 261.5872, 261.4743, 262.7297, 262.0242, 
    263.0837, 263.0253, 262.5453, 263.0319, 258.2798, 258.143, 257.6664, 
    258.0394, 257.3607, 257.7398, 257.9575, 258.8003, 258.9868, 259.1579, 
    259.4972, 259.9311, 260.6917, 261.3634, 261.9694, 261.9251, 261.9406, 
    262.0754, 261.7408, 262.1304, 262.1953, 262.0248, 263.0174, 262.7339, 
    263.024, 262.8396, 258.1876, 258.4179, 258.2934, 258.5273, 258.3621, 
    259.095, 259.3147, 260.3425, 259.9223, 260.5926, 259.9908, 260.0971, 
    260.6121, 260.0237, 261.3258, 260.438, 262.0807, 261.1915, 262.1357, 
    261.9667, 262.247, 262.4974, 262.8135, 263.3951, 263.2607, 263.748, 
    258.7617, 259.0599, 259.0347, 259.3475, 259.5783, 260.0793, 260.8815, 
    260.5803, 261.1346, 261.2545, 260.404, 260.9196, 259.2603, 259.5276, 
    259.3693, 258.7846, 260.6483, 259.6921, 261.4677, 260.9409, 262.4616, 
    261.7086, 263.1864, 263.8155, 264.4126, 265.1046, 259.2238, 259.0211, 
    259.385, 259.8856, 260.3528, 260.9723, 261.0362, 261.1519, 261.4622, 
    261.7149, 261.1875, 261.7783, 259.5875, 260.7317, 258.9434, 259.4814, 
    259.8566, 259.6931, 260.5461, 260.7467, 261.5708, 261.141, 263.6593, 
    262.5488, 265.6352, 264.7719, 258.95, 259.2236, 260.1727, 259.7216, 
    261.0142, 261.3409, 261.6002, 261.9299, 261.9663, 262.1618, 261.8413, 
    262.1495, 260.9736, 261.5042, 260.0655, 260.4129, 260.2534, 260.0778, 
    260.6198, 261.2045, 261.2185, 261.4028, 261.9193, 261.0194, 263.7996, 
    262.0851, 259.5217, 260.0452, 260.122, 259.9189, 261.3091, 260.7993, 
    262.1573, 261.793, 262.3903, 262.0933, 262.0496, 261.6686, 261.431, 
    260.822, 260.3344, 259.9485, 260.0384, 260.4623, 261.2401, 261.9688, 
    261.8089, 262.3449, 260.9204, 261.522, 261.2924, 261.8914, 260.5719, 
    261.6917, 260.2874, 260.4101, 260.7894, 261.5611, 261.7323, 261.9122, 
    261.8015, 261.2599, 261.1629, 260.7806, 260.6743, 260.3835, 260.1419, 
    260.3622, 260.5932, 261.2609, 261.8537, 262.5007, 262.6597, 263.4116, 
    262.7972, 263.8087, 262.9452, 264.4419, 261.7586, 262.9233, 260.8073, 
    261.0346, 261.453, 262.3959, 261.8886, 262.4827, 261.1596, 260.4761, 
    260.3013, 259.9717, 260.3088, 260.2815, 260.6039, 260.5004, 261.2827, 
    260.8584, 262.048, 262.4785, 263.6964, 264.442, 265.2039, 265.5393, 
    265.6416, 265.6842 ;

 FSH_NODYNLNDUSE =
  244.1978, 244.8872, 244.7535, 245.3086, 245.0014, 245.3643, 244.3383, 
    244.9139, 244.5469, 244.2609, 246.3831, 245.3335, 247.4779, 246.8088, 
    248.5007, 247.3728, 248.7267, 248.4701, 249.2464, 249.0241, 250.0138, 
    249.3491, 250.5295, 249.8559, 249.9607, 249.3269, 245.5464, 246.2521, 
    245.5042, 245.6049, 245.5601, 245.0071, 244.7273, 244.1463, 244.2521, 
    244.6794, 245.6503, 245.3219, 246.1528, 246.1341, 247.056, 246.6404, 
    248.1998, 247.7505, 249.0334, 248.7128, 249.0181, 248.9257, 249.0193, 
    248.5491, 248.7505, 248.3373, 246.7179, 247.1907, 245.7787, 244.9258, 
    244.3633, 243.9629, 244.0195, 244.127, 244.6819, 245.205, 245.603, 
    245.869, 246.1313, 246.9195, 247.3401, 248.2881, 248.12, 248.4058, 
    248.681, 249.141, 249.0655, 249.2678, 248.3993, 248.976, 248.0239, 
    248.2841, 246.1971, 245.4107, 245.0717, 244.779, 244.0629, 244.5571, 
    244.3621, 244.8272, 245.1219, 244.9764, 245.8763, 245.5262, 247.365, 
    246.5737, 248.6489, 248.1546, 248.7675, 248.455, 248.9901, 248.5085, 
    249.3436, 249.5248, 249.4008, 249.8788, 248.4817, 249.0176, 244.9721, 
    244.9958, 245.1068, 244.6185, 244.5889, 244.1431, 244.5403, 244.709, 
    245.1395, 245.3929, 245.6342, 246.1649, 246.7554, 247.5825, 248.1866, 
    248.5853, 248.3412, 248.5567, 248.3156, 248.2028, 249.4565, 248.752, 
    249.8101, 249.7517, 249.2724, 249.7583, 245.0125, 244.8759, 244.4, 
    244.7724, 244.0946, 244.4733, 244.6906, 245.5323, 245.7185, 245.8895, 
    246.2283, 246.6617, 247.4213, 248.0921, 248.6972, 248.653, 248.6685, 
    248.8031, 248.4689, 248.858, 248.9228, 248.7526, 249.7439, 249.4607, 
    249.7505, 249.5662, 244.9205, 245.1505, 245.0261, 245.2597, 245.0947, 
    245.8266, 246.0461, 247.0725, 246.6528, 247.3223, 246.7212, 246.8274, 
    247.3418, 246.7541, 248.0545, 247.1679, 248.8083, 247.9204, 248.8633, 
    248.6946, 248.9745, 249.2245, 249.5402, 250.1211, 249.9868, 250.4735, 
    245.4938, 245.7916, 245.7664, 246.0788, 246.3093, 246.8097, 247.6108, 
    247.3099, 247.8635, 247.9833, 247.1339, 247.6488, 245.9917, 246.2587, 
    246.1006, 245.5167, 247.3779, 246.4229, 248.1962, 247.6701, 249.1888, 
    248.4368, 249.9126, 250.5409, 251.1371, 251.8283, 245.9552, 245.7528, 
    246.1162, 246.6162, 247.0828, 247.7014, 247.7653, 247.8809, 248.1907, 
    248.443, 247.9164, 248.5064, 246.3185, 247.4612, 245.6753, 246.2125, 
    246.5872, 246.4239, 247.2758, 247.4762, 248.2992, 247.8699, 250.3849, 
    249.2759, 252.3581, 251.4959, 245.6818, 245.955, 246.9029, 246.4524, 
    247.7433, 248.0696, 248.3285, 248.6578, 248.6941, 248.8894, 248.5693, 
    248.8771, 247.7027, 248.2326, 246.7958, 247.1428, 246.9835, 246.8081, 
    247.3494, 247.9333, 247.9473, 248.1314, 248.6473, 247.7485, 250.525, 
    248.8128, 246.2527, 246.7756, 246.8523, 246.6494, 248.0378, 247.5287, 
    248.8848, 248.5211, 249.1175, 248.821, 248.7773, 248.3968, 248.1595, 
    247.5513, 247.0644, 246.679, 246.7688, 247.1921, 247.9689, 248.6967, 
    248.537, 249.0722, 247.6496, 248.2504, 248.0211, 248.6194, 247.3016, 
    248.42, 247.0174, 247.1399, 247.5188, 248.2895, 248.4605, 248.6401, 
    248.5296, 247.9887, 247.8918, 247.51, 247.4038, 247.1134, 246.8721, 
    247.0921, 247.3228, 247.9896, 248.5817, 249.2279, 249.3866, 250.1376, 
    249.524, 250.5342, 249.6718, 251.1664, 248.4867, 249.6499, 247.5366, 
    247.7636, 248.1816, 249.1232, 248.6166, 249.2099, 247.8885, 247.2059, 
    247.0313, 246.7022, 247.0388, 247.0115, 247.3336, 247.2302, 248.0115, 
    247.5877, 248.7757, 249.2056, 250.4219, 251.1665, 251.9273, 252.2623, 
    252.3644, 252.407 ;

 FSH_R =
  244.1978, 244.8872, 244.7535, 245.3086, 245.0014, 245.3643, 244.3383, 
    244.9139, 244.5469, 244.2609, 246.3831, 245.3335, 247.4779, 246.8088, 
    248.5007, 247.3728, 248.7267, 248.4701, 249.2464, 249.0241, 250.0138, 
    249.3491, 250.5295, 249.8559, 249.9607, 249.3269, 245.5464, 246.2521, 
    245.5042, 245.6049, 245.5601, 245.0071, 244.7273, 244.1463, 244.2521, 
    244.6794, 245.6503, 245.3219, 246.1528, 246.1341, 247.056, 246.6404, 
    248.1998, 247.7505, 249.0334, 248.7128, 249.0181, 248.9257, 249.0193, 
    248.5491, 248.7505, 248.3373, 246.7179, 247.1907, 245.7787, 244.9258, 
    244.3633, 243.9629, 244.0195, 244.127, 244.6819, 245.205, 245.603, 
    245.869, 246.1313, 246.9195, 247.3401, 248.2881, 248.12, 248.4058, 
    248.681, 249.141, 249.0655, 249.2678, 248.3993, 248.976, 248.0239, 
    248.2841, 246.1971, 245.4107, 245.0717, 244.779, 244.0629, 244.5571, 
    244.3621, 244.8272, 245.1219, 244.9764, 245.8763, 245.5262, 247.365, 
    246.5737, 248.6489, 248.1546, 248.7675, 248.455, 248.9901, 248.5085, 
    249.3436, 249.5248, 249.4008, 249.8788, 248.4817, 249.0176, 244.9721, 
    244.9958, 245.1068, 244.6185, 244.5889, 244.1431, 244.5403, 244.709, 
    245.1395, 245.3929, 245.6342, 246.1649, 246.7554, 247.5825, 248.1866, 
    248.5853, 248.3412, 248.5567, 248.3156, 248.2028, 249.4565, 248.752, 
    249.8101, 249.7517, 249.2724, 249.7583, 245.0125, 244.8759, 244.4, 
    244.7724, 244.0946, 244.4733, 244.6906, 245.5323, 245.7185, 245.8895, 
    246.2283, 246.6617, 247.4213, 248.0921, 248.6972, 248.653, 248.6685, 
    248.8031, 248.4689, 248.858, 248.9228, 248.7526, 249.7439, 249.4607, 
    249.7505, 249.5662, 244.9205, 245.1505, 245.0261, 245.2597, 245.0947, 
    245.8266, 246.0461, 247.0725, 246.6528, 247.3223, 246.7212, 246.8274, 
    247.3418, 246.7541, 248.0545, 247.1679, 248.8083, 247.9204, 248.8633, 
    248.6946, 248.9745, 249.2245, 249.5402, 250.1211, 249.9868, 250.4735, 
    245.4938, 245.7916, 245.7664, 246.0788, 246.3093, 246.8097, 247.6108, 
    247.3099, 247.8635, 247.9833, 247.1339, 247.6488, 245.9917, 246.2587, 
    246.1006, 245.5167, 247.3779, 246.4229, 248.1962, 247.6701, 249.1888, 
    248.4368, 249.9126, 250.5409, 251.1371, 251.8283, 245.9552, 245.7528, 
    246.1162, 246.6162, 247.0828, 247.7014, 247.7653, 247.8809, 248.1907, 
    248.443, 247.9164, 248.5064, 246.3185, 247.4612, 245.6753, 246.2125, 
    246.5872, 246.4239, 247.2758, 247.4762, 248.2992, 247.8699, 250.3849, 
    249.2759, 252.3581, 251.4959, 245.6818, 245.955, 246.9029, 246.4524, 
    247.7433, 248.0696, 248.3285, 248.6578, 248.6941, 248.8894, 248.5693, 
    248.8771, 247.7027, 248.2326, 246.7958, 247.1428, 246.9835, 246.8081, 
    247.3494, 247.9333, 247.9473, 248.1314, 248.6473, 247.7485, 250.525, 
    248.8128, 246.2527, 246.7756, 246.8523, 246.6494, 248.0378, 247.5287, 
    248.8848, 248.5211, 249.1175, 248.821, 248.7773, 248.3968, 248.1595, 
    247.5513, 247.0644, 246.679, 246.7688, 247.1921, 247.9689, 248.6967, 
    248.537, 249.0722, 247.6496, 248.2504, 248.0211, 248.6194, 247.3016, 
    248.42, 247.0174, 247.1399, 247.5188, 248.2895, 248.4605, 248.6401, 
    248.5296, 247.9887, 247.8918, 247.51, 247.4038, 247.1134, 246.8721, 
    247.0921, 247.3228, 247.9896, 248.5817, 249.2279, 249.3866, 250.1376, 
    249.524, 250.5342, 249.6718, 251.1664, 248.4867, 249.6499, 247.5366, 
    247.7636, 248.1816, 249.1232, 248.6166, 249.2099, 247.8885, 247.2059, 
    247.0313, 246.7022, 247.0388, 247.0115, 247.3336, 247.2302, 248.0115, 
    247.5877, 248.7757, 249.2056, 250.4219, 251.1665, 251.9273, 252.2623, 
    252.3644, 252.407 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -13.26616, -13.26709, -13.26691, -13.26765, -13.26725, -13.26773, 
    -13.26636, -13.26712, -13.26664, -13.26625, -13.26907, -13.26769, 
    -13.27055, -13.26967, -13.27188, -13.2704, -13.27219, -13.27186, 
    -13.2729, -13.2726, -13.2739, -13.27304, -13.27461, -13.27371, -13.27384, 
    -13.27301, -13.26798, -13.26889, -13.26793, -13.26806, -13.268, 
    -13.26725, -13.26686, -13.2661, -13.26624, -13.26681, -13.26812, 
    -13.26768, -13.26881, -13.26879, -13.27, -13.26945, -13.2715, -13.27093, 
    -13.27262, -13.27218, -13.27259, -13.27247, -13.27259, -13.27196, 
    -13.27223, -13.27168, -13.26955, -13.27018, -13.2683, -13.26712, 
    -13.26639, -13.26585, -13.26593, -13.26607, -13.26681, -13.26753, 
    -13.26807, -13.26843, -13.26878, -13.26979, -13.27036, -13.27161, 
    -13.2714, -13.27177, -13.27214, -13.27275, -13.27266, -13.27292, 
    -13.27177, -13.27253, -13.27127, -13.27161, -13.26882, -13.2678, 
    -13.26732, -13.26694, -13.26598, -13.26664, -13.26638, -13.26702, 
    -13.26741, -13.26722, -13.26844, -13.26796, -13.2704, -13.26936, 
    -13.2721, -13.27144, -13.27226, -13.27184, -13.27255, -13.27191, 
    -13.27303, -13.27326, -13.2731, -13.27375, -13.27188, -13.27259, 
    -13.26721, -13.26724, -13.2674, -13.26672, -13.26669, -13.26609, 
    -13.26663, -13.26685, -13.26744, -13.26778, -13.2681, -13.26882, 
    -13.2696, -13.27069, -13.27148, -13.27202, -13.27169, -13.27198, 
    -13.27166, -13.27151, -13.27317, -13.27223, -13.27365, -13.27358, 
    -13.27293, -13.27359, -13.26727, -13.26708, -13.26644, -13.26694, 
    -13.26603, -13.26653, -13.26682, -13.26796, -13.26822, -13.26845, 
    -13.26891, -13.26948, -13.27048, -13.27135, -13.27217, -13.27211, 
    -13.27213, -13.2723, -13.27186, -13.27238, -13.27246, -13.27224, 
    -13.27357, -13.27319, -13.27358, -13.27333, -13.26715, -13.26745, 
    -13.26729, -13.2676, -13.26737, -13.26835, -13.26864, -13.27001, 
    -13.26947, -13.27035, -13.26956, -13.2697, -13.27035, -13.26961, 
    -13.27129, -13.27013, -13.27231, -13.27112, -13.27239, -13.27216, 
    -13.27254, -13.27287, -13.27329, -13.27406, -13.27389, -13.27454, 
    -13.26792, -13.26831, -13.26829, -13.26871, -13.26901, -13.26968, 
    -13.27074, -13.27034, -13.27108, -13.27121, -13.27011, -13.27078, 
    -13.26858, -13.26893, -13.26873, -13.26794, -13.27042, -13.26915, 
    -13.27149, -13.27082, -13.27282, -13.2718, -13.27379, -13.27461, 
    -13.27545, -13.27636, -13.26854, -13.26827, -13.26876, -13.26941, 
    -13.27004, -13.27086, -13.27095, -13.2711, -13.27149, -13.27183, 
    -13.27113, -13.27191, -13.26899, -13.27053, -13.26816, -13.26887, 
    -13.26938, -13.26917, -13.2703, -13.27056, -13.27162, -13.27109, 
    -13.2744, -13.27292, -13.2771, -13.27592, -13.26817, -13.26854, 
    -13.26979, -13.26921, -13.27092, -13.27133, -13.27168, -13.27211, 
    -13.27216, -13.27242, -13.272, -13.27241, -13.27086, -13.27155, 
    -13.26966, -13.27012, -13.26991, -13.26968, -13.2704, -13.27113, 
    -13.27117, -13.2714, -13.27204, -13.27092, -13.27455, -13.27226, 
    -13.26894, -13.26962, -13.26973, -13.26947, -13.27128, -13.27063, 
    -13.27241, -13.27193, -13.27273, -13.27233, -13.27227, -13.27177, 
    -13.27145, -13.27066, -13.27001, -13.26951, -13.26963, -13.27018, 
    -13.27118, -13.27216, -13.27194, -13.27267, -13.27079, -13.27156, 
    -13.27125, -13.27206, -13.27033, -13.27174, -13.26996, -13.27012, 
    -13.27062, -13.2716, -13.27185, -13.27208, -13.27194, -13.27121, 
    -13.27111, -13.27061, -13.27046, -13.27009, -13.26977, -13.27005, 
    -13.27035, -13.27122, -13.272, -13.27287, -13.27309, -13.27406, 
    -13.27324, -13.27456, -13.2734, -13.27544, -13.27185, -13.2734, 
    -13.27065, -13.27095, -13.27146, -13.27271, -13.27206, -13.27283, 
    -13.27111, -13.27019, -13.26998, -13.26954, -13.26999, -13.26995, 
    -13.27038, -13.27024, -13.27125, -13.27071, -13.27226, -13.27283, 
    -13.27447, -13.27547, -13.27652, -13.27698, -13.27712, -13.27718 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658 ;

 FSRND =
  0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004 ;

 FSRNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSRNI =
  0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284 ;

 FSRVD =
  0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081 ;

 FSRVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSRVI =
  0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  1.095659e-14, 1.099812e-14, 1.099e-14, 1.102352e-14, 1.10049e-14, 
    1.102682e-14, 1.096491e-14, 1.099965e-14, 1.097744e-14, 1.096016e-14, 
    1.108844e-14, 1.102487e-14, 1.115442e-14, 1.111384e-14, 1.121569e-14, 
    1.114807e-14, 1.12293e-14, 1.121367e-14, 1.126058e-14, 1.124711e-14, 
    1.130714e-14, 1.126674e-14, 1.133822e-14, 1.129745e-14, 1.130381e-14, 
    1.126532e-14, 1.103777e-14, 1.108067e-14, 1.10352e-14, 1.104132e-14, 
    1.103855e-14, 1.100521e-14, 1.098843e-14, 1.095324e-14, 1.095959e-14, 
    1.098542e-14, 1.104393e-14, 1.102402e-14, 1.107408e-14, 1.107296e-14, 
    1.11287e-14, 1.110355e-14, 1.119731e-14, 1.117062e-14, 1.124765e-14, 
    1.122825e-14, 1.124671e-14, 1.124108e-14, 1.124673e-14, 1.121832e-14, 
    1.123045e-14, 1.120545e-14, 1.110848e-14, 1.113707e-14, 1.105174e-14, 
    1.100046e-14, 1.096636e-14, 1.09422e-14, 1.094558e-14, 1.095209e-14, 
    1.098554e-14, 1.101696e-14, 1.104094e-14, 1.105695e-14, 1.107274e-14, 
    1.112065e-14, 1.114595e-14, 1.120267e-14, 1.11924e-14, 1.120974e-14, 
    1.12263e-14, 1.125411e-14, 1.124952e-14, 1.126176e-14, 1.120917e-14, 
    1.124411e-14, 1.11864e-14, 1.120218e-14, 1.107728e-14, 1.102947e-14, 
    1.10092e-14, 1.09914e-14, 1.094819e-14, 1.097802e-14, 1.096624e-14, 
    1.099417e-14, 1.101194e-14, 1.100312e-14, 1.105737e-14, 1.103625e-14, 
    1.114742e-14, 1.109952e-14, 1.122439e-14, 1.119447e-14, 1.12315e-14, 
    1.121259e-14, 1.124496e-14, 1.12158e-14, 1.126628e-14, 1.12773e-14, 
    1.126973e-14, 1.129861e-14, 1.121407e-14, 1.124653e-14, 1.100298e-14, 
    1.100442e-14, 1.101107e-14, 1.098169e-14, 1.097989e-14, 1.095295e-14, 
    1.097687e-14, 1.098707e-14, 1.101292e-14, 1.10282e-14, 1.104273e-14, 
    1.107475e-14, 1.111049e-14, 1.116047e-14, 1.119638e-14, 1.122044e-14, 
    1.120566e-14, 1.121868e-14, 1.120409e-14, 1.119723e-14, 1.127312e-14, 
    1.12305e-14, 1.129441e-14, 1.129087e-14, 1.126191e-14, 1.129122e-14, 
    1.100539e-14, 1.09971e-14, 1.096846e-14, 1.099084e-14, 1.094999e-14, 
    1.097285e-14, 1.098598e-14, 1.103667e-14, 1.104778e-14, 1.105813e-14, 
    1.107852e-14, 1.11047e-14, 1.115068e-14, 1.119067e-14, 1.122719e-14, 
    1.122448e-14, 1.122542e-14, 1.123355e-14, 1.121333e-14, 1.123684e-14, 
    1.124077e-14, 1.123044e-14, 1.129034e-14, 1.127322e-14, 1.129072e-14, 
    1.127954e-14, 1.099977e-14, 1.101362e-14, 1.10061e-14, 1.102021e-14, 
    1.101024e-14, 1.105445e-14, 1.106768e-14, 1.112969e-14, 1.110419e-14, 
    1.114472e-14, 1.110826e-14, 1.111472e-14, 1.114601e-14, 1.111018e-14, 
    1.118842e-14, 1.113536e-14, 1.123385e-14, 1.118088e-14, 1.123713e-14, 
    1.122688e-14, 1.124378e-14, 1.125895e-14, 1.127798e-14, 1.131319e-14, 
    1.1305e-14, 1.133444e-14, 1.10343e-14, 1.105229e-14, 1.105069e-14, 
    1.106951e-14, 1.108344e-14, 1.111366e-14, 1.116213e-14, 1.114386e-14, 
    1.117731e-14, 1.118404e-14, 1.113314e-14, 1.116438e-14, 1.106416e-14, 
    1.108033e-14, 1.107067e-14, 1.103545e-14, 1.114792e-14, 1.109017e-14, 
    1.119676e-14, 1.116545e-14, 1.125673e-14, 1.121133e-14, 1.13005e-14, 
    1.133867e-14, 1.137452e-14, 1.141648e-14, 1.10621e-14, 1.104983e-14, 
    1.107172e-14, 1.110207e-14, 1.113015e-14, 1.116758e-14, 1.117138e-14, 
    1.117836e-14, 1.119649e-14, 1.121177e-14, 1.118055e-14, 1.121555e-14, 
    1.108408e-14, 1.115292e-14, 1.104497e-14, 1.107748e-14, 1.110001e-14, 
    1.10901e-14, 1.114153e-14, 1.115364e-14, 1.120293e-14, 1.117743e-14, 
    1.13292e-14, 1.126203e-14, 1.144838e-14, 1.139629e-14, 1.104553e-14, 
    1.106197e-14, 1.111931e-14, 1.109202e-14, 1.117002e-14, 1.118924e-14, 
    1.120482e-14, 1.12248e-14, 1.122691e-14, 1.123875e-14, 1.121931e-14, 
    1.123794e-14, 1.116746e-14, 1.119894e-14, 1.111254e-14, 1.113353e-14, 
    1.112385e-14, 1.111321e-14, 1.114593e-14, 1.118083e-14, 1.118154e-14, 
    1.11927e-14, 1.122428e-14, 1.116999e-14, 1.133784e-14, 1.123416e-14, 
    1.107992e-14, 1.111165e-14, 1.111614e-14, 1.110385e-14, 1.118726e-14, 
    1.115702e-14, 1.123846e-14, 1.121641e-14, 1.125246e-14, 1.123454e-14, 
    1.123186e-14, 1.120884e-14, 1.119447e-14, 1.115827e-14, 1.112877e-14, 
    1.110541e-14, 1.11108e-14, 1.113647e-14, 1.118291e-14, 1.122688e-14, 
    1.121723e-14, 1.124949e-14, 1.116398e-14, 1.119984e-14, 1.118594e-14, 
    1.122206e-14, 1.11433e-14, 1.121075e-14, 1.112605e-14, 1.113344e-14, 
    1.115637e-14, 1.120256e-14, 1.121271e-14, 1.122363e-14, 1.121685e-14, 
    1.118422e-14, 1.117885e-14, 1.115569e-14, 1.114928e-14, 1.113166e-14, 
    1.111703e-14, 1.113037e-14, 1.114433e-14, 1.118409e-14, 1.12199e-14, 
    1.125894e-14, 1.126849e-14, 1.131416e-14, 1.127697e-14, 1.133833e-14, 
    1.128617e-14, 1.13764e-14, 1.121458e-14, 1.128498e-14, 1.115741e-14, 
    1.117112e-14, 1.119597e-14, 1.125293e-14, 1.122212e-14, 1.125812e-14, 
    1.117862e-14, 1.11374e-14, 1.112669e-14, 1.110681e-14, 1.112711e-14, 
    1.112546e-14, 1.11449e-14, 1.113862e-14, 1.118535e-14, 1.116024e-14, 
    1.123156e-14, 1.125761e-14, 1.133115e-14, 1.137623e-14, 1.142212e-14, 
    1.144236e-14, 1.144852e-14, 1.145108e-14 ;

 F_DENIT_vr =
  6.256325e-13, 6.280041e-13, 6.275405e-13, 6.294542e-13, 6.28391e-13, 
    6.296427e-13, 6.261076e-13, 6.280915e-13, 6.268232e-13, 6.258365e-13, 
    6.331615e-13, 6.295313e-13, 6.369291e-13, 6.346117e-13, 6.404274e-13, 
    6.365665e-13, 6.412048e-13, 6.403123e-13, 6.42991e-13, 6.422217e-13, 
    6.456496e-13, 6.433425e-13, 6.474238e-13, 6.450962e-13, 6.454593e-13, 
    6.432614e-13, 6.302681e-13, 6.327176e-13, 6.301212e-13, 6.304706e-13, 
    6.303124e-13, 6.284089e-13, 6.274508e-13, 6.254411e-13, 6.25804e-13, 
    6.272788e-13, 6.306201e-13, 6.29483e-13, 6.323416e-13, 6.322772e-13, 
    6.354605e-13, 6.340244e-13, 6.39378e-13, 6.378539e-13, 6.422525e-13, 
    6.411446e-13, 6.421986e-13, 6.418771e-13, 6.421998e-13, 6.405775e-13, 
    6.412703e-13, 6.398427e-13, 6.343059e-13, 6.359382e-13, 6.310659e-13, 
    6.281375e-13, 6.261904e-13, 6.248109e-13, 6.250037e-13, 6.253759e-13, 
    6.272854e-13, 6.2908e-13, 6.304489e-13, 6.313636e-13, 6.322649e-13, 
    6.350007e-13, 6.364454e-13, 6.396839e-13, 6.390979e-13, 6.400877e-13, 
    6.410333e-13, 6.426213e-13, 6.423591e-13, 6.43058e-13, 6.400554e-13, 
    6.420505e-13, 6.387553e-13, 6.396562e-13, 6.325241e-13, 6.297939e-13, 
    6.286367e-13, 6.276202e-13, 6.25153e-13, 6.268562e-13, 6.261835e-13, 
    6.277784e-13, 6.28793e-13, 6.282893e-13, 6.313874e-13, 6.301811e-13, 
    6.365295e-13, 6.337942e-13, 6.409243e-13, 6.392156e-13, 6.413304e-13, 
    6.402506e-13, 6.420991e-13, 6.404336e-13, 6.433163e-13, 6.439452e-13, 
    6.435134e-13, 6.451626e-13, 6.403348e-13, 6.421885e-13, 6.282814e-13, 
    6.283636e-13, 6.287435e-13, 6.270661e-13, 6.269629e-13, 6.25425e-13, 
    6.267903e-13, 6.273729e-13, 6.288489e-13, 6.297218e-13, 6.305516e-13, 
    6.323796e-13, 6.344204e-13, 6.372742e-13, 6.393251e-13, 6.406989e-13, 
    6.398549e-13, 6.40598e-13, 6.397651e-13, 6.393732e-13, 6.437068e-13, 
    6.41273e-13, 6.449223e-13, 6.447204e-13, 6.430666e-13, 6.447401e-13, 
    6.28419e-13, 6.279461e-13, 6.263105e-13, 6.275885e-13, 6.252555e-13, 
    6.265612e-13, 6.273108e-13, 6.302056e-13, 6.308399e-13, 6.314307e-13, 
    6.325949e-13, 6.340899e-13, 6.367155e-13, 6.389987e-13, 6.410839e-13, 
    6.409294e-13, 6.409828e-13, 6.414475e-13, 6.402925e-13, 6.416349e-13, 
    6.418594e-13, 6.412695e-13, 6.446902e-13, 6.437125e-13, 6.447119e-13, 
    6.440733e-13, 6.28098e-13, 6.288893e-13, 6.284595e-13, 6.292656e-13, 
    6.286958e-13, 6.312205e-13, 6.319761e-13, 6.355166e-13, 6.340606e-13, 
    6.363751e-13, 6.342933e-13, 6.346622e-13, 6.364485e-13, 6.344027e-13, 
    6.3887e-13, 6.358404e-13, 6.414644e-13, 6.384397e-13, 6.416519e-13, 
    6.410663e-13, 6.420314e-13, 6.428977e-13, 6.439843e-13, 6.459949e-13, 
    6.455269e-13, 6.47208e-13, 6.300701e-13, 6.310974e-13, 6.310058e-13, 
    6.320807e-13, 6.328756e-13, 6.346014e-13, 6.373689e-13, 6.363258e-13, 
    6.382358e-13, 6.3862e-13, 6.357135e-13, 6.374974e-13, 6.317749e-13, 
    6.32698e-13, 6.321466e-13, 6.301355e-13, 6.365579e-13, 6.332599e-13, 
    6.393465e-13, 6.375585e-13, 6.427712e-13, 6.401788e-13, 6.4527e-13, 
    6.474497e-13, 6.494968e-13, 6.518927e-13, 6.316572e-13, 6.309564e-13, 
    6.322064e-13, 6.339394e-13, 6.355433e-13, 6.376802e-13, 6.378972e-13, 
    6.382961e-13, 6.393314e-13, 6.402037e-13, 6.384207e-13, 6.404192e-13, 
    6.329126e-13, 6.368435e-13, 6.306789e-13, 6.325355e-13, 6.338223e-13, 
    6.332564e-13, 6.36193e-13, 6.368842e-13, 6.396986e-13, 6.382428e-13, 
    6.469092e-13, 6.430737e-13, 6.537141e-13, 6.507401e-13, 6.307111e-13, 
    6.316501e-13, 6.349239e-13, 6.333656e-13, 6.378195e-13, 6.389172e-13, 
    6.398065e-13, 6.409477e-13, 6.410681e-13, 6.417443e-13, 6.406344e-13, 
    6.416982e-13, 6.376735e-13, 6.39471e-13, 6.345373e-13, 6.357363e-13, 
    6.351833e-13, 6.345761e-13, 6.36444e-13, 6.384372e-13, 6.384774e-13, 
    6.39115e-13, 6.409179e-13, 6.378182e-13, 6.474022e-13, 6.414824e-13, 
    6.326747e-13, 6.344867e-13, 6.347431e-13, 6.340411e-13, 6.388041e-13, 
    6.370776e-13, 6.417276e-13, 6.404685e-13, 6.425273e-13, 6.415038e-13, 
    6.41351e-13, 6.400363e-13, 6.392157e-13, 6.371486e-13, 6.354643e-13, 
    6.341304e-13, 6.344382e-13, 6.35904e-13, 6.385558e-13, 6.410666e-13, 
    6.405154e-13, 6.423575e-13, 6.374749e-13, 6.395222e-13, 6.38729e-13, 
    6.407914e-13, 6.36294e-13, 6.401456e-13, 6.35309e-13, 6.357311e-13, 
    6.370403e-13, 6.396776e-13, 6.402573e-13, 6.408808e-13, 6.404937e-13, 
    6.386308e-13, 6.383238e-13, 6.370012e-13, 6.366357e-13, 6.356293e-13, 
    6.347941e-13, 6.355556e-13, 6.363529e-13, 6.386229e-13, 6.406678e-13, 
    6.428971e-13, 6.434423e-13, 6.460503e-13, 6.439269e-13, 6.474301e-13, 
    6.444518e-13, 6.496041e-13, 6.403643e-13, 6.443839e-13, 6.370997e-13, 
    6.378823e-13, 6.393013e-13, 6.425538e-13, 6.407945e-13, 6.428502e-13, 
    6.38311e-13, 6.359568e-13, 6.353456e-13, 6.342102e-13, 6.353695e-13, 
    6.352752e-13, 6.363855e-13, 6.360266e-13, 6.386952e-13, 6.372611e-13, 
    6.413334e-13, 6.428212e-13, 6.470201e-13, 6.495943e-13, 6.522146e-13, 
    6.533706e-13, 6.537224e-13, 6.538685e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  3.319626e-16, 3.320568e-16, 3.320374e-16, 3.321117e-16, 3.320699e-16, 
    3.321174e-16, 3.319789e-16, 3.320569e-16, 3.320065e-16, 3.319661e-16, 
    3.322452e-16, 3.321105e-16, 3.323737e-16, 3.322936e-16, 3.324849e-16, 
    3.323604e-16, 3.325082e-16, 3.324794e-16, 3.325604e-16, 3.325367e-16, 
    3.326363e-16, 3.325694e-16, 3.326836e-16, 3.326194e-16, 3.326292e-16, 
    3.325646e-16, 3.321416e-16, 3.322331e-16, 3.321351e-16, 3.321485e-16, 
    3.321417e-16, 3.320687e-16, 3.320315e-16, 3.319498e-16, 3.319638e-16, 
    3.32023e-16, 3.321505e-16, 3.321066e-16, 3.322118e-16, 3.322096e-16, 
    3.323208e-16, 3.32271e-16, 3.324494e-16, 3.323993e-16, 3.325371e-16, 
    3.325027e-16, 3.325345e-16, 3.32524e-16, 3.325331e-16, 3.324837e-16, 
    3.325039e-16, 3.324596e-16, 3.32287e-16, 3.323425e-16, 3.321695e-16, 
    3.320585e-16, 3.319802e-16, 3.319242e-16, 3.31931e-16, 3.319464e-16, 
    3.320223e-16, 3.320908e-16, 3.321423e-16, 3.321754e-16, 3.322076e-16, 
    3.323057e-16, 3.323537e-16, 3.324582e-16, 3.32439e-16, 3.324699e-16, 
    3.324987e-16, 3.325461e-16, 3.325379e-16, 3.325581e-16, 3.324658e-16, 
    3.325275e-16, 3.324234e-16, 3.324524e-16, 3.322239e-16, 3.321206e-16, 
    3.320771e-16, 3.320362e-16, 3.319368e-16, 3.320056e-16, 3.319781e-16, 
    3.320401e-16, 3.320793e-16, 3.32059e-16, 3.321757e-16, 3.321302e-16, 
    3.323557e-16, 3.322614e-16, 3.32496e-16, 3.324416e-16, 3.32507e-16, 
    3.324736e-16, 3.325295e-16, 3.324784e-16, 3.325645e-16, 3.325832e-16, 
    3.325694e-16, 3.326168e-16, 3.324722e-16, 3.325293e-16, 3.320617e-16, 
    3.320651e-16, 3.32079e-16, 3.320131e-16, 3.320088e-16, 3.319461e-16, 
    3.320003e-16, 3.320236e-16, 3.320799e-16, 3.321125e-16, 3.321431e-16, 
    3.322103e-16, 3.322824e-16, 3.323786e-16, 3.324446e-16, 3.324868e-16, 
    3.324602e-16, 3.324826e-16, 3.324564e-16, 3.324431e-16, 3.325748e-16, 
    3.325021e-16, 3.326085e-16, 3.326028e-16, 3.325544e-16, 3.326019e-16, 
    3.320662e-16, 3.320469e-16, 3.319823e-16, 3.32032e-16, 3.319382e-16, 
    3.319911e-16, 3.320203e-16, 3.321308e-16, 3.321533e-16, 3.321754e-16, 
    3.32217e-16, 3.322694e-16, 3.323593e-16, 3.324332e-16, 3.324981e-16, 
    3.324925e-16, 3.324939e-16, 3.325075e-16, 3.324716e-16, 3.325122e-16, 
    3.325185e-16, 3.325005e-16, 3.326005e-16, 3.325724e-16, 3.326005e-16, 
    3.325813e-16, 3.320522e-16, 3.320821e-16, 3.320649e-16, 3.32096e-16, 
    3.320732e-16, 3.321687e-16, 3.321958e-16, 3.3232e-16, 3.322684e-16, 
    3.323483e-16, 3.322755e-16, 3.322886e-16, 3.323498e-16, 3.322778e-16, 
    3.324278e-16, 3.323272e-16, 3.325074e-16, 3.324125e-16, 3.325121e-16, 
    3.324933e-16, 3.32522e-16, 3.325482e-16, 3.325788e-16, 3.326363e-16, 
    3.326219e-16, 3.326683e-16, 3.321264e-16, 3.321642e-16, 3.321602e-16, 
    3.321989e-16, 3.32227e-16, 3.322879e-16, 3.323812e-16, 3.323454e-16, 
    3.324079e-16, 3.324206e-16, 3.323229e-16, 3.323832e-16, 3.321837e-16, 
    3.322168e-16, 3.321962e-16, 3.321212e-16, 3.323495e-16, 3.322348e-16, 
    3.324392e-16, 3.323805e-16, 3.32543e-16, 3.324644e-16, 3.326144e-16, 
    3.326752e-16, 3.327275e-16, 3.327872e-16, 3.32184e-16, 3.321572e-16, 
    3.322024e-16, 3.32265e-16, 3.32319e-16, 3.323907e-16, 3.32397e-16, 
    3.324093e-16, 3.324417e-16, 3.324694e-16, 3.324124e-16, 3.324746e-16, 
    3.322246e-16, 3.323587e-16, 3.321404e-16, 3.32209e-16, 3.322534e-16, 
    3.322333e-16, 3.323342e-16, 3.323566e-16, 3.324476e-16, 3.324008e-16, 
    3.326592e-16, 3.325501e-16, 3.328288e-16, 3.327578e-16, 3.321476e-16, 
    3.321814e-16, 3.322976e-16, 3.322429e-16, 3.323936e-16, 3.324294e-16, 
    3.324564e-16, 3.324924e-16, 3.324947e-16, 3.325156e-16, 3.324803e-16, 
    3.325131e-16, 3.32385e-16, 3.32443e-16, 3.322781e-16, 3.323188e-16, 
    3.322995e-16, 3.322777e-16, 3.323409e-16, 3.324073e-16, 3.324074e-16, 
    3.324273e-16, 3.324854e-16, 3.323841e-16, 3.326716e-16, 3.325007e-16, 
    3.32218e-16, 3.32282e-16, 3.322897e-16, 3.322652e-16, 3.324243e-16, 
    3.323681e-16, 3.32515e-16, 3.324754e-16, 3.325375e-16, 3.325068e-16, 
    3.32501e-16, 3.324604e-16, 3.324334e-16, 3.323665e-16, 3.323086e-16, 
    3.322622e-16, 3.322719e-16, 3.323227e-16, 3.324095e-16, 3.324886e-16, 
    3.32471e-16, 3.32526e-16, 3.323718e-16, 3.324384e-16, 3.32412e-16, 
    3.324769e-16, 3.323424e-16, 3.324692e-16, 3.323081e-16, 3.323218e-16, 
    3.323653e-16, 3.324514e-16, 3.324678e-16, 3.324876e-16, 3.324742e-16, 
    3.324157e-16, 3.324049e-16, 3.323605e-16, 3.323479e-16, 3.323137e-16, 
    3.322839e-16, 3.323103e-16, 3.323364e-16, 3.324111e-16, 3.324753e-16, 
    3.32542e-16, 3.325576e-16, 3.326324e-16, 3.325716e-16, 3.326699e-16, 
    3.325871e-16, 3.327254e-16, 3.324739e-16, 3.325945e-16, 3.323672e-16, 
    3.323922e-16, 3.324384e-16, 3.32538e-16, 3.324832e-16, 3.325461e-16, 
    3.324041e-16, 3.323256e-16, 3.323035e-16, 3.322644e-16, 3.323034e-16, 
    3.323002e-16, 3.323372e-16, 3.323243e-16, 3.32412e-16, 3.323651e-16, 
    3.324938e-16, 3.32539e-16, 3.326575e-16, 3.327249e-16, 3.327891e-16, 
    3.328157e-16, 3.328237e-16, 3.328265e-16 ;

 F_N2O_NIT =
  2.414584e-14, 2.435388e-14, 2.431336e-14, 2.448168e-14, 2.438823e-14, 
    2.449855e-14, 2.418793e-14, 2.436214e-14, 2.425085e-14, 2.416451e-14, 
    2.481004e-14, 2.448918e-14, 2.514558e-14, 2.493927e-14, 2.545918e-14, 
    2.511342e-14, 2.552919e-14, 2.544916e-14, 2.56904e-14, 2.562116e-14, 
    2.593103e-14, 2.572238e-14, 2.60924e-14, 2.588111e-14, 2.591411e-14, 
    2.57155e-14, 2.455359e-14, 2.477e-14, 2.45408e-14, 2.457159e-14, 
    2.455777e-14, 2.439015e-14, 2.430591e-14, 2.412995e-14, 2.416184e-14, 
    2.42911e-14, 2.458542e-14, 2.44853e-14, 2.473802e-14, 2.473229e-14, 
    2.501519e-14, 2.488743e-14, 2.53654e-14, 2.522907e-14, 2.562405e-14, 
    2.552441e-14, 2.561936e-14, 2.559054e-14, 2.561973e-14, 2.547369e-14, 
    2.55362e-14, 2.540789e-14, 2.491136e-14, 2.505678e-14, 2.462437e-14, 
    2.436624e-14, 2.419555e-14, 2.407481e-14, 2.409185e-14, 2.412438e-14, 
    2.429185e-14, 2.444985e-14, 2.457061e-14, 2.465157e-14, 2.473146e-14, 
    2.497415e-14, 2.510308e-14, 2.539301e-14, 2.534055e-14, 2.542944e-14, 
    2.551451e-14, 2.565766e-14, 2.563407e-14, 2.569724e-14, 2.542708e-14, 
    2.560646e-14, 2.531067e-14, 2.53914e-14, 2.475326e-14, 2.45123e-14, 
    2.441027e-14, 2.432112e-14, 2.410497e-14, 2.425413e-14, 2.419527e-14, 
    2.433541e-14, 2.442468e-14, 2.43805e-14, 2.465378e-14, 2.454734e-14, 
    2.511072e-14, 2.486725e-14, 2.550458e-14, 2.53513e-14, 2.554138e-14, 
    2.54443e-14, 2.561076e-14, 2.546091e-14, 2.572077e-14, 2.577754e-14, 
    2.573873e-14, 2.588793e-14, 2.54526e-14, 2.561933e-14, 2.437928e-14, 
    2.438648e-14, 2.442004e-14, 2.427268e-14, 2.426368e-14, 2.412906e-14, 
    2.424882e-14, 2.429991e-14, 2.442985e-14, 2.450688e-14, 2.458022e-14, 
    2.474187e-14, 2.492306e-14, 2.517756e-14, 2.536122e-14, 2.548472e-14, 
    2.540895e-14, 2.547584e-14, 2.540107e-14, 2.536606e-14, 2.575625e-14, 
    2.553677e-14, 2.586643e-14, 2.584814e-14, 2.569872e-14, 2.585019e-14, 
    2.439153e-14, 2.43501e-14, 2.420654e-14, 2.431885e-14, 2.411442e-14, 
    2.422874e-14, 2.42946e-14, 2.454957e-14, 2.460576e-14, 2.465794e-14, 
    2.476115e-14, 2.489394e-14, 2.512777e-14, 2.533214e-14, 2.551945e-14, 
    2.55057e-14, 2.551054e-14, 2.555247e-14, 2.544866e-14, 2.556953e-14, 
    2.558984e-14, 2.553674e-14, 2.584568e-14, 2.575722e-14, 2.584774e-14, 
    2.579011e-14, 2.436356e-14, 2.443331e-14, 2.43956e-14, 2.446653e-14, 
    2.441654e-14, 2.463918e-14, 2.470614e-14, 2.502067e-14, 2.489132e-14, 
    2.509733e-14, 2.49122e-14, 2.494496e-14, 2.510407e-14, 2.492218e-14, 
    2.532085e-14, 2.505021e-14, 2.55541e-14, 2.528256e-14, 2.557116e-14, 
    2.551862e-14, 2.560562e-14, 2.568369e-14, 2.578205e-14, 2.596409e-14, 
    2.592187e-14, 2.607448e-14, 2.453748e-14, 2.46283e-14, 2.462029e-14, 
    2.471551e-14, 2.478605e-14, 2.493929e-14, 2.51861e-14, 2.509314e-14, 
    2.526393e-14, 2.529829e-14, 2.503886e-14, 2.519798e-14, 2.468916e-14, 
    2.4771e-14, 2.472225e-14, 2.45446e-14, 2.511453e-14, 2.482119e-14, 
    2.536423e-14, 2.520429e-14, 2.567254e-14, 2.543911e-14, 2.589865e-14, 
    2.609641e-14, 2.628322e-14, 2.650243e-14, 2.467794e-14, 2.461614e-14, 
    2.472684e-14, 2.488043e-14, 2.502337e-14, 2.521406e-14, 2.523361e-14, 
    2.526943e-14, 2.536233e-14, 2.544059e-14, 2.528076e-14, 2.546021e-14, 
    2.479001e-14, 2.514007e-14, 2.459276e-14, 2.475692e-14, 2.487133e-14, 
    2.48211e-14, 2.508249e-14, 2.51443e-14, 2.53963e-14, 2.526587e-14, 
    2.604753e-14, 2.570018e-14, 2.666996e-14, 2.639708e-14, 2.459456e-14, 
    2.467771e-14, 2.496825e-14, 2.482979e-14, 2.522681e-14, 2.532503e-14, 
    2.540502e-14, 2.550747e-14, 2.551854e-14, 2.557935e-14, 2.547973e-14, 
    2.557541e-14, 2.521444e-14, 2.537542e-14, 2.493492e-14, 2.504176e-14, 
    2.499258e-14, 2.493868e-14, 2.51052e-14, 2.528324e-14, 2.528704e-14, 
    2.534427e-14, 2.550592e-14, 2.522837e-14, 2.609254e-14, 2.555708e-14, 
    2.476855e-14, 2.492944e-14, 2.495245e-14, 2.489003e-14, 2.531517e-14, 
    2.51607e-14, 2.557787e-14, 2.546477e-14, 2.565021e-14, 2.555797e-14, 
    2.554441e-14, 2.542623e-14, 2.535279e-14, 2.516775e-14, 2.50177e-14, 
    2.489905e-14, 2.492661e-14, 2.505704e-14, 2.529414e-14, 2.551951e-14, 
    2.547005e-14, 2.563606e-14, 2.519785e-14, 2.538113e-14, 2.531021e-14, 
    2.549533e-14, 2.509066e-14, 2.543512e-14, 2.5003e-14, 2.504073e-14, 
    2.515763e-14, 2.539363e-14, 2.544598e-14, 2.550196e-14, 2.54674e-14, 
    2.530019e-14, 2.527285e-14, 2.515476e-14, 2.512221e-14, 2.503249e-14, 
    2.495833e-14, 2.502608e-14, 2.509733e-14, 2.530024e-14, 2.548383e-14, 
    2.568477e-14, 2.573406e-14, 2.597013e-14, 2.577788e-14, 2.609552e-14, 
    2.582535e-14, 2.629394e-14, 2.545513e-14, 2.581747e-14, 2.516295e-14, 
    2.523304e-14, 2.536008e-14, 2.565269e-14, 2.549449e-14, 2.567954e-14, 
    2.527178e-14, 2.506155e-14, 2.500729e-14, 2.490625e-14, 2.50096e-14, 
    2.500119e-14, 2.510027e-14, 2.50684e-14, 2.530698e-14, 2.517868e-14, 
    2.554404e-14, 2.567805e-14, 2.605844e-14, 2.629307e-14, 2.653301e-14, 
    2.66393e-14, 2.66717e-14, 2.668524e-14 ;

 F_NIT =
  4.024307e-11, 4.05898e-11, 4.052226e-11, 4.080281e-11, 4.064705e-11, 
    4.083092e-11, 4.031322e-11, 4.060357e-11, 4.041808e-11, 4.027418e-11, 
    4.135007e-11, 4.081531e-11, 4.19093e-11, 4.156545e-11, 4.243196e-11, 
    4.18557e-11, 4.254865e-11, 4.241526e-11, 4.281734e-11, 4.270194e-11, 
    4.321838e-11, 4.287063e-11, 4.348734e-11, 4.313519e-11, 4.319018e-11, 
    4.285917e-11, 4.092265e-11, 4.128333e-11, 4.090133e-11, 4.095265e-11, 
    4.092961e-11, 4.065025e-11, 4.050985e-11, 4.021659e-11, 4.026974e-11, 
    4.048516e-11, 4.09757e-11, 4.080883e-11, 4.123003e-11, 4.122049e-11, 
    4.169198e-11, 4.147905e-11, 4.227567e-11, 4.204844e-11, 4.270675e-11, 
    4.254069e-11, 4.269893e-11, 4.265091e-11, 4.269955e-11, 4.245615e-11, 
    4.256033e-11, 4.234648e-11, 4.151894e-11, 4.17613e-11, 4.104061e-11, 
    4.06104e-11, 4.032591e-11, 4.012468e-11, 4.015309e-11, 4.020729e-11, 
    4.048642e-11, 4.074975e-11, 4.095102e-11, 4.108594e-11, 4.12191e-11, 
    4.162358e-11, 4.183846e-11, 4.232168e-11, 4.223425e-11, 4.23824e-11, 
    4.252418e-11, 4.276277e-11, 4.272345e-11, 4.282874e-11, 4.237846e-11, 
    4.267744e-11, 4.218445e-11, 4.2319e-11, 4.125543e-11, 4.085383e-11, 
    4.068378e-11, 4.05352e-11, 4.017494e-11, 4.042355e-11, 4.032545e-11, 
    4.055901e-11, 4.070779e-11, 4.063417e-11, 4.108963e-11, 4.091224e-11, 
    4.18512e-11, 4.144541e-11, 4.250764e-11, 4.225217e-11, 4.256897e-11, 
    4.240716e-11, 4.26846e-11, 4.243486e-11, 4.286795e-11, 4.296256e-11, 
    4.289788e-11, 4.314655e-11, 4.242101e-11, 4.269889e-11, 4.063213e-11, 
    4.064414e-11, 4.070007e-11, 4.045447e-11, 4.043947e-11, 4.021511e-11, 
    4.04147e-11, 4.049985e-11, 4.071641e-11, 4.08448e-11, 4.096703e-11, 
    4.123646e-11, 4.153843e-11, 4.19626e-11, 4.226871e-11, 4.247454e-11, 
    4.234825e-11, 4.245973e-11, 4.233511e-11, 4.227677e-11, 4.292709e-11, 
    4.256129e-11, 4.311072e-11, 4.308023e-11, 4.283121e-11, 4.308365e-11, 
    4.065255e-11, 4.05835e-11, 4.034424e-11, 4.053141e-11, 4.01907e-11, 
    4.038123e-11, 4.049099e-11, 4.091595e-11, 4.100961e-11, 4.109657e-11, 
    4.126859e-11, 4.14899e-11, 4.187962e-11, 4.222023e-11, 4.253242e-11, 
    4.25095e-11, 4.251756e-11, 4.258745e-11, 4.241443e-11, 4.261588e-11, 
    4.264973e-11, 4.256123e-11, 4.307613e-11, 4.29287e-11, 4.307956e-11, 
    4.298352e-11, 4.060593e-11, 4.072218e-11, 4.065933e-11, 4.077754e-11, 
    4.069424e-11, 4.106531e-11, 4.117689e-11, 4.170111e-11, 4.148554e-11, 
    4.182888e-11, 4.152034e-11, 4.157492e-11, 4.184011e-11, 4.153696e-11, 
    4.220141e-11, 4.175035e-11, 4.259016e-11, 4.21376e-11, 4.26186e-11, 
    4.253103e-11, 4.267604e-11, 4.280614e-11, 4.297009e-11, 4.327349e-11, 
    4.320312e-11, 4.345747e-11, 4.08958e-11, 4.104717e-11, 4.103382e-11, 
    4.119251e-11, 4.131008e-11, 4.156549e-11, 4.197684e-11, 4.18219e-11, 
    4.210655e-11, 4.216381e-11, 4.173143e-11, 4.199664e-11, 4.114859e-11, 
    4.1285e-11, 4.120375e-11, 4.090767e-11, 4.185755e-11, 4.136866e-11, 
    4.227372e-11, 4.200714e-11, 4.278757e-11, 4.239853e-11, 4.316442e-11, 
    4.349402e-11, 4.380537e-11, 4.417072e-11, 4.11299e-11, 4.102689e-11, 
    4.12114e-11, 4.146739e-11, 4.170561e-11, 4.202343e-11, 4.205601e-11, 
    4.211571e-11, 4.227055e-11, 4.240098e-11, 4.213459e-11, 4.243369e-11, 
    4.131668e-11, 4.190012e-11, 4.098794e-11, 4.126154e-11, 4.145221e-11, 
    4.13685e-11, 4.180415e-11, 4.190717e-11, 4.232717e-11, 4.210978e-11, 
    4.341254e-11, 4.283363e-11, 4.444993e-11, 4.399513e-11, 4.099094e-11, 
    4.112952e-11, 4.161375e-11, 4.138299e-11, 4.204468e-11, 4.220839e-11, 
    4.23417e-11, 4.251246e-11, 4.25309e-11, 4.263226e-11, 4.246622e-11, 
    4.262568e-11, 4.202406e-11, 4.229236e-11, 4.15582e-11, 4.173627e-11, 
    4.165429e-11, 4.156447e-11, 4.1842e-11, 4.213873e-11, 4.214506e-11, 
    4.224044e-11, 4.250986e-11, 4.204729e-11, 4.348756e-11, 4.259513e-11, 
    4.128092e-11, 4.154906e-11, 4.158742e-11, 4.148339e-11, 4.219195e-11, 
    4.193449e-11, 4.262979e-11, 4.244128e-11, 4.275035e-11, 4.259662e-11, 
    4.257402e-11, 4.237705e-11, 4.225464e-11, 4.194625e-11, 4.169617e-11, 
    4.149842e-11, 4.154434e-11, 4.176173e-11, 4.21569e-11, 4.253252e-11, 
    4.245009e-11, 4.272676e-11, 4.199643e-11, 4.230188e-11, 4.218368e-11, 
    4.249221e-11, 4.181777e-11, 4.239186e-11, 4.167167e-11, 4.173455e-11, 
    4.192938e-11, 4.232271e-11, 4.240996e-11, 4.250326e-11, 4.244567e-11, 
    4.216699e-11, 4.212141e-11, 4.192461e-11, 4.187035e-11, 4.172082e-11, 
    4.159722e-11, 4.171013e-11, 4.182888e-11, 4.216706e-11, 4.247305e-11, 
    4.280794e-11, 4.28901e-11, 4.328354e-11, 4.296314e-11, 4.349254e-11, 
    4.304225e-11, 4.382324e-11, 4.242522e-11, 4.302911e-11, 4.193825e-11, 
    4.205507e-11, 4.22668e-11, 4.275448e-11, 4.249082e-11, 4.279924e-11, 
    4.211963e-11, 4.176925e-11, 4.167882e-11, 4.151042e-11, 4.168267e-11, 
    4.166864e-11, 4.183379e-11, 4.178068e-11, 4.217831e-11, 4.196447e-11, 
    4.257339e-11, 4.279674e-11, 4.343073e-11, 4.382178e-11, 4.422169e-11, 
    4.439884e-11, 4.445283e-11, 4.447541e-11 ;

 F_NIT_vr =
  2.396062e-10, 2.406568e-10, 2.404519e-10, 2.412998e-10, 2.408291e-10, 
    2.41384e-10, 2.398179e-10, 2.406968e-10, 2.401353e-10, 2.396986e-10, 
    2.429449e-10, 2.413357e-10, 2.446185e-10, 2.435901e-10, 2.461737e-10, 
    2.444578e-10, 2.465197e-10, 2.461235e-10, 2.473151e-10, 2.469732e-10, 
    2.484984e-10, 2.474721e-10, 2.492894e-10, 2.482528e-10, 2.484146e-10, 
    2.47437e-10, 2.416611e-10, 2.427464e-10, 2.415964e-10, 2.417511e-10, 
    2.416813e-10, 2.408377e-10, 2.40413e-10, 2.395237e-10, 2.396846e-10, 
    2.403376e-10, 2.418188e-10, 2.413153e-10, 2.425834e-10, 2.425548e-10, 
    2.439678e-10, 2.433303e-10, 2.457083e-10, 2.450316e-10, 2.469872e-10, 
    2.464946e-10, 2.469636e-10, 2.468209e-10, 2.469647e-10, 2.46243e-10, 
    2.465516e-10, 2.459168e-10, 2.434527e-10, 2.441777e-10, 2.420155e-10, 
    2.407171e-10, 2.398553e-10, 2.392445e-10, 2.393303e-10, 2.39495e-10, 
    2.403409e-10, 2.411368e-10, 2.417438e-10, 2.421497e-10, 2.425499e-10, 
    2.437631e-10, 2.444052e-10, 2.458446e-10, 2.455845e-10, 2.460246e-10, 
    2.464454e-10, 2.47152e-10, 2.470355e-10, 2.473467e-10, 2.460116e-10, 
    2.468986e-10, 2.454342e-10, 2.458345e-10, 2.426614e-10, 2.414521e-10, 
    2.409386e-10, 2.40489e-10, 2.393965e-10, 2.401507e-10, 2.39853e-10, 
    2.405601e-10, 2.410098e-10, 2.407869e-10, 2.421606e-10, 2.416259e-10, 
    2.444429e-10, 2.432287e-10, 2.463966e-10, 2.456373e-10, 2.465779e-10, 
    2.460977e-10, 2.469201e-10, 2.461795e-10, 2.474622e-10, 2.477418e-10, 
    2.475502e-10, 2.482844e-10, 2.461369e-10, 2.46961e-10, 2.407822e-10, 
    2.408185e-10, 2.409872e-10, 2.40244e-10, 2.401984e-10, 2.395177e-10, 
    2.401227e-10, 2.403807e-10, 2.410352e-10, 2.414224e-10, 2.417906e-10, 
    2.426013e-10, 2.43507e-10, 2.447746e-10, 2.456862e-10, 2.462974e-10, 
    2.459222e-10, 2.462529e-10, 2.458827e-10, 2.457088e-10, 2.476363e-10, 
    2.465535e-10, 2.48178e-10, 2.480881e-10, 2.473521e-10, 2.480975e-10, 
    2.408435e-10, 2.406343e-10, 2.399097e-10, 2.404763e-10, 2.394431e-10, 
    2.400212e-10, 2.403533e-10, 2.416367e-10, 2.419187e-10, 2.421805e-10, 
    2.426974e-10, 2.43361e-10, 2.445267e-10, 2.455414e-10, 2.464688e-10, 
    2.464005e-10, 2.464243e-10, 2.466312e-10, 2.461177e-10, 2.46715e-10, 
    2.46815e-10, 2.465527e-10, 2.480753e-10, 2.4764e-10, 2.480852e-10, 
    2.478013e-10, 2.407019e-10, 2.410528e-10, 2.408627e-10, 2.412198e-10, 
    2.409677e-10, 2.420867e-10, 2.424221e-10, 2.439937e-10, 2.433479e-10, 
    2.443754e-10, 2.434517e-10, 2.436153e-10, 2.44408e-10, 2.435009e-10, 
    2.454847e-10, 2.44139e-10, 2.46639e-10, 2.45294e-10, 2.467228e-10, 
    2.464627e-10, 2.468923e-10, 2.472775e-10, 2.477616e-10, 2.486565e-10, 
    2.484486e-10, 2.491973e-10, 2.415765e-10, 2.420322e-10, 2.419919e-10, 
    2.42469e-10, 2.428219e-10, 2.435878e-10, 2.44817e-10, 2.443541e-10, 
    2.452029e-10, 2.453734e-10, 2.440829e-10, 2.448749e-10, 2.423349e-10, 
    2.427445e-10, 2.425003e-10, 2.416086e-10, 2.444586e-10, 2.429947e-10, 
    2.456982e-10, 2.449041e-10, 2.472218e-10, 2.460685e-10, 2.483344e-10, 
    2.493045e-10, 2.502178e-10, 2.512858e-10, 2.422809e-10, 2.419705e-10, 
    2.425252e-10, 2.432937e-10, 2.440065e-10, 2.449556e-10, 2.450524e-10, 
    2.452299e-10, 2.456903e-10, 2.46078e-10, 2.452855e-10, 2.461745e-10, 
    2.428393e-10, 2.445856e-10, 2.4185e-10, 2.426731e-10, 2.432448e-10, 
    2.429938e-10, 2.442979e-10, 2.446052e-10, 2.458558e-10, 2.452091e-10, 
    2.490643e-10, 2.47357e-10, 2.520994e-10, 2.507723e-10, 2.418619e-10, 
    2.422788e-10, 2.437315e-10, 2.430399e-10, 2.450182e-10, 2.455058e-10, 
    2.459017e-10, 2.464088e-10, 2.46463e-10, 2.467636e-10, 2.462706e-10, 
    2.467436e-10, 2.449549e-10, 2.457536e-10, 2.435625e-10, 2.44095e-10, 
    2.438497e-10, 2.435804e-10, 2.444102e-10, 2.45295e-10, 2.453136e-10, 
    2.455971e-10, 2.463973e-10, 2.450216e-10, 2.492839e-10, 2.466494e-10, 
    2.427335e-10, 2.435374e-10, 2.43652e-10, 2.433404e-10, 2.454561e-10, 
    2.44689e-10, 2.467562e-10, 2.461967e-10, 2.471126e-10, 2.466573e-10, 
    2.465897e-10, 2.460052e-10, 2.456408e-10, 2.447222e-10, 2.439746e-10, 
    2.433826e-10, 2.435197e-10, 2.441702e-10, 2.453484e-10, 2.464648e-10, 
    2.462199e-10, 2.470397e-10, 2.448694e-10, 2.457789e-10, 2.454267e-10, 
    2.463438e-10, 2.443408e-10, 2.460509e-10, 2.439038e-10, 2.440914e-10, 
    2.446731e-10, 2.458445e-10, 2.461032e-10, 2.463802e-10, 2.462087e-10, 
    2.453803e-10, 2.452444e-10, 2.446572e-10, 2.44495e-10, 2.440482e-10, 
    2.436779e-10, 2.440158e-10, 2.443701e-10, 2.453786e-10, 2.462878e-10, 
    2.472798e-10, 2.475227e-10, 2.48683e-10, 2.47738e-10, 2.492973e-10, 
    2.47971e-10, 2.502671e-10, 2.461492e-10, 2.479373e-10, 2.446996e-10, 
    2.450476e-10, 2.456777e-10, 2.471243e-10, 2.463426e-10, 2.472565e-10, 
    2.452389e-10, 2.441931e-10, 2.439224e-10, 2.434182e-10, 2.439334e-10, 
    2.438915e-10, 2.443849e-10, 2.442258e-10, 2.454114e-10, 2.447743e-10, 
    2.465847e-10, 2.472463e-10, 2.491159e-10, 2.502631e-10, 2.514322e-10, 
    2.519483e-10, 2.521054e-10, 2.521708e-10,
  1.336014e-10, 1.346103e-10, 1.34414e-10, 1.352293e-10, 1.347768e-10, 
    1.35311e-10, 1.338058e-10, 1.346504e-10, 1.34111e-10, 1.336922e-10, 
    1.368166e-10, 1.352657e-10, 1.384346e-10, 1.374404e-10, 1.399427e-10, 
    1.382797e-10, 1.402789e-10, 1.398946e-10, 1.410523e-10, 1.407203e-10, 
    1.422048e-10, 1.412057e-10, 1.429765e-10, 1.41966e-10, 1.421239e-10, 
    1.411727e-10, 1.355773e-10, 1.366232e-10, 1.355154e-10, 1.356644e-10, 
    1.355975e-10, 1.347861e-10, 1.343779e-10, 1.335245e-10, 1.336793e-10, 
    1.343061e-10, 1.357314e-10, 1.35247e-10, 1.36469e-10, 1.364414e-10, 
    1.378065e-10, 1.371904e-10, 1.394922e-10, 1.388366e-10, 1.407342e-10, 
    1.402561e-10, 1.407117e-10, 1.405735e-10, 1.407135e-10, 1.400125e-10, 
    1.403127e-10, 1.396965e-10, 1.373057e-10, 1.380068e-10, 1.359196e-10, 
    1.346702e-10, 1.338428e-10, 1.332567e-10, 1.333395e-10, 1.334974e-10, 
    1.343098e-10, 1.350754e-10, 1.356598e-10, 1.360513e-10, 1.364374e-10, 
    1.376085e-10, 1.382299e-10, 1.396249e-10, 1.393728e-10, 1.398e-10, 
    1.402085e-10, 1.408954e-10, 1.407823e-10, 1.410852e-10, 1.397887e-10, 
    1.406499e-10, 1.392292e-10, 1.396173e-10, 1.365424e-10, 1.353776e-10, 
    1.348835e-10, 1.344517e-10, 1.334032e-10, 1.341269e-10, 1.338415e-10, 
    1.34521e-10, 1.349535e-10, 1.347395e-10, 1.36062e-10, 1.355473e-10, 
    1.382668e-10, 1.37093e-10, 1.401609e-10, 1.394245e-10, 1.403376e-10, 
    1.398714e-10, 1.406705e-10, 1.399512e-10, 1.41198e-10, 1.4147e-10, 
    1.412841e-10, 1.419987e-10, 1.399114e-10, 1.407117e-10, 1.347335e-10, 
    1.347684e-10, 1.34931e-10, 1.342169e-10, 1.341733e-10, 1.335202e-10, 
    1.341013e-10, 1.34349e-10, 1.349786e-10, 1.353515e-10, 1.357063e-10, 
    1.364877e-10, 1.373623e-10, 1.385887e-10, 1.394722e-10, 1.400656e-10, 
    1.397016e-10, 1.400229e-10, 1.396638e-10, 1.394955e-10, 1.413681e-10, 
    1.403155e-10, 1.418959e-10, 1.418083e-10, 1.410924e-10, 1.418181e-10, 
    1.347929e-10, 1.345922e-10, 1.338962e-10, 1.344408e-10, 1.334492e-10, 
    1.340039e-10, 1.343232e-10, 1.35558e-10, 1.358299e-10, 1.360821e-10, 
    1.365809e-10, 1.372219e-10, 1.38349e-10, 1.393324e-10, 1.402323e-10, 
    1.401663e-10, 1.401896e-10, 1.403909e-10, 1.398924e-10, 1.404727e-10, 
    1.405702e-10, 1.403154e-10, 1.417965e-10, 1.413728e-10, 1.418064e-10, 
    1.415305e-10, 1.346574e-10, 1.349953e-10, 1.348127e-10, 1.351561e-10, 
    1.349141e-10, 1.359914e-10, 1.36315e-10, 1.378329e-10, 1.372093e-10, 
    1.382024e-10, 1.3731e-10, 1.37468e-10, 1.382348e-10, 1.373582e-10, 
    1.392781e-10, 1.379754e-10, 1.403987e-10, 1.39094e-10, 1.404806e-10, 
    1.402284e-10, 1.40646e-10, 1.410204e-10, 1.414918e-10, 1.423632e-10, 
    1.421613e-10, 1.428911e-10, 1.354995e-10, 1.359388e-10, 1.359001e-10, 
    1.363604e-10, 1.367011e-10, 1.374407e-10, 1.386299e-10, 1.381822e-10, 
    1.390044e-10, 1.391696e-10, 1.379208e-10, 1.386871e-10, 1.362331e-10, 
    1.366285e-10, 1.36393e-10, 1.355342e-10, 1.382853e-10, 1.368709e-10, 
    1.394868e-10, 1.387176e-10, 1.40967e-10, 1.398466e-10, 1.420501e-10, 
    1.429958e-10, 1.438879e-10, 1.449329e-10, 1.361788e-10, 1.358801e-10, 
    1.364151e-10, 1.371567e-10, 1.37846e-10, 1.387644e-10, 1.388585e-10, 
    1.390309e-10, 1.394776e-10, 1.398536e-10, 1.390854e-10, 1.39948e-10, 
    1.367202e-10, 1.384084e-10, 1.357672e-10, 1.365605e-10, 1.371129e-10, 
    1.368705e-10, 1.381311e-10, 1.384288e-10, 1.39641e-10, 1.390139e-10, 
    1.427622e-10, 1.410995e-10, 1.457303e-10, 1.444309e-10, 1.357758e-10, 
    1.361778e-10, 1.375803e-10, 1.369123e-10, 1.388258e-10, 1.392983e-10, 
    1.396828e-10, 1.401748e-10, 1.40228e-10, 1.405199e-10, 1.400417e-10, 
    1.40501e-10, 1.387664e-10, 1.395406e-10, 1.374198e-10, 1.379349e-10, 
    1.376978e-10, 1.37438e-10, 1.382405e-10, 1.390974e-10, 1.391158e-10, 
    1.393909e-10, 1.401673e-10, 1.388336e-10, 1.429772e-10, 1.40413e-10, 
    1.366167e-10, 1.373931e-10, 1.375042e-10, 1.372031e-10, 1.392509e-10, 
    1.385076e-10, 1.405128e-10, 1.399698e-10, 1.408599e-10, 1.404173e-10, 
    1.403523e-10, 1.397848e-10, 1.394318e-10, 1.385417e-10, 1.378189e-10, 
    1.372468e-10, 1.373797e-10, 1.380085e-10, 1.391499e-10, 1.402328e-10, 
    1.399953e-10, 1.407921e-10, 1.386868e-10, 1.395682e-10, 1.392272e-10, 
    1.401168e-10, 1.381704e-10, 1.398272e-10, 1.37748e-10, 1.379298e-10, 
    1.384929e-10, 1.39628e-10, 1.398796e-10, 1.401484e-10, 1.399826e-10, 
    1.391789e-10, 1.390475e-10, 1.384792e-10, 1.383225e-10, 1.378902e-10, 
    1.375327e-10, 1.378593e-10, 1.382026e-10, 1.391793e-10, 1.400615e-10, 
    1.410257e-10, 1.41262e-10, 1.423921e-10, 1.414719e-10, 1.429916e-10, 
    1.416991e-10, 1.439391e-10, 1.399234e-10, 1.416612e-10, 1.385186e-10, 
    1.388559e-10, 1.394668e-10, 1.408717e-10, 1.401126e-10, 1.410005e-10, 
    1.390423e-10, 1.380302e-10, 1.377688e-10, 1.372815e-10, 1.3778e-10, 
    1.377394e-10, 1.382169e-10, 1.380634e-10, 1.392117e-10, 1.385945e-10, 
    1.403506e-10, 1.409935e-10, 1.428146e-10, 1.43935e-10, 1.450787e-10, 
    1.455846e-10, 1.457387e-10, 1.458032e-10,
  1.249146e-10, 1.260187e-10, 1.258037e-10, 1.266966e-10, 1.26201e-10, 
    1.267861e-10, 1.251382e-10, 1.260626e-10, 1.254721e-10, 1.250139e-10, 
    1.284367e-10, 1.267365e-10, 1.302131e-10, 1.291213e-10, 1.318713e-10, 
    1.300429e-10, 1.322413e-10, 1.318185e-10, 1.330929e-10, 1.327272e-10, 
    1.343628e-10, 1.332617e-10, 1.352139e-10, 1.340995e-10, 1.342736e-10, 
    1.332255e-10, 1.270779e-10, 1.282245e-10, 1.270101e-10, 1.271733e-10, 
    1.271001e-10, 1.262112e-10, 1.257642e-10, 1.248305e-10, 1.249998e-10, 
    1.256857e-10, 1.272467e-10, 1.267159e-10, 1.280555e-10, 1.280252e-10, 
    1.295233e-10, 1.288469e-10, 1.313758e-10, 1.306549e-10, 1.327425e-10, 
    1.322162e-10, 1.327178e-10, 1.325656e-10, 1.327197e-10, 1.319482e-10, 
    1.322785e-10, 1.316005e-10, 1.289734e-10, 1.297432e-10, 1.274531e-10, 
    1.260843e-10, 1.251786e-10, 1.245377e-10, 1.246282e-10, 1.248009e-10, 
    1.256898e-10, 1.26528e-10, 1.271683e-10, 1.275974e-10, 1.280208e-10, 
    1.293059e-10, 1.299883e-10, 1.315217e-10, 1.312445e-10, 1.317143e-10, 
    1.321639e-10, 1.329201e-10, 1.327955e-10, 1.331291e-10, 1.317019e-10, 
    1.326497e-10, 1.310866e-10, 1.315134e-10, 1.281359e-10, 1.26859e-10, 
    1.263179e-10, 1.25845e-10, 1.246978e-10, 1.254896e-10, 1.251772e-10, 
    1.259209e-10, 1.263945e-10, 1.261602e-10, 1.276091e-10, 1.27045e-10, 
    1.300288e-10, 1.2874e-10, 1.321114e-10, 1.313013e-10, 1.323059e-10, 
    1.317929e-10, 1.326724e-10, 1.318808e-10, 1.332533e-10, 1.33553e-10, 
    1.333482e-10, 1.341356e-10, 1.318369e-10, 1.327177e-10, 1.261536e-10, 
    1.261918e-10, 1.263698e-10, 1.255881e-10, 1.255403e-10, 1.248258e-10, 
    1.254615e-10, 1.257326e-10, 1.26422e-10, 1.268304e-10, 1.272193e-10, 
    1.28076e-10, 1.290356e-10, 1.303825e-10, 1.313538e-10, 1.320066e-10, 
    1.316061e-10, 1.319596e-10, 1.315645e-10, 1.313795e-10, 1.334407e-10, 
    1.322816e-10, 1.340223e-10, 1.339257e-10, 1.33137e-10, 1.339366e-10, 
    1.262186e-10, 1.259989e-10, 1.252371e-10, 1.258331e-10, 1.247481e-10, 
    1.253549e-10, 1.257044e-10, 1.270568e-10, 1.273547e-10, 1.276313e-10, 
    1.281782e-10, 1.288815e-10, 1.301191e-10, 1.312e-10, 1.321901e-10, 
    1.321174e-10, 1.32143e-10, 1.323645e-10, 1.31816e-10, 1.324547e-10, 
    1.32562e-10, 1.322815e-10, 1.339128e-10, 1.334459e-10, 1.339236e-10, 
    1.336196e-10, 1.260703e-10, 1.264403e-10, 1.262403e-10, 1.266164e-10, 
    1.263514e-10, 1.275318e-10, 1.278866e-10, 1.295523e-10, 1.288676e-10, 
    1.29958e-10, 1.289782e-10, 1.291516e-10, 1.299936e-10, 1.290311e-10, 
    1.311403e-10, 1.297087e-10, 1.323732e-10, 1.309379e-10, 1.324633e-10, 
    1.321858e-10, 1.326454e-10, 1.330576e-10, 1.33577e-10, 1.345375e-10, 
    1.343148e-10, 1.351197e-10, 1.269927e-10, 1.274741e-10, 1.274317e-10, 
    1.279363e-10, 1.2831e-10, 1.291216e-10, 1.304277e-10, 1.299359e-10, 
    1.308394e-10, 1.310211e-10, 1.296487e-10, 1.304906e-10, 1.277968e-10, 
    1.282304e-10, 1.279721e-10, 1.270306e-10, 1.300492e-10, 1.284963e-10, 
    1.313699e-10, 1.305241e-10, 1.329988e-10, 1.317657e-10, 1.341923e-10, 
    1.352352e-10, 1.362199e-10, 1.373743e-10, 1.277372e-10, 1.274097e-10, 
    1.279964e-10, 1.288099e-10, 1.295667e-10, 1.305756e-10, 1.306791e-10, 
    1.308685e-10, 1.313597e-10, 1.317734e-10, 1.309284e-10, 1.318771e-10, 
    1.28331e-10, 1.301843e-10, 1.27286e-10, 1.281558e-10, 1.287619e-10, 
    1.284959e-10, 1.298798e-10, 1.302068e-10, 1.315394e-10, 1.308499e-10, 
    1.349775e-10, 1.331448e-10, 1.382559e-10, 1.368196e-10, 1.272954e-10, 
    1.277361e-10, 1.292749e-10, 1.285418e-10, 1.306431e-10, 1.311625e-10, 
    1.315854e-10, 1.321268e-10, 1.321853e-10, 1.325066e-10, 1.319803e-10, 
    1.324858e-10, 1.305778e-10, 1.31429e-10, 1.290986e-10, 1.296642e-10, 
    1.294039e-10, 1.291186e-10, 1.3e-10, 1.309417e-10, 1.309619e-10, 
    1.312644e-10, 1.321186e-10, 1.306517e-10, 1.352148e-10, 1.323889e-10, 
    1.282174e-10, 1.290694e-10, 1.291913e-10, 1.288609e-10, 1.311104e-10, 
    1.302934e-10, 1.324988e-10, 1.319012e-10, 1.328809e-10, 1.323937e-10, 
    1.323221e-10, 1.316976e-10, 1.313094e-10, 1.303308e-10, 1.295369e-10, 
    1.289088e-10, 1.290547e-10, 1.297451e-10, 1.309994e-10, 1.321906e-10, 
    1.319293e-10, 1.328063e-10, 1.304903e-10, 1.314593e-10, 1.310844e-10, 
    1.320629e-10, 1.299229e-10, 1.317442e-10, 1.29459e-10, 1.296587e-10, 
    1.302772e-10, 1.315252e-10, 1.31802e-10, 1.320977e-10, 1.319152e-10, 
    1.310313e-10, 1.308867e-10, 1.302622e-10, 1.3009e-10, 1.296152e-10, 
    1.292227e-10, 1.295813e-10, 1.299583e-10, 1.310317e-10, 1.320021e-10, 
    1.330635e-10, 1.333238e-10, 1.345694e-10, 1.33555e-10, 1.352305e-10, 
    1.338054e-10, 1.362764e-10, 1.318502e-10, 1.337637e-10, 1.303054e-10, 
    1.306762e-10, 1.313478e-10, 1.328939e-10, 1.320583e-10, 1.330357e-10, 
    1.308811e-10, 1.297689e-10, 1.294819e-10, 1.289469e-10, 1.294941e-10, 
    1.294496e-10, 1.29974e-10, 1.298054e-10, 1.310674e-10, 1.303889e-10, 
    1.323203e-10, 1.33028e-10, 1.350353e-10, 1.362719e-10, 1.375355e-10, 
    1.380948e-10, 1.382653e-10, 1.383365e-10,
  1.281121e-10, 1.293278e-10, 1.29091e-10, 1.300747e-10, 1.295286e-10, 
    1.301733e-10, 1.283581e-10, 1.293762e-10, 1.287258e-10, 1.282213e-10, 
    1.319939e-10, 1.301187e-10, 1.339553e-10, 1.327494e-10, 1.357886e-10, 
    1.337673e-10, 1.361979e-10, 1.357301e-10, 1.371405e-10, 1.367357e-10, 
    1.385474e-10, 1.373275e-10, 1.394909e-10, 1.382556e-10, 1.384485e-10, 
    1.372874e-10, 1.30495e-10, 1.317598e-10, 1.304203e-10, 1.306002e-10, 
    1.305194e-10, 1.295399e-10, 1.290476e-10, 1.280194e-10, 1.282058e-10, 
    1.289611e-10, 1.306811e-10, 1.30096e-10, 1.315731e-10, 1.315396e-10, 
    1.331932e-10, 1.324464e-10, 1.352405e-10, 1.344435e-10, 1.367526e-10, 
    1.361701e-10, 1.367252e-10, 1.365568e-10, 1.367274e-10, 1.358736e-10, 
    1.362391e-10, 1.35489e-10, 1.325861e-10, 1.334361e-10, 1.309087e-10, 
    1.294001e-10, 1.284027e-10, 1.276972e-10, 1.277968e-10, 1.279868e-10, 
    1.289655e-10, 1.298889e-10, 1.305947e-10, 1.310678e-10, 1.315348e-10, 
    1.329533e-10, 1.337069e-10, 1.354019e-10, 1.350952e-10, 1.356149e-10, 
    1.361122e-10, 1.369492e-10, 1.368113e-10, 1.371806e-10, 1.356012e-10, 
    1.366499e-10, 1.349207e-10, 1.353926e-10, 1.31662e-10, 1.302538e-10, 
    1.296574e-10, 1.291365e-10, 1.278734e-10, 1.287451e-10, 1.284011e-10, 
    1.292201e-10, 1.297418e-10, 1.294836e-10, 1.310808e-10, 1.304587e-10, 
    1.337517e-10, 1.323285e-10, 1.360542e-10, 1.351581e-10, 1.362694e-10, 
    1.357018e-10, 1.36675e-10, 1.35799e-10, 1.373182e-10, 1.376501e-10, 
    1.374232e-10, 1.382956e-10, 1.357505e-10, 1.367252e-10, 1.294764e-10, 
    1.295185e-10, 1.297146e-10, 1.288535e-10, 1.288009e-10, 1.280143e-10, 
    1.287141e-10, 1.290127e-10, 1.29772e-10, 1.302222e-10, 1.306509e-10, 
    1.315957e-10, 1.326547e-10, 1.341425e-10, 1.352161e-10, 1.359382e-10, 
    1.354952e-10, 1.358862e-10, 1.354492e-10, 1.352445e-10, 1.375257e-10, 
    1.362425e-10, 1.381699e-10, 1.380629e-10, 1.371894e-10, 1.38075e-10, 
    1.29548e-10, 1.293059e-10, 1.28467e-10, 1.291233e-10, 1.279288e-10, 
    1.285968e-10, 1.289816e-10, 1.304717e-10, 1.308002e-10, 1.311052e-10, 
    1.317084e-10, 1.324846e-10, 1.338514e-10, 1.350462e-10, 1.361412e-10, 
    1.360608e-10, 1.360891e-10, 1.363343e-10, 1.357274e-10, 1.36434e-10, 
    1.365528e-10, 1.362424e-10, 1.380486e-10, 1.375314e-10, 1.380607e-10, 
    1.377238e-10, 1.293846e-10, 1.297922e-10, 1.295719e-10, 1.299864e-10, 
    1.296943e-10, 1.309955e-10, 1.313868e-10, 1.332253e-10, 1.324693e-10, 
    1.336735e-10, 1.325914e-10, 1.327828e-10, 1.337129e-10, 1.326497e-10, 
    1.349802e-10, 1.333981e-10, 1.363438e-10, 1.347564e-10, 1.364436e-10, 
    1.361365e-10, 1.366452e-10, 1.371015e-10, 1.376767e-10, 1.38741e-10, 
    1.384942e-10, 1.393864e-10, 1.304011e-10, 1.309319e-10, 1.308851e-10, 
    1.314416e-10, 1.318539e-10, 1.327497e-10, 1.341924e-10, 1.33649e-10, 
    1.346474e-10, 1.348483e-10, 1.333317e-10, 1.342619e-10, 1.312877e-10, 
    1.317661e-10, 1.314812e-10, 1.304429e-10, 1.337741e-10, 1.320595e-10, 
    1.352339e-10, 1.342989e-10, 1.370364e-10, 1.356717e-10, 1.383584e-10, 
    1.395146e-10, 1.406069e-10, 1.418887e-10, 1.31222e-10, 1.308608e-10, 
    1.315079e-10, 1.324056e-10, 1.332411e-10, 1.343559e-10, 1.344702e-10, 
    1.346796e-10, 1.352227e-10, 1.356802e-10, 1.347458e-10, 1.35795e-10, 
    1.318772e-10, 1.339235e-10, 1.307244e-10, 1.316839e-10, 1.323526e-10, 
    1.32059e-10, 1.33587e-10, 1.339483e-10, 1.354215e-10, 1.34659e-10, 
    1.392289e-10, 1.37198e-10, 1.428682e-10, 1.412727e-10, 1.307348e-10, 
    1.312208e-10, 1.32919e-10, 1.321097e-10, 1.344304e-10, 1.350046e-10, 
    1.354723e-10, 1.360712e-10, 1.36136e-10, 1.364915e-10, 1.359091e-10, 
    1.364685e-10, 1.343582e-10, 1.352993e-10, 1.327243e-10, 1.333489e-10, 
    1.330614e-10, 1.327464e-10, 1.337197e-10, 1.347605e-10, 1.347828e-10, 
    1.351173e-10, 1.360623e-10, 1.344399e-10, 1.39492e-10, 1.363615e-10, 
    1.317517e-10, 1.326921e-10, 1.328267e-10, 1.324618e-10, 1.34947e-10, 
    1.34044e-10, 1.364828e-10, 1.358216e-10, 1.369058e-10, 1.363665e-10, 
    1.362873e-10, 1.355964e-10, 1.351671e-10, 1.340853e-10, 1.332083e-10, 
    1.325147e-10, 1.326758e-10, 1.334382e-10, 1.348243e-10, 1.361418e-10, 
    1.358527e-10, 1.368233e-10, 1.342615e-10, 1.353329e-10, 1.349183e-10, 
    1.360006e-10, 1.336346e-10, 1.356482e-10, 1.331222e-10, 1.333428e-10, 
    1.340261e-10, 1.354057e-10, 1.357118e-10, 1.360391e-10, 1.358371e-10, 
    1.348596e-10, 1.346997e-10, 1.340095e-10, 1.338192e-10, 1.332947e-10, 
    1.328613e-10, 1.332573e-10, 1.336738e-10, 1.3486e-10, 1.359333e-10, 
    1.37108e-10, 1.373962e-10, 1.387764e-10, 1.376524e-10, 1.395096e-10, 
    1.3793e-10, 1.406698e-10, 1.357652e-10, 1.378836e-10, 1.340572e-10, 
    1.34467e-10, 1.352096e-10, 1.369203e-10, 1.359955e-10, 1.370773e-10, 
    1.346935e-10, 1.334646e-10, 1.331475e-10, 1.325568e-10, 1.33161e-10, 
    1.331118e-10, 1.33691e-10, 1.335047e-10, 1.348994e-10, 1.341494e-10, 
    1.362853e-10, 1.370688e-10, 1.392928e-10, 1.406647e-10, 1.420677e-10, 
    1.426892e-10, 1.428786e-10, 1.429578e-10,
  1.381727e-10, 1.394605e-10, 1.392096e-10, 1.402522e-10, 1.396732e-10, 
    1.403568e-10, 1.384332e-10, 1.395118e-10, 1.388226e-10, 1.382883e-10, 
    1.422883e-10, 1.402988e-10, 1.443716e-10, 1.430903e-10, 1.463214e-10, 
    1.441718e-10, 1.46757e-10, 1.46259e-10, 1.477606e-10, 1.473295e-10, 
    1.492601e-10, 1.479598e-10, 1.502664e-10, 1.489489e-10, 1.491546e-10, 
    1.479171e-10, 1.406978e-10, 1.420398e-10, 1.406185e-10, 1.408094e-10, 
    1.407237e-10, 1.396852e-10, 1.391636e-10, 1.380745e-10, 1.382718e-10, 
    1.390719e-10, 1.408953e-10, 1.402747e-10, 1.418414e-10, 1.418059e-10, 
    1.435617e-10, 1.427685e-10, 1.457381e-10, 1.448905e-10, 1.473475e-10, 
    1.467274e-10, 1.473184e-10, 1.47139e-10, 1.473207e-10, 1.464118e-10, 
    1.468008e-10, 1.460025e-10, 1.429169e-10, 1.438198e-10, 1.411366e-10, 
    1.395372e-10, 1.384804e-10, 1.377333e-10, 1.378388e-10, 1.3804e-10, 
    1.390766e-10, 1.400551e-10, 1.408035e-10, 1.413053e-10, 1.418008e-10, 
    1.43307e-10, 1.441076e-10, 1.459099e-10, 1.455836e-10, 1.461365e-10, 
    1.466657e-10, 1.475569e-10, 1.4741e-10, 1.478034e-10, 1.461219e-10, 
    1.472382e-10, 1.453979e-10, 1.459e-10, 1.41936e-10, 1.404419e-10, 
    1.398099e-10, 1.392578e-10, 1.3792e-10, 1.388431e-10, 1.384788e-10, 
    1.393463e-10, 1.398992e-10, 1.396256e-10, 1.413191e-10, 1.406593e-10, 
    1.441552e-10, 1.426434e-10, 1.46604e-10, 1.456505e-10, 1.46833e-10, 
    1.462289e-10, 1.472649e-10, 1.463323e-10, 1.479499e-10, 1.483036e-10, 
    1.480619e-10, 1.489915e-10, 1.462807e-10, 1.473184e-10, 1.396179e-10, 
    1.396625e-10, 1.398704e-10, 1.389579e-10, 1.389022e-10, 1.380691e-10, 
    1.388102e-10, 1.391265e-10, 1.399313e-10, 1.404085e-10, 1.408631e-10, 
    1.418655e-10, 1.429898e-10, 1.445705e-10, 1.457122e-10, 1.464805e-10, 
    1.460091e-10, 1.464252e-10, 1.459601e-10, 1.457424e-10, 1.48171e-10, 
    1.468045e-10, 1.488576e-10, 1.487435e-10, 1.478128e-10, 1.487564e-10, 
    1.396939e-10, 1.394372e-10, 1.385485e-10, 1.392438e-10, 1.379785e-10, 
    1.38686e-10, 1.390937e-10, 1.406732e-10, 1.410215e-10, 1.41345e-10, 
    1.419851e-10, 1.428091e-10, 1.442611e-10, 1.455314e-10, 1.466966e-10, 
    1.46611e-10, 1.466411e-10, 1.469021e-10, 1.462561e-10, 1.470083e-10, 
    1.471348e-10, 1.468043e-10, 1.487282e-10, 1.481771e-10, 1.487411e-10, 
    1.483821e-10, 1.395206e-10, 1.399527e-10, 1.397191e-10, 1.401585e-10, 
    1.398489e-10, 1.412287e-10, 1.416439e-10, 1.435959e-10, 1.427928e-10, 
    1.44072e-10, 1.429225e-10, 1.431258e-10, 1.44114e-10, 1.429844e-10, 
    1.454613e-10, 1.437795e-10, 1.469123e-10, 1.452233e-10, 1.470185e-10, 
    1.466915e-10, 1.472331e-10, 1.477191e-10, 1.483319e-10, 1.494664e-10, 
    1.492032e-10, 1.501549e-10, 1.405982e-10, 1.411612e-10, 1.411115e-10, 
    1.41702e-10, 1.421395e-10, 1.430906e-10, 1.446236e-10, 1.44046e-10, 
    1.451073e-10, 1.453209e-10, 1.437089e-10, 1.446975e-10, 1.415387e-10, 
    1.420464e-10, 1.417439e-10, 1.406426e-10, 1.44179e-10, 1.423579e-10, 
    1.457311e-10, 1.447368e-10, 1.476498e-10, 1.46197e-10, 1.490585e-10, 
    1.502918e-10, 1.514575e-10, 1.528269e-10, 1.41469e-10, 1.410858e-10, 
    1.417722e-10, 1.427253e-10, 1.436126e-10, 1.447973e-10, 1.449188e-10, 
    1.451415e-10, 1.457192e-10, 1.462059e-10, 1.45212e-10, 1.463281e-10, 
    1.421644e-10, 1.443377e-10, 1.409411e-10, 1.419591e-10, 1.42669e-10, 
    1.423573e-10, 1.4398e-10, 1.44364e-10, 1.459307e-10, 1.451196e-10, 
    1.499869e-10, 1.47822e-10, 1.538742e-10, 1.521687e-10, 1.409521e-10, 
    1.414676e-10, 1.432704e-10, 1.42411e-10, 1.448766e-10, 1.454872e-10, 
    1.459847e-10, 1.466221e-10, 1.46691e-10, 1.470695e-10, 1.464495e-10, 
    1.47045e-10, 1.447999e-10, 1.458007e-10, 1.430636e-10, 1.437271e-10, 
    1.434216e-10, 1.430871e-10, 1.441211e-10, 1.452276e-10, 1.452512e-10, 
    1.456071e-10, 1.466129e-10, 1.448866e-10, 1.502678e-10, 1.469313e-10, 
    1.42031e-10, 1.430295e-10, 1.431724e-10, 1.427849e-10, 1.454259e-10, 
    1.444658e-10, 1.470603e-10, 1.463564e-10, 1.475106e-10, 1.469364e-10, 
    1.468521e-10, 1.461167e-10, 1.4566e-10, 1.445098e-10, 1.435777e-10, 
    1.42841e-10, 1.430121e-10, 1.43822e-10, 1.452955e-10, 1.466973e-10, 
    1.463896e-10, 1.474227e-10, 1.44697e-10, 1.458364e-10, 1.453955e-10, 
    1.465469e-10, 1.440307e-10, 1.461721e-10, 1.434863e-10, 1.437206e-10, 
    1.444468e-10, 1.45914e-10, 1.462396e-10, 1.465879e-10, 1.463729e-10, 
    1.45333e-10, 1.45163e-10, 1.444291e-10, 1.442269e-10, 1.436695e-10, 
    1.432091e-10, 1.436298e-10, 1.440723e-10, 1.453334e-10, 1.464753e-10, 
    1.477261e-10, 1.480331e-10, 1.495044e-10, 1.483062e-10, 1.502866e-10, 
    1.486021e-10, 1.515248e-10, 1.462966e-10, 1.485525e-10, 1.444798e-10, 
    1.449154e-10, 1.457054e-10, 1.475262e-10, 1.465414e-10, 1.476934e-10, 
    1.451563e-10, 1.438501e-10, 1.435131e-10, 1.428858e-10, 1.435274e-10, 
    1.434752e-10, 1.440906e-10, 1.438927e-10, 1.453753e-10, 1.445778e-10, 
    1.4685e-10, 1.476843e-10, 1.50055e-10, 1.515193e-10, 1.530181e-10, 
    1.536826e-10, 1.538852e-10, 1.539699e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24532.39, 24552.28, 24548.38, 24564.66, 24555.6, 24566.3, 24536.39, 
    24553.08, 24542.39, 24534.16, 24596.99, 24565.39, 24630.84, 24609.91, 
    24662.94, 24627.55, 24670.21, 24661.91, 24687.12, 24679.83, 24712.87, 
    24690.51, 24730.47, 24707.48, 24711.04, 24689.79, 24571.68, 24593.01, 
    24570.43, 24573.45, 24572.09, 24555.78, 24547.67, 24530.89, 24533.91, 
    24546.25, 24574.81, 24565.02, 24589.85, 24589.28, 24617.57, 24604.71, 
    24653.28, 24639.37, 24680.13, 24669.71, 24679.64, 24676.62, 24679.68, 
    24664.45, 24670.94, 24657.65, 24607.1, 24621.78, 24578.63, 24553.47, 
    24537.12, 24525.67, 24527.28, 24530.36, 24546.32, 24561.57, 24573.35, 
    24581.32, 24589.2, 24613.42, 24626.5, 24656.12, 24650.73, 24659.87, 
    24668.68, 24683.67, 24681.19, 24687.85, 24659.63, 24678.29, 24647.67, 
    24655.95, 24591.36, 24567.65, 24557.73, 24549.13, 24528.52, 24542.71, 
    24537.09, 24550.5, 24559.12, 24554.85, 24581.54, 24571.07, 24627.28, 
    24602.69, 24667.65, 24651.83, 24671.48, 24661.41, 24678.74, 24663.12, 
    24690.34, 24696.38, 24692.25, 24708.22, 24662.27, 24679.64, 24554.73, 
    24555.43, 24558.68, 24544.48, 24543.62, 24530.8, 24542.2, 24547.09, 
    24559.63, 24567.12, 24574.3, 24590.23, 24608.28, 24634.12, 24652.85, 
    24665.59, 24657.76, 24664.67, 24656.95, 24653.35, 24694.12, 24671, 
    24705.91, 24703.94, 24688.01, 24704.16, 24555.92, 24551.92, 24538.16, 
    24548.91, 24529.42, 24540.28, 24546.58, 24571.29, 24576.81, 24581.95, 
    24592.14, 24605.36, 24629.02, 24649.87, 24669.2, 24667.77, 24668.27, 
    24672.64, 24661.86, 24674.42, 24676.55, 24671, 24703.68, 24694.22, 
    24703.9, 24697.73, 24553.21, 24559.96, 24556.31, 24563.19, 24558.34, 
    24580.1, 24586.7, 24618.12, 24605.1, 24625.92, 24607.19, 24610.48, 
    24626.61, 24608.2, 24648.71, 24621.12, 24672.81, 24644.81, 24674.59, 
    24669.11, 24678.2, 24686.42, 24696.87, 24716.46, 24711.89, 24728.51, 
    24570.11, 24579.03, 24578.24, 24587.62, 24594.61, 24609.91, 24635, 
    24625.49, 24642.91, 24646.41, 24619.97, 24636.22, 24585.03, 24593.12, 
    24588.29, 24570.81, 24627.67, 24598.1, 24653.16, 24636.86, 24685.24, 
    24660.88, 24709.38, 24730.92, 24751.62, 24776.28, 24583.92, 24577.83, 
    24588.74, 24604.01, 24618.4, 24637.85, 24639.83, 24643.47, 24652.96, 
    24661.02, 24644.62, 24663.05, 24595, 24630.29, 24575.53, 24591.72, 
    24603.1, 24598.09, 24624.41, 24630.72, 24656.46, 24643.11, 24725.55, 
    24688.17, 24795.25, 24764.45, 24575.71, 24583.9, 24612.83, 24598.96, 
    24639.14, 24649.14, 24657.35, 24667.95, 24669.1, 24675.45, 24665.07, 
    24675.04, 24637.89, 24654.31, 24609.48, 24620.27, 24615.29, 24609.86, 
    24626.72, 24644.88, 24645.27, 24651.12, 24667.8, 24639.3, 24730.5, 
    24673.13, 24592.87, 24608.92, 24611.24, 24604.97, 24648.13, 24632.4, 
    24675.29, 24663.53, 24682.89, 24673.21, 24671.8, 24659.54, 24651.99, 
    24633.12, 24617.83, 24605.88, 24608.64, 24621.82, 24645.99, 24669.21, 
    24664.08, 24681.4, 24636.21, 24654.9, 24647.63, 24666.7, 24625.24, 
    24660.46, 24616.34, 24620.16, 24632.08, 24656.18, 24661.58, 24667.38, 
    24663.8, 24646.61, 24643.82, 24631.79, 24628.46, 24619.33, 24611.83, 
    24618.68, 24625.92, 24646.61, 24665.5, 24686.54, 24691.76, 24717.12, 
    24696.43, 24730.83, 24701.51, 24752.83, 24662.53, 24700.65, 24632.63, 
    24639.77, 24652.74, 24683.15, 24666.61, 24685.98, 24643.71, 24622.28, 
    24616.78, 24606.6, 24617.01, 24616.16, 24626.22, 24622.97, 24647.3, 
    24634.25, 24671.77, 24685.83, 24726.75, 24752.73, 24779.72, 24791.76, 
    24795.46, 24797 ;

 GC_ICE1 =
  17606.64, 17638.41, 17632.18, 17658.19, 17643.71, 17660.81, 17613.03, 
    17639.69, 17622.62, 17609.47, 17709.79, 17659.36, 17763.81, 17730.41, 
    17814.93, 17758.57, 17826.49, 17813.28, 17853.4, 17841.79, 17894.37, 
    17858.79, 17922.36, 17885.8, 17891.46, 17857.64, 17669.4, 17703.45, 
    17667.4, 17672.22, 17670.05, 17644.01, 17631.04, 17604.24, 17609.07, 
    17628.78, 17674.39, 17658.75, 17698.4, 17697.5, 17742.63, 17722.11, 
    17799.54, 17777.4, 17842.28, 17825.7, 17841.49, 17836.69, 17841.56, 
    17817.32, 17827.65, 17806.5, 17725.94, 17749.36, 17680.5, 17640.32, 
    17614.19, 17595.91, 17598.49, 17603.4, 17628.89, 17653.25, 17672.07, 
    17684.79, 17697.37, 17736.02, 17756.88, 17804.06, 17795.48, 17810.04, 
    17824.06, 17847.91, 17843.96, 17854.56, 17809.65, 17839.34, 17790.62, 
    17803.8, 17700.81, 17662.95, 17647.12, 17633.38, 17600.46, 17623.12, 
    17614.15, 17635.57, 17649.35, 17642.52, 17685.14, 17668.43, 17758.13, 
    17718.89, 17822.42, 17797.24, 17828.51, 17812.48, 17840.06, 17815.21, 
    17858.53, 17868.13, 17861.56, 17886.97, 17813.85, 17841.49, 17642.33, 
    17643.44, 17648.63, 17625.96, 17624.58, 17604.11, 17622.31, 17630.13, 
    17650.15, 17662.11, 17673.57, 17699.01, 17727.82, 17769.05, 17798.86, 
    17819.14, 17806.67, 17817.67, 17805.38, 17799.65, 17864.53, 17827.75, 
    17883.29, 17880.16, 17854.81, 17880.51, 17644.22, 17637.83, 17615.87, 
    17633.03, 17601.9, 17619.25, 17629.31, 17668.78, 17677.58, 17685.8, 
    17702.05, 17723.16, 17760.91, 17794.12, 17824.88, 17822.6, 17823.4, 
    17830.35, 17813.2, 17833.19, 17836.57, 17827.75, 17879.74, 17864.69, 
    17880.09, 17870.27, 17639.91, 17650.68, 17644.85, 17655.84, 17648.09, 
    17682.84, 17693.38, 17743.52, 17722.74, 17755.95, 17726.08, 17731.33, 
    17757.05, 17727.68, 17792.28, 17748.31, 17830.62, 17786.06, 17833.46, 
    17824.74, 17839.21, 17852.28, 17868.9, 17900.07, 17892.8, 17919.24, 
    17666.89, 17681.13, 17679.87, 17694.86, 17705.99, 17730.42, 17770.45, 
    17755.27, 17783.04, 17788.61, 17746.46, 17772.39, 17690.72, 17703.62, 
    17695.92, 17668.01, 17758.76, 17711.57, 17799.36, 17773.41, 17850.41, 
    17811.63, 17888.81, 17923.07, 17955.99, 17995.14, 17688.95, 17679.21, 
    17696.64, 17721, 17743.96, 17774.98, 17778.13, 17783.93, 17799.04, 
    17811.87, 17785.77, 17815.1, 17706.63, 17762.92, 17675.55, 17701.39, 
    17719.55, 17711.56, 17753.54, 17763.61, 17804.61, 17783.36, 17914.54, 
    17855.06, 18025.23, 17976.38, 17675.82, 17688.92, 17735.07, 17712.93, 
    17777.04, 17792.96, 17806.03, 17822.9, 17824.73, 17834.83, 17818.32, 
    17834.17, 17775.04, 17801.19, 17729.72, 17746.94, 17738.99, 17730.33, 
    17757.24, 17786.17, 17786.79, 17796.1, 17822.66, 17777.3, 17922.4, 
    17831.13, 17703.22, 17728.84, 17732.53, 17722.53, 17791.36, 17766.29, 
    17834.58, 17815.85, 17846.66, 17831.27, 17829.02, 17809.51, 17797.49, 
    17767.45, 17743.05, 17723.98, 17728.39, 17749.41, 17787.94, 17824.9, 
    17816.73, 17844.3, 17772.38, 17802.12, 17790.56, 17820.9, 17754.87, 
    17810.98, 17740.67, 17746.77, 17765.79, 17804.17, 17812.76, 17821.99, 
    17816.29, 17788.92, 17784.49, 17765.32, 17760.01, 17745.44, 17733.48, 
    17744.4, 17755.96, 17788.93, 17819, 17852.47, 17860.78, 17901.12, 
    17868.21, 17922.93, 17876.29, 17957.91, 17814.27, 17874.93, 17766.66, 
    17778.04, 17798.68, 17847.08, 17820.76, 17851.59, 17784.31, 17750.15, 
    17741.37, 17725.13, 17741.74, 17740.38, 17756.44, 17751.26, 17790.03, 
    17769.24, 17828.96, 17851.34, 17916.44, 17957.75, 18000.62, 18019.7, 
    18025.55, 18028 ;

 GC_LIQ1 =
  5232.799, 5234.828, 5234.43, 5236.092, 5235.167, 5236.259, 5233.207, 
    5234.91, 5233.819, 5232.98, 5239.4, 5236.167, 5242.88, 5240.728, 5246.23, 
    5242.542, 5246.992, 5246.121, 5248.765, 5248, 5251.466, 5249.12, 
    5253.315, 5250.9, 5251.274, 5249.044, 5236.808, 5238.992, 5236.681, 
    5236.988, 5236.85, 5235.186, 5234.357, 5232.646, 5232.954, 5234.212, 
    5237.127, 5236.128, 5238.667, 5238.608, 5241.515, 5240.194, 5245.218, 
    5243.762, 5248.032, 5246.939, 5247.98, 5247.663, 5247.984, 5246.388, 
    5247.068, 5245.675, 5240.44, 5241.949, 5237.518, 5234.95, 5233.281, 
    5232.114, 5232.278, 5232.592, 5234.22, 5235.776, 5236.979, 5237.792, 
    5238.6, 5241.089, 5242.434, 5245.515, 5244.951, 5245.908, 5246.832, 
    5248.403, 5248.142, 5248.841, 5245.883, 5247.838, 5244.631, 5245.498, 
    5238.822, 5236.396, 5235.384, 5234.507, 5232.405, 5233.852, 5233.278, 
    5234.647, 5235.527, 5235.09, 5237.814, 5236.746, 5242.514, 5239.986, 
    5246.723, 5245.066, 5247.125, 5246.069, 5247.886, 5246.249, 5249.103, 
    5249.736, 5249.303, 5250.978, 5246.159, 5247.98, 5235.078, 5235.149, 
    5235.481, 5234.033, 5233.945, 5232.637, 5233.8, 5234.299, 5235.578, 
    5236.343, 5237.075, 5238.706, 5240.561, 5243.217, 5245.173, 5246.507, 
    5245.687, 5246.411, 5245.602, 5245.225, 5249.498, 5247.075, 5250.735, 
    5250.528, 5248.858, 5250.552, 5235.199, 5234.791, 5233.388, 5234.484, 
    5232.496, 5233.604, 5234.247, 5236.769, 5237.332, 5237.856, 5238.902, 
    5240.261, 5242.693, 5244.861, 5246.885, 5246.735, 5246.788, 5247.246, 
    5246.116, 5247.433, 5247.656, 5247.074, 5250.501, 5249.509, 5250.524, 
    5249.877, 5234.924, 5235.612, 5235.239, 5235.941, 5235.446, 5237.667, 
    5238.344, 5241.573, 5240.234, 5242.374, 5240.449, 5240.787, 5242.444, 
    5240.552, 5244.741, 5241.881, 5247.264, 5244.332, 5247.451, 5246.876, 
    5247.829, 5248.691, 5249.787, 5251.843, 5251.363, 5253.109, 5236.647, 
    5237.558, 5237.478, 5238.438, 5239.156, 5240.729, 5243.308, 5242.33, 
    5244.133, 5244.499, 5241.762, 5243.433, 5238.172, 5239.002, 5238.507, 
    5236.719, 5242.554, 5239.515, 5245.206, 5243.5, 5248.568, 5246.013, 
    5251.099, 5253.363, 5255.544, 5258.163, 5238.058, 5237.436, 5238.553, 
    5240.122, 5241.601, 5243.604, 5243.811, 5244.191, 5245.185, 5246.029, 
    5244.312, 5246.242, 5239.197, 5242.823, 5237.201, 5238.859, 5240.029, 
    5239.514, 5242.218, 5242.867, 5245.551, 5244.154, 5252.799, 5248.875, 
    5260.208, 5256.896, 5237.219, 5238.056, 5241.028, 5239.603, 5243.738, 
    5244.785, 5245.645, 5246.755, 5246.875, 5247.541, 5246.453, 5247.498, 
    5243.608, 5245.326, 5240.684, 5241.793, 5241.281, 5240.723, 5242.456, 
    5244.339, 5244.379, 5244.992, 5246.739, 5243.756, 5253.318, 5247.298, 
    5238.978, 5240.627, 5240.865, 5240.221, 5244.68, 5243.04, 5247.524, 
    5246.291, 5248.321, 5247.307, 5247.158, 5245.874, 5245.083, 5243.114, 
    5241.542, 5240.314, 5240.598, 5241.952, 5244.456, 5246.887, 5246.349, 
    5248.165, 5243.433, 5245.388, 5244.627, 5246.624, 5242.304, 5245.97, 
    5241.389, 5241.782, 5243.007, 5245.522, 5246.087, 5246.695, 5246.32, 
    5244.52, 5244.228, 5242.977, 5242.635, 5241.696, 5240.926, 5241.629, 
    5242.374, 5244.521, 5246.499, 5248.704, 5249.251, 5251.913, 5249.741, 
    5253.353, 5250.273, 5255.672, 5246.187, 5250.184, 5243.063, 5243.805, 
    5245.161, 5248.348, 5246.614, 5248.646, 5244.217, 5242, 5241.434, 
    5240.388, 5241.458, 5241.371, 5242.405, 5242.071, 5244.593, 5243.23, 
    5247.155, 5248.629, 5252.925, 5255.661, 5258.533, 5259.831, 5260.229, 
    5260.396 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.958688e-09, 8.998072e-09, 8.990416e-09, 9.022181e-09, 9.004559e-09, 
    9.02536e-09, 8.966672e-09, 8.999636e-09, 8.978592e-09, 8.962233e-09, 
    9.083827e-09, 9.023598e-09, 9.146384e-09, 9.107973e-09, 9.20446e-09, 
    9.140408e-09, 9.217374e-09, 9.202611e-09, 9.247044e-09, 9.234315e-09, 
    9.29115e-09, 9.252919e-09, 9.32061e-09, 9.28202e-09, 9.288057e-09, 
    9.251658e-09, 9.035718e-09, 9.076329e-09, 9.033312e-09, 9.039103e-09, 
    9.036504e-09, 9.004924e-09, 8.98901e-09, 8.955677e-09, 8.961728e-09, 
    8.98621e-09, 9.041707e-09, 9.022868e-09, 9.070344e-09, 9.069272e-09, 
    9.122129e-09, 9.098297e-09, 9.187134e-09, 9.161885e-09, 9.234846e-09, 
    9.216497e-09, 9.233984e-09, 9.228682e-09, 9.234054e-09, 9.207143e-09, 
    9.218673e-09, 9.194992e-09, 9.10276e-09, 9.129868e-09, 9.049021e-09, 
    9.000409e-09, 8.968118e-09, 8.945205e-09, 8.948444e-09, 8.954619e-09, 
    8.986353e-09, 9.016188e-09, 9.038924e-09, 9.054133e-09, 9.069119e-09, 
    9.114481e-09, 9.138486e-09, 9.19224e-09, 9.182538e-09, 9.198973e-09, 
    9.214672e-09, 9.24103e-09, 9.236692e-09, 9.248305e-09, 9.198538e-09, 
    9.231614e-09, 9.177012e-09, 9.191947e-09, 9.073196e-09, 9.02795e-09, 
    9.008721e-09, 8.991887e-09, 8.950934e-09, 8.979216e-09, 8.968067e-09, 
    8.994589e-09, 9.011442e-09, 9.003107e-09, 9.054549e-09, 9.03455e-09, 
    9.139909e-09, 9.094528e-09, 9.212841e-09, 9.18453e-09, 9.219627e-09, 
    9.201717e-09, 9.232404e-09, 9.204786e-09, 9.252627e-09, 9.263045e-09, 
    9.255926e-09, 9.283271e-09, 9.203255e-09, 9.233984e-09, 9.002874e-09, 
    9.004233e-09, 9.010567e-09, 8.982727e-09, 8.981025e-09, 8.955512e-09, 
    8.978213e-09, 8.98788e-09, 9.012419e-09, 9.026935e-09, 9.040733e-09, 
    9.071071e-09, 9.104952e-09, 9.15233e-09, 9.186365e-09, 9.209179e-09, 
    9.195189e-09, 9.207541e-09, 9.193734e-09, 9.187262e-09, 9.259141e-09, 
    9.21878e-09, 9.279337e-09, 9.275986e-09, 9.248581e-09, 9.276365e-09, 
    9.005188e-09, 8.997365e-09, 8.970204e-09, 8.99146e-09, 8.952733e-09, 
    8.974411e-09, 8.986876e-09, 9.034969e-09, 9.045534e-09, 9.055332e-09, 
    9.074683e-09, 9.099517e-09, 9.143081e-09, 9.180985e-09, 9.215585e-09, 
    9.21305e-09, 9.213942e-09, 9.221672e-09, 9.202525e-09, 9.224816e-09, 
    9.228557e-09, 9.218775e-09, 9.275538e-09, 9.259321e-09, 9.275915e-09, 
    9.265356e-09, 8.999907e-09, 9.01307e-09, 9.005958e-09, 9.019333e-09, 
    9.00991e-09, 9.051811e-09, 9.064373e-09, 9.123153e-09, 9.099028e-09, 
    9.137421e-09, 9.102928e-09, 9.10904e-09, 9.138676e-09, 9.104792e-09, 
    9.178896e-09, 9.128657e-09, 9.221973e-09, 9.171807e-09, 9.225117e-09, 
    9.215436e-09, 9.231464e-09, 9.245819e-09, 9.263879e-09, 9.297202e-09, 
    9.289486e-09, 9.317352e-09, 9.032694e-09, 9.049767e-09, 9.048263e-09, 
    9.06613e-09, 9.079343e-09, 9.107982e-09, 9.153915e-09, 9.136643e-09, 
    9.168352e-09, 9.174718e-09, 9.126543e-09, 9.156122e-09, 9.061193e-09, 
    9.076532e-09, 9.067398e-09, 9.034041e-09, 9.140624e-09, 9.085927e-09, 
    9.186928e-09, 9.157296e-09, 9.243773e-09, 9.200767e-09, 9.285237e-09, 
    9.32135e-09, 9.355333e-09, 9.39505e-09, 9.059084e-09, 9.047484e-09, 
    9.068255e-09, 9.096993e-09, 9.123656e-09, 9.159104e-09, 9.16273e-09, 
    9.169371e-09, 9.186572e-09, 9.201035e-09, 9.171472e-09, 9.20466e-09, 
    9.08009e-09, 9.145372e-09, 9.043098e-09, 9.073896e-09, 9.0953e-09, 
    9.08591e-09, 9.134668e-09, 9.14616e-09, 9.192859e-09, 9.168718e-09, 
    9.312438e-09, 9.248852e-09, 9.425289e-09, 9.375984e-09, 9.04343e-09, 
    9.059044e-09, 9.113386e-09, 9.08753e-09, 9.16147e-09, 9.17967e-09, 
    9.194465e-09, 9.213379e-09, 9.21542e-09, 9.226626e-09, 9.208263e-09, 
    9.2259e-09, 9.159179e-09, 9.188995e-09, 9.107173e-09, 9.127089e-09, 
    9.117927e-09, 9.107877e-09, 9.138893e-09, 9.171937e-09, 9.172642e-09, 
    9.183238e-09, 9.213099e-09, 9.161769e-09, 9.320647e-09, 9.222531e-09, 
    9.07607e-09, 9.106146e-09, 9.11044e-09, 9.09879e-09, 9.177845e-09, 
    9.149201e-09, 9.226352e-09, 9.205501e-09, 9.239665e-09, 9.222688e-09, 
    9.220191e-09, 9.198386e-09, 9.184811e-09, 9.150515e-09, 9.122608e-09, 
    9.100479e-09, 9.105625e-09, 9.129934e-09, 9.173958e-09, 9.215605e-09, 
    9.206483e-09, 9.237069e-09, 9.156109e-09, 9.190058e-09, 9.176937e-09, 
    9.211148e-09, 9.136183e-09, 9.200025e-09, 9.119866e-09, 9.126894e-09, 
    9.148633e-09, 9.192362e-09, 9.202034e-09, 9.212364e-09, 9.205989e-09, 
    9.175076e-09, 9.170011e-09, 9.148104e-09, 9.142056e-09, 9.125364e-09, 
    9.111544e-09, 9.124171e-09, 9.137431e-09, 9.175088e-09, 9.209025e-09, 
    9.246024e-09, 9.255078e-09, 9.298311e-09, 9.263119e-09, 9.321194e-09, 
    9.271822e-09, 9.357285e-09, 9.203722e-09, 9.270368e-09, 9.149622e-09, 
    9.16263e-09, 9.186159e-09, 9.240122e-09, 9.210988e-09, 9.245059e-09, 
    9.169812e-09, 9.130773e-09, 9.12067e-09, 9.101825e-09, 9.121101e-09, 
    9.119534e-09, 9.137979e-09, 9.132052e-09, 9.176339e-09, 9.15255e-09, 
    9.220129e-09, 9.24479e-09, 9.314432e-09, 9.357126e-09, 9.400582e-09, 
    9.419768e-09, 9.425607e-09, 9.428049e-09 ;

 H2OCAN =
  0.07672506, 0.07670978, 0.07671268, 0.07670048, 0.07670714, 0.07669923, 
    0.07672183, 0.07670929, 0.07671722, 0.07672349, 0.07667709, 0.0766999, 
    0.07665224, 0.07666693, 0.0766295, 0.07665472, 0.07662432, 0.07662991, 
    0.07661226, 0.07661731, 0.07659526, 0.07660992, 0.07658322, 0.0765986, 
    0.07659632, 0.07661045, 0.07669501, 0.07668001, 0.07669597, 0.07669382, 
    0.07669471, 0.07670711, 0.07671354, 0.076726, 0.07672369, 0.07671441, 
    0.07669284, 0.07669998, 0.07668134, 0.07668176, 0.0766614, 0.07667059, 
    0.076636, 0.0766458, 0.07661709, 0.07662439, 0.07661749, 0.07661954, 
    0.07661746, 0.07662815, 0.0766236, 0.07663287, 0.07666893, 0.07665846, 
    0.07668988, 0.0767093, 0.07672133, 0.07673008, 0.07672884, 0.07672656, 
    0.07671437, 0.07670258, 0.07669366, 0.07668773, 0.07668182, 0.07666495, 
    0.07665532, 0.07663417, 0.07663774, 0.07663148, 0.07662511, 0.07661473, 
    0.07661641, 0.07661188, 0.07663145, 0.07661857, 0.07663982, 0.07663406, 
    0.07668129, 0.07669801, 0.07670599, 0.07671216, 0.07672792, 0.07671711, 
    0.0767214, 0.07671095, 0.07670444, 0.07670762, 0.07668757, 0.07669542, 
    0.07665475, 0.07667221, 0.07662585, 0.07663698, 0.07662313, 0.07663016, 
    0.0766182, 0.07662896, 0.07661012, 0.07660612, 0.07660887, 0.07659789, 
    0.07662959, 0.07661759, 0.07670776, 0.07670725, 0.07670474, 0.07671577, 
    0.07671638, 0.07672612, 0.07671736, 0.0767137, 0.07670398, 0.07669841, 
    0.07669304, 0.07668116, 0.07666823, 0.07664977, 0.07663627, 0.07662722, 
    0.07663271, 0.07662787, 0.07663332, 0.07663582, 0.07660768, 0.07662362, 
    0.07659948, 0.07660078, 0.07661182, 0.07660063, 0.07670687, 0.07670984, 
    0.07672049, 0.07671216, 0.07672717, 0.07671891, 0.07671423, 0.07669549, 
    0.0766911, 0.07668735, 0.07667971, 0.07667013, 0.07665333, 0.07663849, 
    0.07662469, 0.07662568, 0.07662535, 0.07662236, 0.07662989, 0.07662112, 
    0.07661974, 0.07662349, 0.07660096, 0.07660741, 0.07660081, 0.07660498, 
    0.07670885, 0.07670379, 0.07670654, 0.07670143, 0.07670512, 0.07668897, 
    0.07668411, 0.07666127, 0.07667037, 0.07665558, 0.07666879, 0.07666651, 
    0.07665554, 0.07666801, 0.07663952, 0.07665925, 0.07662224, 0.07664254, 
    0.076621, 0.07662475, 0.07661842, 0.07661285, 0.07660562, 0.07659253, 
    0.07659552, 0.07658436, 0.07669614, 0.07668963, 0.07669001, 0.07668304, 
    0.07667797, 0.07666679, 0.07664902, 0.07665564, 0.07664325, 0.07664083, 
    0.07665954, 0.07664825, 0.07668512, 0.07667934, 0.07668263, 0.07669574, 
    0.0766544, 0.07667567, 0.07663608, 0.07664765, 0.07661366, 0.07663085, 
    0.07659722, 0.07658322, 0.07656902, 0.07655343, 0.07668586, 0.07669031, 
    0.07668216, 0.07667136, 0.07666078, 0.07664698, 0.07664546, 0.07664293, 
    0.0766361, 0.07663044, 0.07664232, 0.076629, 0.07667841, 0.07665245, 
    0.07669217, 0.07668041, 0.07667191, 0.07667543, 0.07665635, 0.07665192, 
    0.07663387, 0.0766431, 0.07658686, 0.07661195, 0.0765408, 0.07656103, 
    0.07669191, 0.07668578, 0.0766649, 0.07667477, 0.07664596, 0.07663891, 
    0.07663299, 0.07662573, 0.0766248, 0.07662045, 0.07662758, 0.07662065, 
    0.07664696, 0.07663521, 0.07666705, 0.07665944, 0.07666288, 0.07666678, 
    0.07665473, 0.07664219, 0.0766416, 0.07663761, 0.07662692, 0.07664584, 
    0.07658421, 0.07662304, 0.07667913, 0.07666789, 0.07666589, 0.07667032, 
    0.07663963, 0.07665082, 0.07662051, 0.07662868, 0.07661519, 0.07662193, 
    0.07662294, 0.07663148, 0.07663687, 0.07665037, 0.07666122, 0.07666963, 
    0.07666766, 0.07665839, 0.07664134, 0.07662486, 0.07662852, 0.07661622, 
    0.07664807, 0.07663494, 0.07664013, 0.07662651, 0.07665589, 0.07663187, 
    0.07666212, 0.07665941, 0.07665104, 0.07663427, 0.07663005, 0.07662613, 
    0.07662848, 0.07664084, 0.07664271, 0.07665116, 0.07665365, 0.07665998, 
    0.07666535, 0.07666052, 0.0766555, 0.0766407, 0.07662746, 0.07661282, 
    0.07660909, 0.07659265, 0.07660649, 0.07658406, 0.07660383, 0.07656916, 
    0.07663, 0.07660374, 0.07665055, 0.07664548, 0.07663663, 0.07661546, 
    0.07662657, 0.07661341, 0.07664277, 0.07665823, 0.07666183, 0.07666919, 
    0.07666166, 0.07666226, 0.07665507, 0.07665736, 0.07664021, 0.07664942, 
    0.07662305, 0.07661343, 0.07658566, 0.07656866, 0.07655071, 0.07654291, 
    0.07654051, 0.07653952 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  3.864273, 3.877373, 3.874824, 3.885409, 3.879536, 3.88647, 3.866928, 
    3.877892, 3.870891, 3.865453, 3.906011, 3.885882, 3.927028, 3.914122, 
    3.946614, 3.925015, 3.950981, 3.945994, 3.96103, 3.956718, 3.975991, 
    3.963022, 3.986018, 3.972893, 3.974942, 3.962594, 3.88993, 3.903499, 
    3.889126, 3.891059, 3.890193, 3.879656, 3.874352, 3.863276, 3.865286, 
    3.873423, 3.891928, 3.885641, 3.90151, 3.901151, 3.918876, 3.910876, 
    3.940767, 3.932254, 3.956898, 3.950689, 3.956606, 3.954811, 3.956629, 
    3.947525, 3.951423, 3.943421, 3.912373, 3.921476, 3.894374, 3.878145, 
    3.867407, 3.859799, 3.860874, 3.862923, 3.873471, 3.883413, 3.891003, 
    3.896086, 3.9011, 3.916298, 3.924371, 3.942488, 3.939218, 3.944763, 
    3.950071, 3.958992, 3.957523, 3.961456, 3.944619, 3.955801, 3.937355, 
    3.942393, 3.902449, 3.887337, 3.880916, 3.875313, 3.8617, 3.871096, 
    3.86739, 3.876216, 3.88183, 3.879053, 3.896224, 3.889541, 3.92485, 
    3.90961, 3.949452, 3.939889, 3.951747, 3.945693, 3.956069, 3.94673, 
    3.962922, 3.966453, 3.964039, 3.973321, 3.946213, 3.956604, 3.878975, 
    3.879427, 3.881539, 3.872264, 3.871698, 3.86322, 3.870764, 3.87398, 
    3.882157, 3.886998, 3.891606, 3.901752, 3.913106, 3.929032, 3.940508, 
    3.948215, 3.943489, 3.947661, 3.942997, 3.940813, 3.965128, 3.951459, 
    3.971985, 3.970848, 3.961549, 3.970976, 3.879745, 3.87714, 3.868101, 
    3.875174, 3.862298, 3.869499, 3.873643, 3.889677, 3.893211, 3.896485, 
    3.902962, 3.911285, 3.92592, 3.938691, 3.950381, 3.949524, 3.949826, 
    3.952439, 3.945966, 3.953502, 3.954767, 3.951459, 3.970695, 3.965192, 
    3.970824, 3.96724, 3.877987, 3.882374, 3.880003, 3.884461, 3.881319, 
    3.895304, 3.899505, 3.919216, 3.91112, 3.924015, 3.91243, 3.91448, 
    3.92443, 3.913056, 3.937983, 3.921064, 3.95254, 3.935589, 3.953604, 
    3.95033, 3.955754, 3.960614, 3.966738, 3.978053, 3.975431, 3.984911, 
    3.888921, 3.894623, 3.894123, 3.900099, 3.904522, 3.914127, 3.929568, 
    3.923757, 3.934434, 3.936579, 3.920362, 3.93031, 3.898444, 3.903576, 
    3.900522, 3.889369, 3.925091, 3.906724, 3.940698, 3.930708, 3.95992, 
    3.945368, 3.973988, 3.986265, 3.997859, 4.011427, 3.89774, 3.893863, 
    3.90081, 3.910435, 3.91939, 3.931316, 3.932539, 3.934776, 3.94058, 
    3.945463, 3.935481, 3.946688, 3.904761, 3.92669, 3.892395, 3.902693, 
    3.909868, 3.906722, 3.923094, 3.926959, 3.942698, 3.934557, 3.98323, 
    3.961637, 4.02179, 4.004908, 3.892508, 3.897728, 3.915938, 3.907265, 
    3.932114, 3.938249, 3.943244, 3.949632, 3.950325, 3.954114, 3.947905, 
    3.95387, 3.931341, 3.941396, 3.913856, 3.920543, 3.917467, 3.914092, 
    3.924514, 3.935638, 3.93588, 3.939451, 3.949522, 3.932215, 3.986016, 
    3.952714, 3.903427, 3.913504, 3.914951, 3.911043, 3.937634, 3.927981, 
    3.954022, 3.946972, 3.95853, 3.952783, 3.951938, 3.944568, 3.939984, 
    3.928423, 3.919037, 3.91161, 3.913336, 3.921499, 3.93632, 3.950385, 
    3.9473, 3.957651, 3.930308, 3.941753, 3.937325, 3.94888, 3.923601, 
    3.945106, 3.918118, 3.920479, 3.92779, 3.942527, 3.9458, 3.949289, 
    3.947137, 3.936698, 3.934991, 3.927613, 3.925576, 3.919966, 3.915323, 
    3.919563, 3.924019, 3.936704, 3.94816, 3.960682, 3.963753, 3.978422, 
    3.966472, 3.986201, 3.969414, 3.998513, 3.946362, 3.96893, 3.928125, 
    3.932506, 3.940435, 3.958678, 3.948826, 3.960352, 3.934925, 3.921778, 
    3.918388, 3.91206, 3.918533, 3.918006, 3.924207, 3.922214, 3.937125, 
    3.92911, 3.951916, 3.960262, 3.983915, 3.998466, 4.013327, 4.019899, 
    4.021902, 4.022739,
  3.292639, 3.30539, 3.30291, 3.313153, 3.307498, 3.314159, 3.295225, 
    3.305894, 3.299082, 3.29379, 3.332687, 3.313602, 3.352645, 3.340398, 
    3.371245, 3.350732, 3.375395, 3.370661, 3.384948, 3.380851, 3.399157, 
    3.386841, 3.408693, 3.396218, 3.398163, 3.386433, 3.317445, 3.330303, 
    3.316682, 3.318513, 3.317693, 3.307613, 3.302446, 3.291672, 3.293627, 
    3.301545, 3.319337, 3.313377, 3.328433, 3.328092, 3.344911, 3.337319, 
    3.365697, 3.357614, 3.381022, 3.375121, 3.380743, 3.379039, 3.380765, 
    3.372115, 3.375819, 3.368218, 3.338738, 3.347377, 3.321659, 3.306137, 
    3.295691, 3.288288, 3.289333, 3.291326, 3.301591, 3.311264, 3.318463, 
    3.323285, 3.328043, 3.342454, 3.350123, 3.367329, 3.364226, 3.36949, 
    3.374535, 3.383009, 3.381614, 3.38535, 3.369356, 3.379976, 3.362458, 
    3.367241, 3.329306, 3.314986, 3.308835, 3.303386, 3.290137, 3.29928, 
    3.295673, 3.304266, 3.309732, 3.307029, 3.323417, 3.317076, 3.350578, 
    3.336114, 3.373946, 3.364864, 3.376127, 3.370378, 3.380232, 3.371362, 
    3.386744, 3.390097, 3.387805, 3.396628, 3.37087, 3.38074, 3.306952, 
    3.307392, 3.309448, 3.300417, 3.299866, 3.291617, 3.298959, 3.302088, 
    3.310051, 3.314664, 3.319034, 3.32866, 3.339432, 3.35455, 3.365451, 
    3.372773, 3.368284, 3.372247, 3.367816, 3.365742, 3.388838, 3.375851, 
    3.395358, 3.394277, 3.385438, 3.394399, 3.307702, 3.305166, 3.296366, 
    3.303252, 3.29072, 3.297726, 3.301759, 3.317202, 3.320558, 3.323663, 
    3.329809, 3.337707, 3.351596, 3.363724, 3.37483, 3.374016, 3.374302, 
    3.376784, 3.370636, 3.377795, 3.378994, 3.375854, 3.394132, 3.388902, 
    3.394254, 3.390849, 3.305991, 3.310261, 3.307953, 3.312257, 3.309232, 
    3.322538, 3.326523, 3.345229, 3.33755, 3.349787, 3.338794, 3.340738, 
    3.350174, 3.339389, 3.363048, 3.346982, 3.37688, 3.360771, 3.377891, 
    3.374782, 3.379934, 3.384551, 3.390371, 3.401122, 3.398632, 3.407643, 
    3.316489, 3.321894, 3.321424, 3.327092, 3.331288, 3.340405, 3.355062, 
    3.349546, 3.359684, 3.36172, 3.346323, 3.355764, 3.325521, 3.330386, 
    3.327493, 3.316911, 3.350808, 3.333374, 3.365631, 3.356144, 3.383891, 
    3.370064, 3.39726, 3.408924, 3.419957, 3.432855, 3.324854, 3.321177, 
    3.327769, 3.336895, 3.345399, 3.356721, 3.357885, 3.360008, 3.36552, 
    3.370158, 3.360674, 3.371322, 3.331503, 3.352327, 3.319782, 3.329547, 
    3.33636, 3.333376, 3.348917, 3.352587, 3.367529, 3.359802, 3.406037, 
    3.385518, 3.44272, 3.426655, 3.319891, 3.324844, 3.34212, 3.333892, 
    3.357481, 3.363306, 3.368052, 3.374116, 3.374776, 3.378375, 3.372478, 
    3.378144, 3.356745, 3.366295, 3.340149, 3.346494, 3.343576, 3.340373, 
    3.350266, 3.360821, 3.361057, 3.364446, 3.373994, 3.357578, 3.408675, 
    3.377029, 3.330251, 3.339808, 3.341186, 3.337478, 3.362721, 3.353556, 
    3.378289, 3.371592, 3.382572, 3.377111, 3.376308, 3.369308, 3.364954, 
    3.353974, 3.345064, 3.338017, 3.339655, 3.3474, 3.36147, 3.374831, 
    3.3719, 3.381737, 3.355766, 3.366632, 3.362426, 3.373403, 3.349397, 
    3.369802, 3.344194, 3.346435, 3.353374, 3.367363, 3.370479, 3.373791, 
    3.371748, 3.36183, 3.360211, 3.353208, 3.351271, 3.345948, 3.341541, 
    3.345565, 3.349793, 3.361838, 3.372718, 3.384615, 3.387535, 3.401464, 
    3.390109, 3.40885, 3.392892, 3.420563, 3.371002, 3.392442, 3.353693, 
    3.357853, 3.365377, 3.382705, 3.373352, 3.384298, 3.360149, 3.347663, 
    3.34445, 3.338444, 3.344588, 3.344088, 3.349974, 3.348083, 3.362239, 
    3.354629, 3.376286, 3.384214, 3.406695, 3.420528, 3.43467, 3.440923, 
    3.442829, 3.443625,
  3.019191, 3.033293, 3.030548, 3.04195, 3.035621, 3.043092, 3.022047, 
    3.033854, 3.026313, 3.020459, 3.064165, 3.042459, 3.086834, 3.072903, 
    3.107873, 3.084663, 3.112446, 3.10722, 3.122973, 3.118454, 3.138665, 
    3.12506, 3.149182, 3.135412, 3.137563, 3.124612, 3.046819, 3.061456, 
    3.045953, 3.048037, 3.047101, 3.035752, 3.030043, 3.018116, 3.020279, 
    3.029041, 3.048974, 3.042197, 3.059299, 3.058912, 3.078032, 3.0694, 
    3.101668, 3.092472, 3.118642, 3.112137, 3.118336, 3.116456, 3.118361, 
    3.108824, 3.112907, 3.104525, 3.071015, 3.080839, 3.051609, 3.03413, 
    3.022564, 3.014375, 3.015532, 3.017737, 3.029092, 3.039797, 3.047973, 
    3.053451, 3.058856, 3.075258, 3.083966, 3.103529, 3.099993, 3.105932, 
    3.11149, 3.120837, 3.119297, 3.12342, 3.10578, 3.117495, 3.097979, 
    3.103423, 3.060325, 3.044024, 3.037113, 3.031075, 3.016421, 3.026535, 
    3.022545, 3.032045, 3.038092, 3.0351, 3.053601, 3.046399, 3.084483, 
    3.068036, 3.110842, 3.100718, 3.113245, 3.106904, 3.117775, 3.10799, 
    3.124956, 3.128659, 3.126128, 3.135859, 3.107448, 3.118336, 3.035017, 
    3.035504, 3.037778, 3.027793, 3.027183, 3.018056, 3.026177, 3.029639, 
    3.038443, 3.043659, 3.048624, 3.059561, 3.071808, 3.088996, 3.101388, 
    3.109545, 3.104595, 3.108965, 3.104075, 3.101715, 3.12727, 3.112945, 
    3.134458, 3.133265, 3.123518, 3.133399, 3.035847, 3.03304, 3.02331, 
    3.030923, 3.017064, 3.024815, 3.029279, 3.046549, 3.050353, 3.053883, 
    3.060865, 3.069842, 3.085635, 3.099426, 3.111814, 3.110916, 3.111232, 
    3.11397, 3.10719, 3.115085, 3.116411, 3.112944, 3.133105, 3.127336, 
    3.13324, 3.129482, 3.033952, 3.038677, 3.036123, 3.040927, 3.037542, 
    3.052613, 3.057142, 3.078402, 3.069665, 3.08358, 3.071076, 3.073289, 
    3.084033, 3.071751, 3.098664, 3.080398, 3.114077, 3.096081, 3.115191, 
    3.111761, 3.117442, 3.122537, 3.128956, 3.140825, 3.138074, 3.148019, 
    3.045731, 3.051877, 3.051336, 3.057778, 3.062548, 3.072906, 3.089573, 
    3.083298, 3.094826, 3.097143, 3.079633, 3.090375, 3.055996, 3.061531, 
    3.058235, 3.046215, 3.084743, 3.064926, 3.101592, 3.090803, 3.12181, 
    3.106567, 3.13656, 3.149445, 3.161612, 3.17587, 3.055236, 3.051055, 
    3.058545, 3.068928, 3.078586, 3.09146, 3.09278, 3.095196, 3.101463, 
    3.106663, 3.09596, 3.107946, 3.062815, 3.086467, 3.049475, 3.06058, 
    3.068315, 3.06492, 3.082582, 3.086755, 3.103755, 3.094959, 3.146261, 
    3.123613, 3.18676, 3.169019, 3.049595, 3.055222, 3.074863, 3.065506, 
    3.092321, 3.098947, 3.104339, 3.111031, 3.111755, 3.115726, 3.109221, 
    3.115469, 3.091487, 3.102347, 3.072614, 3.079831, 3.076509, 3.072869, 
    3.084115, 3.09613, 3.096387, 3.100247, 3.110927, 3.09243, 3.149191, 
    3.11427, 3.061366, 3.07224, 3.073796, 3.069579, 3.098283, 3.08786, 
    3.115629, 3.108243, 3.120353, 3.114331, 3.113445, 3.105726, 3.100821, 
    3.088337, 3.078206, 3.07019, 3.072053, 3.080863, 3.096866, 3.11182, 
    3.108589, 3.119431, 3.090371, 3.102734, 3.097951, 3.110242, 3.083131, 
    3.1063, 3.077212, 3.079761, 3.087653, 3.103573, 3.107016, 3.110672, 
    3.108416, 3.097273, 3.095429, 3.087461, 3.085263, 3.079206, 3.074197, 
    3.078773, 3.083584, 3.097278, 3.10949, 3.12261, 3.125827, 3.141217, 
    3.128683, 3.149386, 3.131776, 3.162307, 3.107611, 3.131261, 3.088013, 
    3.092743, 3.101311, 3.120512, 3.110185, 3.122266, 3.095357, 3.081167, 
    3.077504, 3.070677, 3.07766, 3.077092, 3.083784, 3.081632, 3.097733, 
    3.089077, 3.113423, 3.122171, 3.146975, 3.162252, 3.177862, 3.184771, 
    3.186876, 3.187756,
  2.8934, 2.908718, 2.905735, 2.918126, 2.911247, 2.919368, 2.8965, 2.909328, 
    2.901133, 2.894776, 2.942291, 2.918679, 2.966968, 2.951796, 2.989996, 
    2.964604, 2.994977, 2.989283, 3.006443, 3.001519, 3.023555, 3.008718, 
    3.035027, 3.020006, 3.022352, 3.008229, 2.923418, 2.939344, 2.922477, 
    2.924743, 2.923726, 2.911389, 2.905188, 2.892231, 2.89458, 2.904098, 
    2.925763, 2.918394, 2.936991, 2.93657, 2.95738, 2.947983, 2.983129, 
    2.973107, 3.001724, 2.994637, 3.001391, 2.999342, 3.001418, 2.99103, 
    2.995477, 2.986254, 2.949741, 2.960437, 2.928627, 2.90963, 2.897062, 
    2.88817, 2.889426, 2.891821, 2.904154, 2.915785, 2.924673, 2.93063, 
    2.936509, 2.954363, 2.963844, 2.98516, 2.981303, 2.987838, 2.993933, 
    3.004116, 3.002438, 3.006931, 2.987664, 3.000475, 2.979108, 2.985042, 
    2.938113, 2.92038, 2.912871, 2.906308, 2.890391, 2.901376, 2.897042, 
    2.90736, 2.913932, 2.91068, 2.930793, 2.922961, 2.964406, 2.946499, 
    2.993227, 2.982094, 2.995845, 2.988929, 3.000781, 2.990121, 3.008605, 
    3.012642, 3.009882, 3.020492, 2.989531, 3.001392, 2.910589, 2.911119, 
    2.91359, 2.902742, 2.90208, 2.892167, 2.900986, 2.904748, 2.914313, 
    2.919983, 2.925381, 2.937276, 2.950605, 2.969321, 2.982824, 2.991815, 
    2.986332, 2.991183, 2.985753, 2.98318, 3.011129, 2.995519, 3.018964, 
    3.017663, 3.007038, 3.017809, 2.911492, 2.908442, 2.897872, 2.906141, 
    2.891089, 2.899508, 2.904357, 2.923126, 2.927261, 2.931101, 2.938695, 
    2.948463, 2.965661, 2.980686, 2.994285, 2.993307, 2.993652, 2.996635, 
    2.98925, 2.997849, 2.999294, 2.995517, 3.017488, 3.011198, 3.017635, 
    3.013538, 2.909433, 2.914568, 2.911792, 2.917013, 2.913335, 2.929721, 
    2.934647, 2.957785, 2.948271, 2.963422, 2.949807, 2.952216, 2.963919, 
    2.950541, 2.979857, 2.959959, 2.996751, 2.977044, 2.997965, 2.994228, 
    3.000417, 3.005969, 3.012965, 3.025908, 3.022907, 3.033756, 2.922235, 
    2.92892, 2.92833, 2.935336, 2.940526, 2.951799, 2.969949, 2.963114, 
    2.975671, 2.978198, 2.959123, 2.970824, 2.933399, 2.939422, 2.935834, 
    2.922762, 2.964689, 2.943115, 2.983047, 2.971289, 3.005177, 2.988552, 
    3.021256, 3.035316, 3.048593, 3.064171, 2.932572, 2.928024, 2.93617, 
    2.94747, 2.957983, 2.972005, 2.973442, 2.976076, 2.982906, 2.988658, 
    2.97691, 2.990073, 2.940821, 2.966567, 2.926307, 2.938387, 2.946803, 
    2.943108, 2.962333, 2.966879, 2.985405, 2.975817, 3.031842, 3.007144, 
    3.076072, 3.056685, 2.926437, 2.932556, 2.95393, 2.943745, 2.972943, 
    2.980164, 2.986044, 2.993434, 2.994222, 2.998548, 2.991461, 2.998267, 
    2.972035, 2.983869, 2.95148, 2.959338, 2.955721, 2.951757, 2.964004, 
    2.977095, 2.977374, 2.981581, 2.993329, 2.973061, 3.035043, 2.996969, 
    2.93924, 2.951076, 2.952768, 2.948177, 2.979439, 2.968083, 2.998442, 
    2.990397, 3.003588, 2.997027, 2.996063, 2.987604, 2.982206, 2.968603, 
    2.957569, 2.948842, 2.95087, 2.960463, 2.977897, 2.994293, 2.990776, 
    3.002584, 2.970818, 2.984292, 2.979079, 2.992574, 2.962933, 2.988258, 
    2.956486, 2.959261, 2.967858, 2.985208, 2.989055, 2.993043, 2.990585, 
    2.97834, 2.97633, 2.967648, 2.965255, 2.958657, 2.953203, 2.958186, 
    2.963426, 2.978345, 2.991755, 3.006048, 3.009554, 3.026341, 3.012671, 
    3.035257, 3.016049, 3.049359, 2.989712, 3.015483, 2.968249, 2.973402, 
    2.982742, 3.003765, 2.992512, 3.005675, 2.976251, 2.960794, 2.956804, 
    2.949373, 2.956974, 2.956355, 2.963642, 2.961299, 2.978841, 2.969408, 
    2.996039, 3.005571, 3.032618, 3.049295, 3.066344, 3.073896, 3.076197, 
    3.07716,
  2.944195, 2.960307, 2.957167, 2.970212, 2.962969, 2.971521, 2.947454, 
    2.960949, 2.952327, 2.945641, 2.995688, 2.970795, 3.021753, 3.005721, 
    3.04615, 3.019253, 3.051601, 3.045369, 3.06416, 3.058765, 3.082829, 
    3.066653, 3.095021, 3.079031, 3.081551, 3.066118, 2.975787, 2.992579, 
    2.974796, 2.977184, 2.976111, 2.963119, 2.956593, 2.942966, 2.945435, 
    2.955445, 2.978258, 2.970494, 2.990096, 2.989651, 3.011619, 3.001695, 
    3.038851, 3.028245, 3.05899, 3.05123, 3.058625, 3.056381, 3.058655, 
    3.047281, 3.052149, 3.042159, 3.003551, 3.014849, 2.981277, 2.961267, 
    2.948045, 2.938697, 2.940017, 2.942535, 2.955504, 2.967746, 2.977109, 
    2.983388, 2.989588, 3.008433, 3.01845, 3.041, 3.036917, 3.043836, 
    3.050459, 3.06161, 3.059772, 3.064695, 3.043653, 3.057622, 3.034594, 
    3.040876, 2.991281, 2.972586, 2.964679, 2.957771, 2.941032, 2.952582, 
    2.948024, 2.958878, 2.965796, 2.962372, 2.98356, 2.975306, 3.019045, 
    3.000129, 3.049685, 3.037755, 3.052552, 3.044992, 3.057957, 3.046286, 
    3.066529, 3.070955, 3.06793, 3.079564, 3.045641, 3.058626, 2.962276, 
    2.962835, 2.965436, 2.954019, 2.953322, 2.942898, 2.952171, 2.956129, 
    2.966197, 2.972168, 2.977855, 2.990396, 3.004464, 3.024241, 3.038527, 
    3.04814, 3.042241, 3.047448, 3.041628, 3.038904, 3.069296, 3.052195, 
    3.077888, 3.076461, 3.064812, 3.076621, 2.963227, 2.960016, 2.948897, 
    2.957595, 2.941765, 2.950617, 2.955718, 2.975479, 2.979837, 2.983884, 
    2.991893, 3.002202, 3.02037, 3.036265, 3.050844, 3.049773, 3.05015, 
    3.053416, 3.045333, 3.054745, 3.056329, 3.052192, 3.076269, 3.069372, 
    3.07643, 3.071937, 2.961059, 2.966465, 2.963543, 2.96904, 2.965167, 
    2.98243, 2.987624, 3.012047, 3.001999, 3.018004, 3.003621, 3.006165, 
    3.01853, 3.004396, 3.035387, 3.014344, 3.053543, 3.03241, 3.054873, 
    3.050781, 3.057558, 3.063641, 3.071309, 3.085329, 3.08214, 3.09367, 
    2.974541, 2.981585, 2.980963, 2.988351, 2.993825, 3.005724, 3.024905, 
    3.017678, 3.030957, 3.033631, 3.01346, 3.02583, 2.986308, 2.99266, 
    2.988876, 2.975096, 3.019343, 2.996557, 3.038764, 3.026321, 3.062773, 
    3.044593, 3.080386, 3.09533, 3.109456, 3.126053, 2.985435, 2.980641, 
    2.98923, 3.001154, 3.012256, 3.027079, 3.028599, 3.031386, 3.038614, 
    3.044704, 3.032268, 3.046233, 2.994138, 3.021328, 2.978832, 2.991569, 
    3.000449, 2.996549, 3.016853, 3.021658, 3.041261, 3.031111, 3.091635, 
    3.064929, 3.138747, 3.118075, 2.978968, 2.985419, 3.007975, 2.997222, 
    3.028071, 3.035712, 3.041936, 3.049913, 3.050774, 3.055511, 3.047753, 
    3.055204, 3.027111, 3.039634, 3.005387, 3.013688, 3.009866, 3.00568, 
    3.018619, 3.032464, 3.032759, 3.037212, 3.049799, 3.028196, 3.095041, 
    3.053783, 2.992468, 3.004961, 3.006747, 3.001899, 3.034945, 3.022931, 
    3.055395, 3.046588, 3.061031, 3.053846, 3.05279, 3.043588, 3.037874, 
    3.023481, 3.011819, 3.002602, 3.004743, 3.014876, 3.033313, 3.050853, 
    3.047003, 3.059931, 3.025824, 3.040081, 3.034564, 3.048971, 3.017487, 
    3.044282, 3.010675, 3.013607, 3.022693, 3.041052, 3.045126, 3.049484, 
    3.046794, 3.033782, 3.031654, 3.022471, 3.019942, 3.012968, 3.007207, 
    3.01247, 3.018008, 3.033786, 3.048075, 3.063728, 3.067569, 3.085789, 
    3.070988, 3.095268, 3.074693, 3.110273, 3.04584, 3.074071, 3.023106, 
    3.028557, 3.038441, 3.061227, 3.048903, 3.063319, 3.031571, 3.015227, 
    3.01101, 3.003162, 3.01119, 3.010536, 3.018236, 3.01576, 3.034312, 
    3.024333, 3.052764, 3.063205, 3.09246, 3.110204, 3.12837, 3.136425, 
    3.13888, 3.139908,
  2.969919, 2.988319, 2.984731, 2.999653, 2.991363, 3.001151, 2.973637, 
    2.989053, 2.9792, 2.971569, 3.028875, 3.00032, 3.058885, 3.040413, 
    3.087081, 3.056003, 3.093395, 3.086177, 3.107961, 3.1017, 3.129779, 
    3.110856, 3.144458, 3.125246, 3.128242, 3.110234, 3.006038, 3.025303, 
    3.004902, 3.007638, 3.00641, 2.991535, 2.984074, 2.968517, 2.971334, 
    2.982763, 3.00887, 2.999975, 3.022451, 3.021941, 3.047204, 3.035781, 
    3.078634, 3.066378, 3.101961, 3.092964, 3.101538, 3.098935, 3.101572, 
    3.08839, 3.094029, 3.082461, 3.037917, 3.050925, 3.012331, 2.989418, 
    2.974312, 2.96365, 2.965155, 2.968025, 2.98283, 2.99683, 3.007553, 
    3.014753, 3.021868, 3.043535, 3.055076, 3.081121, 3.076398, 3.084402, 
    3.092071, 3.105001, 3.102868, 3.108582, 3.08419, 3.100375, 3.073713, 
    3.080977, 3.023812, 3.002371, 2.99332, 2.98542, 2.966312, 2.979492, 
    2.974288, 2.986686, 2.994597, 2.990681, 3.01495, 3.005486, 3.055762, 
    3.03398, 3.091175, 3.077367, 3.094496, 3.08574, 3.100763, 3.087238, 
    3.110712, 3.115854, 3.112339, 3.125865, 3.086491, 3.101539, 2.990572, 
    2.99121, 2.994185, 2.981134, 2.980337, 2.96844, 2.979023, 2.983544, 
    2.995056, 3.001893, 3.008409, 3.022796, 3.038966, 3.061756, 3.078259, 
    3.089385, 3.082556, 3.088584, 3.081847, 3.078696, 3.113926, 3.094082, 
    3.123915, 3.122255, 3.108719, 3.122442, 2.991658, 2.987987, 2.975285, 
    2.985219, 2.967148, 2.977248, 2.983075, 3.005685, 3.01068, 3.015322, 
    3.024515, 3.036364, 3.057291, 3.075644, 3.092517, 3.091277, 3.091714, 
    3.095498, 3.086135, 3.097039, 3.098874, 3.094079, 3.122033, 3.114014, 
    3.12222, 3.116995, 2.989179, 2.995363, 2.99202, 2.998311, 2.993878, 
    3.013654, 3.019614, 3.047697, 3.036131, 3.054562, 3.037996, 3.040924, 
    3.055169, 3.038888, 3.07463, 3.050344, 3.095645, 3.071189, 3.097186, 
    3.092444, 3.1003, 3.107358, 3.116265, 3.132787, 3.128951, 3.14283, 
    3.00461, 3.012685, 3.011971, 3.020447, 3.026735, 3.040416, 3.062522, 
    3.054186, 3.069511, 3.072599, 3.049325, 3.06359, 3.018103, 3.025396, 
    3.02105, 3.005247, 3.056106, 3.029874, 3.078533, 3.064157, 3.106351, 
    3.085278, 3.126842, 3.14483, 3.161399, 3.180834, 3.017102, 3.011602, 
    3.021457, 3.035159, 3.047938, 3.065032, 3.066787, 3.070005, 3.07836, 
    3.085407, 3.071025, 3.087177, 3.027093, 3.058396, 3.009527, 3.024142, 
    3.034348, 3.029865, 3.053235, 3.058775, 3.081422, 3.069688, 3.140379, 
    3.108853, 3.195733, 3.171485, 3.009684, 3.017082, 3.043007, 3.030638, 
    3.066177, 3.075005, 3.082203, 3.091438, 3.092437, 3.097927, 3.088937, 
    3.09757, 3.065068, 3.07954, 3.040029, 3.049588, 3.045185, 3.040366, 
    3.05527, 3.071251, 3.071592, 3.076739, 3.091307, 3.066322, 3.144481, 
    3.095924, 3.025175, 3.039538, 3.041595, 3.036016, 3.074118, 3.060244, 
    3.097792, 3.087587, 3.10433, 3.095996, 3.094773, 3.084115, 3.077504, 
    3.060879, 3.047435, 3.036824, 3.039287, 3.050956, 3.072232, 3.092528, 
    3.088068, 3.103053, 3.063583, 3.080058, 3.073678, 3.090348, 3.053965, 
    3.084919, 3.046116, 3.049493, 3.05997, 3.08118, 3.085895, 3.090942, 
    3.087826, 3.072774, 3.070316, 3.059714, 3.056796, 3.048758, 3.042123, 
    3.048184, 3.054567, 3.072779, 3.08931, 3.107459, 3.11192, 3.133341, 
    3.115892, 3.144755, 3.120199, 3.162355, 3.086722, 3.119477, 3.060447, 
    3.066738, 3.078161, 3.104556, 3.090269, 3.106985, 3.070219, 3.051361, 
    3.046503, 3.037468, 3.04671, 3.045957, 3.05483, 3.051975, 3.073386, 
    3.061862, 3.094742, 3.106852, 3.141373, 3.162275, 3.18355, 3.193005, 
    3.19589, 3.197097,
  3.25474, 3.278216, 3.273628, 3.292736, 3.282112, 3.294659, 3.259475, 
    3.279155, 3.266567, 3.25684, 3.329906, 3.293593, 3.36768, 3.344389, 
    3.403475, 3.364037, 3.411532, 3.402323, 3.430178, 3.422154, 3.458264, 
    3.433893, 3.477266, 3.452412, 3.456279, 3.433096, 3.300937, 3.32543, 
    3.299477, 3.302995, 3.301415, 3.282331, 3.272789, 3.252956, 3.256541, 
    3.271114, 3.304579, 3.29315, 3.321861, 3.321223, 3.352937, 3.338568, 
    3.39272, 3.377162, 3.422488, 3.410982, 3.421946, 3.418614, 3.42199, 
    3.405144, 3.412343, 3.397589, 3.341251, 3.357627, 3.309035, 3.279622, 
    3.260334, 3.246769, 3.248681, 3.252331, 3.2712, 3.289115, 3.302885, 
    3.312154, 3.321131, 3.348316, 3.362867, 3.395883, 3.389878, 3.400062, 
    3.409841, 3.426383, 3.42365, 3.430976, 3.399791, 3.420457, 3.386467, 
    3.3957, 3.323564, 3.296226, 3.284618, 3.27451, 3.250152, 3.266939, 
    3.260304, 3.276128, 3.286254, 3.281238, 3.312408, 3.300228, 3.363733, 
    3.336308, 3.408698, 3.391109, 3.412939, 3.401766, 3.420953, 3.403676, 
    3.433709, 3.440316, 3.435799, 3.453212, 3.402723, 3.421947, 3.281098, 
    3.281915, 3.285726, 3.269035, 3.268018, 3.252858, 3.26634, 3.272112, 
    3.286842, 3.295611, 3.303986, 3.322293, 3.342571, 3.371311, 3.392244, 
    3.406413, 3.397711, 3.405391, 3.396808, 3.392798, 3.437838, 3.41241, 
    3.450697, 3.448557, 3.43115, 3.448798, 3.282489, 3.277791, 3.261574, 
    3.274253, 3.251215, 3.264076, 3.271513, 3.300484, 3.306908, 3.312887, 
    3.324444, 3.339301, 3.365664, 3.388919, 3.410411, 3.408828, 3.409385, 
    3.41422, 3.402269, 3.416189, 3.418537, 3.412406, 3.44827, 3.437951, 
    3.448511, 3.441785, 3.279317, 3.287235, 3.282952, 3.291014, 3.285331, 
    3.310738, 3.318314, 3.353558, 3.339008, 3.362218, 3.341352, 3.345032, 
    3.362983, 3.342472, 3.387631, 3.356895, 3.414408, 3.383263, 3.416378, 
    3.410318, 3.420361, 3.429405, 3.440845, 3.46215, 3.457194, 3.475154, 
    3.299102, 3.30949, 3.308571, 3.319355, 3.327223, 3.344393, 3.37228, 
    3.361742, 3.381134, 3.385053, 3.35561, 3.373632, 3.316426, 3.325547, 
    3.32011, 3.29992, 3.364168, 3.331157, 3.392592, 3.37435, 3.428113, 
    3.401177, 3.454472, 3.477748, 3.499923, 3.526196, 3.315175, 3.308096, 
    3.320618, 3.337787, 3.353861, 3.375458, 3.377681, 3.381761, 3.392371, 
    3.401342, 3.383055, 3.403597, 3.327673, 3.367061, 3.305425, 3.323977, 
    3.33677, 3.331146, 3.360542, 3.367541, 3.396266, 3.381359, 3.471977, 
    3.431324, 3.546063, 3.513536, 3.305627, 3.31515, 3.347653, 3.332115, 
    3.376908, 3.388107, 3.397261, 3.409034, 3.410308, 3.417325, 3.405841, 
    3.416869, 3.375504, 3.393872, 3.343906, 3.355941, 3.350394, 3.34433, 
    3.363112, 3.383342, 3.383774, 3.390311, 3.408866, 3.377091, 3.477296, 
    3.414763, 3.32527, 3.34329, 3.345875, 3.338864, 3.386981, 3.369398, 
    3.417153, 3.404121, 3.425522, 3.414856, 3.413292, 3.399696, 3.391283, 
    3.370201, 3.353227, 3.339879, 3.342974, 3.357667, 3.384586, 3.410425, 
    3.404733, 3.423887, 3.373622, 3.394531, 3.386421, 3.407641, 3.361464, 
    3.40072, 3.351566, 3.355822, 3.369051, 3.395959, 3.401963, 3.408401, 
    3.404425, 3.385274, 3.382155, 3.368728, 3.365039, 3.354895, 3.34654, 
    3.354172, 3.362223, 3.385281, 3.406317, 3.429534, 3.435261, 3.462866, 
    3.440366, 3.477651, 3.445909, 3.501211, 3.403017, 3.444978, 3.369654, 
    3.377619, 3.392118, 3.425813, 3.407541, 3.428927, 3.382033, 3.358178, 
    3.352053, 3.340688, 3.352314, 3.351366, 3.362556, 3.358952, 3.386052, 
    3.371444, 3.413254, 3.428756, 3.473264, 3.501102, 3.529882, 3.542461, 
    3.54627, 3.547865,
  3.812393, 3.852924, 3.844952, 3.878324, 3.859713, 3.881707, 3.820515, 
    3.854559, 3.83273, 3.815992, 3.945428, 3.879831, 4.016907, 3.972589, 
    4.084889, 4.009922, 4.100391, 4.08268, 4.136661, 4.120984, 4.192374, 
    4.143956, 4.230835, 4.180657, 4.188393, 4.142387, 3.892786, 3.937095, 
    3.890205, 3.896428, 3.893631, 3.860096, 3.843497, 3.80934, 3.815479, 
    3.840594, 3.899235, 3.879052, 3.93047, 3.929288, 3.988761, 3.961638, 
    4.064354, 4.034963, 4.121634, 4.099329, 4.12058, 4.114101, 4.120664, 
    4.088093, 4.101956, 4.073629, 3.96668, 3.997681, 3.907147, 3.855371, 
    3.821991, 3.798779, 3.802038, 3.808271, 3.840742, 3.871965, 3.896233, 
    3.912702, 3.929118, 3.980006, 4.007683, 4.070376, 4.058958, 4.078353, 
    4.097129, 4.129234, 4.123899, 4.138225, 4.077835, 4.117682, 4.052496, 
    4.070027, 3.933629, 3.884468, 3.86409, 3.846481, 3.804549, 3.833373, 
    3.82194, 3.849291, 3.866952, 3.858189, 3.913155, 3.891532, 4.00934, 
    3.957397, 4.094926, 4.061294, 4.103108, 4.081614, 4.118647, 4.085274, 
    4.143593, 4.15662, 4.147705, 4.182254, 4.083448, 4.120581, 3.857945, 
    3.85937, 3.866028, 3.836994, 3.835237, 3.809173, 3.832339, 3.842322, 
    3.867982, 3.883384, 3.898182, 3.931272, 3.969163, 4.023889, 4.06345, 
    4.09053, 4.073862, 4.088568, 4.072139, 4.064504, 4.151726, 4.102087, 
    4.177233, 4.172968, 4.138568, 4.173448, 3.860372, 3.852184, 3.824124, 
    3.846035, 3.806363, 3.828434, 3.841284, 3.891984, 3.903368, 3.91401, 
    3.935263, 3.963014, 4.01304, 4.05714, 4.098228, 4.095177, 4.096251, 
    4.105585, 4.082578, 4.109397, 4.113951, 4.102079, 4.172398, 4.151948, 
    4.172878, 4.159524, 3.85484, 3.86867, 3.86118, 3.875299, 3.865339, 
    3.910178, 3.923903, 3.989941, 3.962463, 4.006441, 3.966868, 3.973802, 
    4.007906, 3.968978, 4.0547, 3.996286, 4.105948, 4.046445, 4.109763, 
    4.098048, 4.117496, 4.135146, 4.157666, 4.200188, 4.190227, 4.226528, 
    3.889542, 3.907957, 3.906323, 3.92583, 3.940431, 3.972598, 4.025756, 
    4.005533, 4.042431, 4.049824, 3.99384, 4.028343, 3.920414, 3.937314, 
    3.927225, 3.890987, 4.010172, 3.947763, 4.064112, 4.029688, 4.132617, 
    4.080487, 4.184773, 4.231818, 4.277538, 4.332246, 3.918106, 3.905478, 
    3.928166, 3.960172, 3.990517, 4.031764, 4.035937, 4.043613, 4.063693, 
    4.080802, 4.046052, 4.085124, 3.941267, 4.015718, 3.900735, 3.934397, 
    3.958264, 3.947742, 4.003239, 4.01664, 4.071107, 4.042855, 4.220065, 
    4.138907, 4.374605, 4.306057, 3.901093, 3.918061, 3.978752, 3.949552, 
    4.034485, 4.055602, 4.073004, 4.095573, 4.09803, 4.111598, 4.089432, 
    4.110715, 4.031851, 4.066545, 3.971679, 3.994471, 3.983939, 3.972478, 
    4.008152, 4.046594, 4.047409, 4.05978, 4.09525, 4.03483, 4.230896, 
    4.106637, 3.936798, 3.970517, 3.975393, 3.962193, 4.053471, 4.020208, 
    4.111266, 4.086128, 4.127552, 4.106816, 4.103791, 4.077653, 4.061625, 
    4.021753, 3.989313, 3.964099, 3.969922, 3.997757, 4.048943, 4.098255, 
    4.087304, 4.124361, 4.028325, 4.067799, 4.052412, 4.092893, 4.005001, 
    4.079612, 3.986161, 3.994245, 4.019541, 4.070521, 4.081992, 4.094354, 
    4.086712, 4.050242, 4.044355, 4.018919, 4.011842, 3.99248, 3.976649, 
    3.991108, 4.006452, 4.050256, 4.090347, 4.1354, 4.146646, 4.201631, 
    4.156718, 4.231621, 4.167703, 4.280221, 4.084012, 4.165855, 4.020701, 
    4.03582, 4.06321, 4.128119, 4.0927, 4.134209, 4.044125, 3.99873, 
    3.987085, 3.965621, 3.98758, 3.985781, 4.007088, 4.000206, 4.051713, 
    4.024145, 4.103716, 4.133875, 4.222682, 4.279996, 4.339895, 4.366773, 
    4.375056, 4.378533,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24814.43, 24834.87, 24830.86, 24847.59, 24838.27, 24849.28, 24818.54, 
    24835.69, 24824.71, 24816.25, 24880.8, 24848.34, 24915.59, 24894.08, 
    24948.58, 24912.21, 24956.05, 24947.52, 24973.43, 24965.93, 24999.9, 
    24976.92, 25017.98, 24994.36, 24998.02, 24976.17, 24854.8, 24876.72, 
    24853.52, 24856.62, 24855.22, 24838.47, 24830.13, 24812.89, 24815.99, 
    24828.67, 24858.01, 24847.95, 24873.46, 24872.88, 24901.95, 24888.74, 
    24938.65, 24924.35, 24966.25, 24955.54, 24965.74, 24962.63, 24965.78, 
    24950.13, 24956.8, 24943.14, 24891.2, 24906.28, 24861.95, 24836.1, 
    24819.29, 24807.53, 24809.19, 24812.35, 24828.74, 24844.41, 24856.52, 
    24864.7, 24872.8, 24897.69, 24911.13, 24941.56, 24936.03, 24945.42, 
    24954.48, 24969.88, 24967.33, 24974.18, 24945.17, 24964.35, 24932.89, 
    24941.4, 24875.02, 24850.66, 24840.47, 24831.63, 24810.46, 24825.03, 
    24819.26, 24833.04, 24841.9, 24837.51, 24864.93, 24854.18, 24911.93, 
    24886.66, 24953.42, 24937.16, 24957.36, 24947, 24964.81, 24948.77, 
    24976.74, 24982.95, 24978.7, 24995.12, 24947.89, 24965.74, 24837.39, 
    24838.1, 24841.44, 24826.86, 24825.97, 24812.8, 24824.51, 24829.54, 
    24842.42, 24850.12, 24857.49, 24873.86, 24892.41, 24918.96, 24938.21, 
    24951.3, 24943.25, 24950.36, 24942.42, 24938.72, 24980.62, 24956.87, 
    24992.74, 24990.71, 24974.34, 24990.94, 24838.61, 24834.5, 24820.36, 
    24831.41, 24811.38, 24822.54, 24829.02, 24854.4, 24860.07, 24865.35, 
    24875.82, 24889.41, 24913.72, 24935.14, 24955.01, 24953.54, 24954.06, 
    24958.55, 24947.47, 24960.38, 24962.56, 24956.86, 24990.44, 24980.72, 
    24990.67, 24984.33, 24835.83, 24842.76, 24839.01, 24846.08, 24841.09, 
    24863.45, 24870.24, 24902.53, 24889.14, 24910.53, 24891.29, 24894.67, 
    24911.24, 24892.32, 24933.96, 24905.61, 24958.72, 24929.95, 24960.55, 
    24954.92, 24964.26, 24972.71, 24983.45, 25003.58, 24998.88, 25015.96, 
    24853.19, 24862.35, 24861.54, 24871.18, 24878.36, 24894.09, 24919.87, 
    24910.09, 24927.99, 24931.59, 24904.42, 24921.12, 24868.52, 24876.83, 
    24871.87, 24853.91, 24912.34, 24881.95, 24938.53, 24921.78, 24971.5, 
    24946.46, 24996.31, 25018.44, 25039.72, 25065.06, 24867.38, 24861.12, 
    24872.33, 24888.02, 24902.8, 24922.79, 24924.83, 24928.57, 24938.33, 
    24946.61, 24929.75, 24948.7, 24878.77, 24915.02, 24858.76, 24875.39, 
    24887.09, 24881.94, 24908.98, 24915.46, 24941.92, 24928.2, 25012.93, 
    24974.51, 25084.57, 25052.9, 24858.94, 24867.36, 24897.08, 24882.83, 
    24924.12, 24934.4, 24942.84, 24953.73, 24954.91, 24961.43, 24950.77, 
    24961.01, 24922.83, 24939.71, 24893.64, 24904.72, 24899.61, 24894.03, 
    24911.36, 24930.02, 24930.41, 24936.43, 24953.57, 24924.29, 25018.01, 
    24959.05, 24876.57, 24893.07, 24895.45, 24889.01, 24933.36, 24917.19, 
    24961.27, 24949.18, 24969.08, 24959.14, 24957.68, 24945.09, 24937.32, 
    24917.93, 24902.22, 24889.94, 24892.78, 24906.32, 24931.16, 24955.02, 
    24949.75, 24967.55, 24921.11, 24940.32, 24932.85, 24952.44, 24909.83, 
    24946.03, 24900.69, 24904.62, 24916.87, 24941.63, 24947.18, 24953.14, 
    24949.46, 24931.79, 24928.93, 24916.57, 24913.14, 24903.76, 24896.06, 
    24903.09, 24910.54, 24931.8, 24951.21, 24972.83, 24978.2, 25004.26, 
    24982.99, 25018.35, 24988.21, 25040.96, 24948.16, 24987.34, 24917.43, 
    24924.77, 24938.09, 24969.35, 24952.35, 24972.26, 24928.81, 24906.79, 
    24901.14, 24890.68, 24901.38, 24900.5, 24910.84, 24907.51, 24932.51, 
    24919.09, 24957.65, 24972.1, 25014.16, 25040.86, 25068.61, 25080.98, 
    25084.78, 25086.37 ;

 HCSOI =
  24814.43, 24834.87, 24830.86, 24847.59, 24838.27, 24849.28, 24818.54, 
    24835.69, 24824.71, 24816.25, 24880.8, 24848.34, 24915.59, 24894.08, 
    24948.58, 24912.21, 24956.05, 24947.52, 24973.43, 24965.93, 24999.9, 
    24976.92, 25017.98, 24994.36, 24998.02, 24976.17, 24854.8, 24876.72, 
    24853.52, 24856.62, 24855.22, 24838.47, 24830.13, 24812.89, 24815.99, 
    24828.67, 24858.01, 24847.95, 24873.46, 24872.88, 24901.95, 24888.74, 
    24938.65, 24924.35, 24966.25, 24955.54, 24965.74, 24962.63, 24965.78, 
    24950.13, 24956.8, 24943.14, 24891.2, 24906.28, 24861.95, 24836.1, 
    24819.29, 24807.53, 24809.19, 24812.35, 24828.74, 24844.41, 24856.52, 
    24864.7, 24872.8, 24897.69, 24911.13, 24941.56, 24936.03, 24945.42, 
    24954.48, 24969.88, 24967.33, 24974.18, 24945.17, 24964.35, 24932.89, 
    24941.4, 24875.02, 24850.66, 24840.47, 24831.63, 24810.46, 24825.03, 
    24819.26, 24833.04, 24841.9, 24837.51, 24864.93, 24854.18, 24911.93, 
    24886.66, 24953.42, 24937.16, 24957.36, 24947, 24964.81, 24948.77, 
    24976.74, 24982.95, 24978.7, 24995.12, 24947.89, 24965.74, 24837.39, 
    24838.1, 24841.44, 24826.86, 24825.97, 24812.8, 24824.51, 24829.54, 
    24842.42, 24850.12, 24857.49, 24873.86, 24892.41, 24918.96, 24938.21, 
    24951.3, 24943.25, 24950.36, 24942.42, 24938.72, 24980.62, 24956.87, 
    24992.74, 24990.71, 24974.34, 24990.94, 24838.61, 24834.5, 24820.36, 
    24831.41, 24811.38, 24822.54, 24829.02, 24854.4, 24860.07, 24865.35, 
    24875.82, 24889.41, 24913.72, 24935.14, 24955.01, 24953.54, 24954.06, 
    24958.55, 24947.47, 24960.38, 24962.56, 24956.86, 24990.44, 24980.72, 
    24990.67, 24984.33, 24835.83, 24842.76, 24839.01, 24846.08, 24841.09, 
    24863.45, 24870.24, 24902.53, 24889.14, 24910.53, 24891.29, 24894.67, 
    24911.24, 24892.32, 24933.96, 24905.61, 24958.72, 24929.95, 24960.55, 
    24954.92, 24964.26, 24972.71, 24983.45, 25003.58, 24998.88, 25015.96, 
    24853.19, 24862.35, 24861.54, 24871.18, 24878.36, 24894.09, 24919.87, 
    24910.09, 24927.99, 24931.59, 24904.42, 24921.12, 24868.52, 24876.83, 
    24871.87, 24853.91, 24912.34, 24881.95, 24938.53, 24921.78, 24971.5, 
    24946.46, 24996.31, 25018.44, 25039.72, 25065.06, 24867.38, 24861.12, 
    24872.33, 24888.02, 24902.8, 24922.79, 24924.83, 24928.57, 24938.33, 
    24946.61, 24929.75, 24948.7, 24878.77, 24915.02, 24858.76, 24875.39, 
    24887.09, 24881.94, 24908.98, 24915.46, 24941.92, 24928.2, 25012.93, 
    24974.51, 25084.57, 25052.9, 24858.94, 24867.36, 24897.08, 24882.83, 
    24924.12, 24934.4, 24942.84, 24953.73, 24954.91, 24961.43, 24950.77, 
    24961.01, 24922.83, 24939.71, 24893.64, 24904.72, 24899.61, 24894.03, 
    24911.36, 24930.02, 24930.41, 24936.43, 24953.57, 24924.29, 25018.01, 
    24959.05, 24876.57, 24893.07, 24895.45, 24889.01, 24933.36, 24917.19, 
    24961.27, 24949.18, 24969.08, 24959.14, 24957.68, 24945.09, 24937.32, 
    24917.93, 24902.22, 24889.94, 24892.78, 24906.32, 24931.16, 24955.02, 
    24949.75, 24967.55, 24921.11, 24940.32, 24932.85, 24952.44, 24909.83, 
    24946.03, 24900.69, 24904.62, 24916.87, 24941.63, 24947.18, 24953.14, 
    24949.46, 24931.79, 24928.93, 24916.57, 24913.14, 24903.76, 24896.06, 
    24903.09, 24910.54, 24931.8, 24951.21, 24972.83, 24978.2, 25004.26, 
    24982.99, 25018.35, 24988.21, 25040.96, 24948.16, 24987.34, 24917.43, 
    24924.77, 24938.09, 24969.35, 24952.35, 24972.26, 24928.81, 24906.79, 
    24901.14, 24890.68, 24901.38, 24900.5, 24910.84, 24907.51, 24932.51, 
    24919.09, 24957.65, 24972.1, 25014.16, 25040.86, 25068.61, 25080.98, 
    25084.78, 25086.37 ;

 HEAT_FROM_AC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 HR =
  6.359163e-08, 6.387121e-08, 6.381686e-08, 6.404235e-08, 6.391726e-08, 
    6.406492e-08, 6.364831e-08, 6.388231e-08, 6.373293e-08, 6.36168e-08, 
    6.447997e-08, 6.405241e-08, 6.492405e-08, 6.465138e-08, 6.533632e-08, 
    6.488163e-08, 6.542801e-08, 6.53232e-08, 6.563863e-08, 6.554826e-08, 
    6.595173e-08, 6.568033e-08, 6.616087e-08, 6.588692e-08, 6.592978e-08, 
    6.567138e-08, 6.413845e-08, 6.442674e-08, 6.412137e-08, 6.416248e-08, 
    6.414403e-08, 6.391985e-08, 6.380688e-08, 6.357025e-08, 6.361321e-08, 
    6.3787e-08, 6.418097e-08, 6.404723e-08, 6.438426e-08, 6.437665e-08, 
    6.475187e-08, 6.458269e-08, 6.521333e-08, 6.503409e-08, 6.555204e-08, 
    6.542178e-08, 6.554592e-08, 6.550827e-08, 6.554641e-08, 6.535537e-08, 
    6.543722e-08, 6.526912e-08, 6.461438e-08, 6.480681e-08, 6.423289e-08, 
    6.38878e-08, 6.365858e-08, 6.349591e-08, 6.351891e-08, 6.356274e-08, 
    6.378801e-08, 6.399981e-08, 6.416121e-08, 6.426918e-08, 6.437556e-08, 
    6.469757e-08, 6.486799e-08, 6.524958e-08, 6.518071e-08, 6.529738e-08, 
    6.540882e-08, 6.559594e-08, 6.556514e-08, 6.564758e-08, 6.529429e-08, 
    6.552909e-08, 6.514148e-08, 6.52475e-08, 6.44045e-08, 6.40833e-08, 
    6.394681e-08, 6.38273e-08, 6.353659e-08, 6.373735e-08, 6.365821e-08, 
    6.384649e-08, 6.396612e-08, 6.390695e-08, 6.427213e-08, 6.413016e-08, 
    6.487809e-08, 6.455593e-08, 6.539582e-08, 6.519484e-08, 6.544399e-08, 
    6.531685e-08, 6.55347e-08, 6.533864e-08, 6.567826e-08, 6.575221e-08, 
    6.570168e-08, 6.58958e-08, 6.532778e-08, 6.554592e-08, 6.39053e-08, 
    6.391495e-08, 6.39599e-08, 6.376228e-08, 6.375019e-08, 6.356908e-08, 
    6.373023e-08, 6.379886e-08, 6.397305e-08, 6.40761e-08, 6.417405e-08, 
    6.438941e-08, 6.462994e-08, 6.496626e-08, 6.520787e-08, 6.536983e-08, 
    6.527052e-08, 6.53582e-08, 6.526018e-08, 6.521424e-08, 6.572451e-08, 
    6.543799e-08, 6.586788e-08, 6.584409e-08, 6.564954e-08, 6.584677e-08, 
    6.392172e-08, 6.386619e-08, 6.367338e-08, 6.382427e-08, 6.354936e-08, 
    6.370324e-08, 6.379173e-08, 6.413313e-08, 6.420814e-08, 6.427769e-08, 
    6.441505e-08, 6.459135e-08, 6.49006e-08, 6.516968e-08, 6.54153e-08, 
    6.539731e-08, 6.540364e-08, 6.545852e-08, 6.53226e-08, 6.548083e-08, 
    6.550739e-08, 6.543795e-08, 6.58409e-08, 6.572579e-08, 6.584358e-08, 
    6.576862e-08, 6.388424e-08, 6.397768e-08, 6.392719e-08, 6.402214e-08, 
    6.395525e-08, 6.425269e-08, 6.434187e-08, 6.475913e-08, 6.458788e-08, 
    6.486043e-08, 6.461556e-08, 6.465896e-08, 6.486933e-08, 6.462879e-08, 
    6.515485e-08, 6.479821e-08, 6.546065e-08, 6.510453e-08, 6.548296e-08, 
    6.541424e-08, 6.552803e-08, 6.562993e-08, 6.575814e-08, 6.59947e-08, 
    6.593991e-08, 6.613774e-08, 6.411698e-08, 6.423819e-08, 6.422751e-08, 
    6.435434e-08, 6.444814e-08, 6.465145e-08, 6.497752e-08, 6.485489e-08, 
    6.508e-08, 6.512519e-08, 6.47832e-08, 6.499319e-08, 6.431929e-08, 
    6.442818e-08, 6.436335e-08, 6.412655e-08, 6.488316e-08, 6.449487e-08, 
    6.521186e-08, 6.500152e-08, 6.56154e-08, 6.531011e-08, 6.590976e-08, 
    6.616612e-08, 6.640736e-08, 6.668932e-08, 6.430432e-08, 6.422197e-08, 
    6.436942e-08, 6.457343e-08, 6.476271e-08, 6.501435e-08, 6.504009e-08, 
    6.508724e-08, 6.520934e-08, 6.531201e-08, 6.510215e-08, 6.533775e-08, 
    6.445345e-08, 6.491686e-08, 6.419084e-08, 6.440948e-08, 6.456141e-08, 
    6.449476e-08, 6.484088e-08, 6.492246e-08, 6.525397e-08, 6.50826e-08, 
    6.610285e-08, 6.565147e-08, 6.690398e-08, 6.655396e-08, 6.41932e-08, 
    6.430404e-08, 6.46898e-08, 6.450625e-08, 6.503114e-08, 6.516034e-08, 
    6.526538e-08, 6.539964e-08, 6.541413e-08, 6.549368e-08, 6.536332e-08, 
    6.548853e-08, 6.501489e-08, 6.522654e-08, 6.46457e-08, 6.478708e-08, 
    6.472204e-08, 6.46507e-08, 6.487087e-08, 6.510545e-08, 6.511046e-08, 
    6.518567e-08, 6.539766e-08, 6.503327e-08, 6.616113e-08, 6.546461e-08, 
    6.44249e-08, 6.463841e-08, 6.466889e-08, 6.458619e-08, 6.514739e-08, 
    6.494405e-08, 6.549174e-08, 6.534372e-08, 6.558625e-08, 6.546573e-08, 
    6.5448e-08, 6.529321e-08, 6.519684e-08, 6.495338e-08, 6.475528e-08, 
    6.459818e-08, 6.463471e-08, 6.480727e-08, 6.51198e-08, 6.541545e-08, 
    6.535068e-08, 6.556781e-08, 6.499309e-08, 6.523408e-08, 6.514095e-08, 
    6.538381e-08, 6.485164e-08, 6.530484e-08, 6.47358e-08, 6.47857e-08, 
    6.494002e-08, 6.525044e-08, 6.53191e-08, 6.539243e-08, 6.534718e-08, 
    6.512773e-08, 6.509178e-08, 6.493626e-08, 6.489333e-08, 6.477483e-08, 
    6.467673e-08, 6.476636e-08, 6.486049e-08, 6.512782e-08, 6.536873e-08, 
    6.563138e-08, 6.569566e-08, 6.600256e-08, 6.575274e-08, 6.616501e-08, 
    6.581453e-08, 6.642122e-08, 6.533109e-08, 6.58042e-08, 6.494704e-08, 
    6.503938e-08, 6.520641e-08, 6.558949e-08, 6.538266e-08, 6.562454e-08, 
    6.509037e-08, 6.481324e-08, 6.474151e-08, 6.460773e-08, 6.474458e-08, 
    6.473344e-08, 6.486439e-08, 6.482231e-08, 6.51367e-08, 6.496782e-08, 
    6.544756e-08, 6.562262e-08, 6.611701e-08, 6.642009e-08, 6.672858e-08, 
    6.686479e-08, 6.690624e-08, 6.692357e-08 ;

 HR_vr =
  2.672496e-07, 2.679569e-07, 2.678195e-07, 2.683896e-07, 2.680734e-07, 
    2.684466e-07, 2.67393e-07, 2.679851e-07, 2.676072e-07, 2.673133e-07, 
    2.694946e-07, 2.68415e-07, 2.706135e-07, 2.699266e-07, 2.716504e-07, 
    2.705067e-07, 2.718807e-07, 2.716174e-07, 2.724095e-07, 2.721827e-07, 
    2.731948e-07, 2.725142e-07, 2.737187e-07, 2.730323e-07, 2.731398e-07, 
    2.724917e-07, 2.686323e-07, 2.693603e-07, 2.685892e-07, 2.686931e-07, 
    2.686465e-07, 2.680799e-07, 2.677943e-07, 2.671954e-07, 2.673042e-07, 
    2.67744e-07, 2.687398e-07, 2.684019e-07, 2.692529e-07, 2.692337e-07, 
    2.701798e-07, 2.697534e-07, 2.713412e-07, 2.708904e-07, 2.721922e-07, 
    2.71865e-07, 2.721768e-07, 2.720823e-07, 2.72178e-07, 2.716982e-07, 
    2.719038e-07, 2.714814e-07, 2.698333e-07, 2.703182e-07, 2.688709e-07, 
    2.67999e-07, 2.67419e-07, 2.670072e-07, 2.670654e-07, 2.671764e-07, 
    2.677466e-07, 2.682821e-07, 2.686898e-07, 2.689625e-07, 2.69231e-07, 
    2.700431e-07, 2.704723e-07, 2.714323e-07, 2.712591e-07, 2.715525e-07, 
    2.718325e-07, 2.723024e-07, 2.722251e-07, 2.72432e-07, 2.715447e-07, 
    2.721346e-07, 2.711605e-07, 2.714271e-07, 2.693042e-07, 2.68493e-07, 
    2.681482e-07, 2.678459e-07, 2.671102e-07, 2.676184e-07, 2.674181e-07, 
    2.678944e-07, 2.681969e-07, 2.680473e-07, 2.689699e-07, 2.686114e-07, 
    2.704978e-07, 2.69686e-07, 2.717998e-07, 2.712947e-07, 2.719208e-07, 
    2.716014e-07, 2.721487e-07, 2.716561e-07, 2.72509e-07, 2.726945e-07, 
    2.725677e-07, 2.730546e-07, 2.716288e-07, 2.721768e-07, 2.680431e-07, 
    2.680675e-07, 2.681812e-07, 2.676815e-07, 2.676509e-07, 2.671925e-07, 
    2.676003e-07, 2.67774e-07, 2.682144e-07, 2.684748e-07, 2.687223e-07, 
    2.692659e-07, 2.698726e-07, 2.707197e-07, 2.713275e-07, 2.717345e-07, 
    2.714849e-07, 2.717053e-07, 2.71459e-07, 2.713435e-07, 2.72625e-07, 
    2.719058e-07, 2.729846e-07, 2.729249e-07, 2.724369e-07, 2.729317e-07, 
    2.680846e-07, 2.679442e-07, 2.674565e-07, 2.678382e-07, 2.671425e-07, 
    2.675321e-07, 2.67756e-07, 2.686189e-07, 2.688083e-07, 2.68984e-07, 
    2.693306e-07, 2.697753e-07, 2.705544e-07, 2.712314e-07, 2.718488e-07, 
    2.718035e-07, 2.718195e-07, 2.719573e-07, 2.716158e-07, 2.720134e-07, 
    2.720801e-07, 2.719057e-07, 2.729169e-07, 2.726282e-07, 2.729237e-07, 
    2.727357e-07, 2.679899e-07, 2.682261e-07, 2.680985e-07, 2.683385e-07, 
    2.681694e-07, 2.689209e-07, 2.69146e-07, 2.701982e-07, 2.697665e-07, 
    2.704533e-07, 2.698363e-07, 2.699457e-07, 2.704758e-07, 2.698696e-07, 
    2.711942e-07, 2.702966e-07, 2.719627e-07, 2.710677e-07, 2.720187e-07, 
    2.718461e-07, 2.721319e-07, 2.723877e-07, 2.727094e-07, 2.733025e-07, 
    2.731652e-07, 2.736608e-07, 2.685781e-07, 2.688842e-07, 2.688573e-07, 
    2.691774e-07, 2.694141e-07, 2.699267e-07, 2.70748e-07, 2.704393e-07, 
    2.710059e-07, 2.711195e-07, 2.702587e-07, 2.707875e-07, 2.69089e-07, 
    2.693638e-07, 2.692002e-07, 2.686023e-07, 2.705105e-07, 2.69532e-07, 
    2.713375e-07, 2.708084e-07, 2.723513e-07, 2.715845e-07, 2.730896e-07, 
    2.737319e-07, 2.743355e-07, 2.750403e-07, 2.690512e-07, 2.688433e-07, 
    2.692155e-07, 2.697302e-07, 2.702071e-07, 2.708407e-07, 2.709055e-07, 
    2.710241e-07, 2.713311e-07, 2.715892e-07, 2.710617e-07, 2.716539e-07, 
    2.694276e-07, 2.705954e-07, 2.687647e-07, 2.693166e-07, 2.696998e-07, 
    2.695317e-07, 2.70404e-07, 2.706094e-07, 2.714434e-07, 2.710124e-07, 
    2.735735e-07, 2.724418e-07, 2.755762e-07, 2.747021e-07, 2.687706e-07, 
    2.690505e-07, 2.700234e-07, 2.695607e-07, 2.70883e-07, 2.712079e-07, 
    2.71472e-07, 2.718094e-07, 2.718458e-07, 2.720456e-07, 2.717182e-07, 
    2.720327e-07, 2.708421e-07, 2.713744e-07, 2.699122e-07, 2.702685e-07, 
    2.701046e-07, 2.699248e-07, 2.704795e-07, 2.710699e-07, 2.710824e-07, 
    2.712717e-07, 2.718046e-07, 2.708883e-07, 2.737195e-07, 2.719728e-07, 
    2.693555e-07, 2.698939e-07, 2.699707e-07, 2.697622e-07, 2.711754e-07, 
    2.706638e-07, 2.720408e-07, 2.716689e-07, 2.72278e-07, 2.719754e-07, 
    2.719309e-07, 2.71542e-07, 2.712997e-07, 2.706873e-07, 2.701884e-07, 
    2.697925e-07, 2.698845e-07, 2.703194e-07, 2.71106e-07, 2.718492e-07, 
    2.716864e-07, 2.722318e-07, 2.707872e-07, 2.713934e-07, 2.711592e-07, 
    2.717697e-07, 2.704311e-07, 2.715714e-07, 2.701393e-07, 2.70265e-07, 
    2.706536e-07, 2.714345e-07, 2.71607e-07, 2.717914e-07, 2.716776e-07, 
    2.711259e-07, 2.710355e-07, 2.706442e-07, 2.705361e-07, 2.702376e-07, 
    2.699904e-07, 2.702163e-07, 2.704534e-07, 2.711261e-07, 2.717318e-07, 
    2.723914e-07, 2.725526e-07, 2.733223e-07, 2.726959e-07, 2.737292e-07, 
    2.72851e-07, 2.743703e-07, 2.716373e-07, 2.72825e-07, 2.706713e-07, 
    2.709037e-07, 2.713238e-07, 2.722863e-07, 2.717668e-07, 2.723742e-07, 
    2.71032e-07, 2.703344e-07, 2.701537e-07, 2.698166e-07, 2.701614e-07, 
    2.701334e-07, 2.704632e-07, 2.703572e-07, 2.711485e-07, 2.707236e-07, 
    2.719298e-07, 2.723694e-07, 2.736089e-07, 2.743674e-07, 2.751383e-07, 
    2.754784e-07, 2.755818e-07, 2.75625e-07,
  2.415711e-07, 2.424821e-07, 2.423051e-07, 2.430394e-07, 2.426322e-07, 
    2.431129e-07, 2.417559e-07, 2.425183e-07, 2.420317e-07, 2.416532e-07, 
    2.444628e-07, 2.430722e-07, 2.459051e-07, 2.450199e-07, 2.47242e-07, 
    2.457674e-07, 2.47539e-07, 2.471995e-07, 2.482211e-07, 2.479285e-07, 
    2.492338e-07, 2.48356e-07, 2.499097e-07, 2.490243e-07, 2.491628e-07, 
    2.48327e-07, 2.433522e-07, 2.442897e-07, 2.432966e-07, 2.434304e-07, 
    2.433704e-07, 2.426406e-07, 2.422726e-07, 2.415014e-07, 2.416415e-07, 
    2.422078e-07, 2.434905e-07, 2.430553e-07, 2.441518e-07, 2.441271e-07, 
    2.453462e-07, 2.447967e-07, 2.468434e-07, 2.462622e-07, 2.479407e-07, 
    2.475189e-07, 2.479209e-07, 2.47799e-07, 2.479225e-07, 2.473037e-07, 
    2.475689e-07, 2.470242e-07, 2.448997e-07, 2.455246e-07, 2.436595e-07, 
    2.425361e-07, 2.417893e-07, 2.41259e-07, 2.41334e-07, 2.414769e-07, 
    2.422111e-07, 2.42901e-07, 2.434263e-07, 2.437775e-07, 2.441235e-07, 
    2.451698e-07, 2.457232e-07, 2.469609e-07, 2.467376e-07, 2.471158e-07, 
    2.474769e-07, 2.480828e-07, 2.479831e-07, 2.4825e-07, 2.471058e-07, 
    2.478664e-07, 2.466105e-07, 2.469541e-07, 2.442174e-07, 2.431728e-07, 
    2.427283e-07, 2.423391e-07, 2.413916e-07, 2.420461e-07, 2.417881e-07, 
    2.424017e-07, 2.427913e-07, 2.425986e-07, 2.437872e-07, 2.433252e-07, 
    2.457559e-07, 2.447098e-07, 2.474348e-07, 2.467835e-07, 2.475908e-07, 
    2.471789e-07, 2.478846e-07, 2.472495e-07, 2.483493e-07, 2.485886e-07, 
    2.484251e-07, 2.49053e-07, 2.472143e-07, 2.479209e-07, 2.425932e-07, 
    2.426246e-07, 2.42771e-07, 2.421273e-07, 2.420879e-07, 2.414976e-07, 
    2.420229e-07, 2.422465e-07, 2.428139e-07, 2.431493e-07, 2.434681e-07, 
    2.441685e-07, 2.449502e-07, 2.460421e-07, 2.468257e-07, 2.473506e-07, 
    2.470288e-07, 2.473129e-07, 2.469953e-07, 2.468464e-07, 2.484989e-07, 
    2.475714e-07, 2.489627e-07, 2.488858e-07, 2.482563e-07, 2.488945e-07, 
    2.426467e-07, 2.424658e-07, 2.418376e-07, 2.423293e-07, 2.414333e-07, 
    2.419349e-07, 2.422232e-07, 2.433349e-07, 2.43579e-07, 2.438052e-07, 
    2.442519e-07, 2.448249e-07, 2.458291e-07, 2.467019e-07, 2.474979e-07, 
    2.474396e-07, 2.474601e-07, 2.476379e-07, 2.471975e-07, 2.477101e-07, 
    2.477961e-07, 2.475713e-07, 2.488755e-07, 2.485031e-07, 2.488842e-07, 
    2.486417e-07, 2.425246e-07, 2.428289e-07, 2.426645e-07, 2.429736e-07, 
    2.427558e-07, 2.437239e-07, 2.440139e-07, 2.453698e-07, 2.448136e-07, 
    2.456986e-07, 2.449035e-07, 2.450444e-07, 2.457274e-07, 2.449465e-07, 
    2.466537e-07, 2.454966e-07, 2.476448e-07, 2.464905e-07, 2.477171e-07, 
    2.474945e-07, 2.47863e-07, 2.481929e-07, 2.486078e-07, 2.493727e-07, 
    2.491957e-07, 2.49835e-07, 2.432824e-07, 2.436767e-07, 2.43642e-07, 
    2.440545e-07, 2.443595e-07, 2.450201e-07, 2.460786e-07, 2.456807e-07, 
    2.464111e-07, 2.465576e-07, 2.45448e-07, 2.461294e-07, 2.439405e-07, 
    2.442945e-07, 2.440838e-07, 2.433135e-07, 2.457724e-07, 2.445113e-07, 
    2.468386e-07, 2.461565e-07, 2.481459e-07, 2.47157e-07, 2.490982e-07, 
    2.499266e-07, 2.507056e-07, 2.51615e-07, 2.438919e-07, 2.43624e-07, 
    2.441035e-07, 2.447666e-07, 2.453814e-07, 2.461981e-07, 2.462817e-07, 
    2.464346e-07, 2.468305e-07, 2.471633e-07, 2.464829e-07, 2.472466e-07, 
    2.443765e-07, 2.458818e-07, 2.435227e-07, 2.442337e-07, 2.447275e-07, 
    2.44511e-07, 2.456352e-07, 2.459e-07, 2.469751e-07, 2.464195e-07, 
    2.497222e-07, 2.482625e-07, 2.523068e-07, 2.511786e-07, 2.435304e-07, 
    2.438909e-07, 2.451446e-07, 2.445483e-07, 2.462527e-07, 2.466716e-07, 
    2.470121e-07, 2.474471e-07, 2.474941e-07, 2.477518e-07, 2.473295e-07, 
    2.477351e-07, 2.461999e-07, 2.468862e-07, 2.450014e-07, 2.454605e-07, 
    2.452494e-07, 2.450177e-07, 2.457326e-07, 2.464936e-07, 2.465098e-07, 
    2.467537e-07, 2.474405e-07, 2.462595e-07, 2.499104e-07, 2.476574e-07, 
    2.442839e-07, 2.449777e-07, 2.450768e-07, 2.448081e-07, 2.466296e-07, 
    2.459701e-07, 2.477455e-07, 2.47266e-07, 2.480515e-07, 2.476612e-07, 
    2.476038e-07, 2.471023e-07, 2.467899e-07, 2.460003e-07, 2.453573e-07, 
    2.448471e-07, 2.449657e-07, 2.455261e-07, 2.465401e-07, 2.474983e-07, 
    2.472885e-07, 2.479918e-07, 2.461292e-07, 2.469106e-07, 2.466087e-07, 
    2.473959e-07, 2.456702e-07, 2.471398e-07, 2.452941e-07, 2.454561e-07, 
    2.45957e-07, 2.469636e-07, 2.471862e-07, 2.474238e-07, 2.472772e-07, 
    2.465658e-07, 2.464493e-07, 2.459448e-07, 2.458054e-07, 2.454208e-07, 
    2.451022e-07, 2.453933e-07, 2.456989e-07, 2.465661e-07, 2.47347e-07, 
    2.481976e-07, 2.484056e-07, 2.493981e-07, 2.485902e-07, 2.499229e-07, 
    2.487899e-07, 2.507502e-07, 2.47225e-07, 2.487567e-07, 2.459797e-07, 
    2.462793e-07, 2.468209e-07, 2.480619e-07, 2.473922e-07, 2.481754e-07, 
    2.464447e-07, 2.455454e-07, 2.453126e-07, 2.448781e-07, 2.453226e-07, 
    2.452864e-07, 2.457115e-07, 2.45575e-07, 2.465949e-07, 2.460472e-07, 
    2.476024e-07, 2.481692e-07, 2.49768e-07, 2.507466e-07, 2.517417e-07, 
    2.521806e-07, 2.523142e-07, 2.5237e-07,
  2.260099e-07, 2.270073e-07, 2.268135e-07, 2.276176e-07, 2.271716e-07, 
    2.27698e-07, 2.262122e-07, 2.270469e-07, 2.265141e-07, 2.260998e-07, 
    2.291768e-07, 2.276535e-07, 2.307575e-07, 2.297872e-07, 2.322235e-07, 
    2.306066e-07, 2.325493e-07, 2.321769e-07, 2.332975e-07, 2.329765e-07, 
    2.344088e-07, 2.334456e-07, 2.351508e-07, 2.341789e-07, 2.343309e-07, 
    2.334138e-07, 2.279602e-07, 2.289872e-07, 2.278993e-07, 2.280458e-07, 
    2.279801e-07, 2.271808e-07, 2.267779e-07, 2.259337e-07, 2.26087e-07, 
    2.26707e-07, 2.281117e-07, 2.27635e-07, 2.288361e-07, 2.28809e-07, 
    2.301449e-07, 2.295427e-07, 2.317863e-07, 2.31149e-07, 2.329899e-07, 
    2.325272e-07, 2.329682e-07, 2.328345e-07, 2.3297e-07, 2.322912e-07, 
    2.325821e-07, 2.319847e-07, 2.296555e-07, 2.303404e-07, 2.282967e-07, 
    2.270665e-07, 2.262488e-07, 2.256683e-07, 2.257504e-07, 2.259069e-07, 
    2.267106e-07, 2.27466e-07, 2.280413e-07, 2.284261e-07, 2.288051e-07, 
    2.299516e-07, 2.305581e-07, 2.319152e-07, 2.316704e-07, 2.320851e-07, 
    2.324812e-07, 2.331459e-07, 2.330365e-07, 2.333292e-07, 2.320741e-07, 
    2.329084e-07, 2.315309e-07, 2.319078e-07, 2.28908e-07, 2.277636e-07, 
    2.272769e-07, 2.268508e-07, 2.258135e-07, 2.265299e-07, 2.262475e-07, 
    2.269192e-07, 2.273459e-07, 2.271349e-07, 2.284366e-07, 2.279306e-07, 
    2.30594e-07, 2.294474e-07, 2.32435e-07, 2.317206e-07, 2.326061e-07, 
    2.321543e-07, 2.329283e-07, 2.322318e-07, 2.334382e-07, 2.337008e-07, 
    2.335213e-07, 2.342104e-07, 2.321931e-07, 2.329682e-07, 2.27129e-07, 
    2.271634e-07, 2.273237e-07, 2.266188e-07, 2.265757e-07, 2.259295e-07, 
    2.265045e-07, 2.267493e-07, 2.273706e-07, 2.277379e-07, 2.280871e-07, 
    2.288544e-07, 2.297109e-07, 2.309077e-07, 2.317669e-07, 2.323426e-07, 
    2.319896e-07, 2.323013e-07, 2.319529e-07, 2.317896e-07, 2.336024e-07, 
    2.325848e-07, 2.341114e-07, 2.340269e-07, 2.333362e-07, 2.340364e-07, 
    2.271875e-07, 2.269895e-07, 2.263017e-07, 2.2684e-07, 2.258591e-07, 
    2.264082e-07, 2.267239e-07, 2.279412e-07, 2.282085e-07, 2.284564e-07, 
    2.289458e-07, 2.295735e-07, 2.306742e-07, 2.316311e-07, 2.325042e-07, 
    2.324402e-07, 2.324628e-07, 2.326577e-07, 2.321747e-07, 2.32737e-07, 
    2.328313e-07, 2.325847e-07, 2.340156e-07, 2.33607e-07, 2.340251e-07, 
    2.337591e-07, 2.270539e-07, 2.273871e-07, 2.27207e-07, 2.275456e-07, 
    2.273071e-07, 2.283673e-07, 2.28685e-07, 2.301707e-07, 2.295612e-07, 
    2.305312e-07, 2.296598e-07, 2.298142e-07, 2.305628e-07, 2.297069e-07, 
    2.315784e-07, 2.303098e-07, 2.326653e-07, 2.313994e-07, 2.327446e-07, 
    2.325004e-07, 2.329047e-07, 2.332666e-07, 2.337218e-07, 2.345613e-07, 
    2.34367e-07, 2.350688e-07, 2.278837e-07, 2.283156e-07, 2.282776e-07, 
    2.287295e-07, 2.290636e-07, 2.297875e-07, 2.309478e-07, 2.305116e-07, 
    2.313123e-07, 2.31473e-07, 2.302565e-07, 2.310035e-07, 2.286046e-07, 
    2.289924e-07, 2.287615e-07, 2.279177e-07, 2.306121e-07, 2.2923e-07, 
    2.317811e-07, 2.310332e-07, 2.33215e-07, 2.321303e-07, 2.3426e-07, 
    2.351693e-07, 2.360247e-07, 2.370235e-07, 2.285513e-07, 2.282579e-07, 
    2.287832e-07, 2.295097e-07, 2.301835e-07, 2.310788e-07, 2.311704e-07, 
    2.31338e-07, 2.317722e-07, 2.321371e-07, 2.31391e-07, 2.322286e-07, 
    2.290823e-07, 2.30732e-07, 2.281469e-07, 2.289258e-07, 2.294669e-07, 
    2.292296e-07, 2.304617e-07, 2.30752e-07, 2.319308e-07, 2.313216e-07, 
    2.349449e-07, 2.33343e-07, 2.377836e-07, 2.365441e-07, 2.281553e-07, 
    2.285503e-07, 2.29924e-07, 2.292706e-07, 2.311386e-07, 2.31598e-07, 
    2.319714e-07, 2.324485e-07, 2.325e-07, 2.327826e-07, 2.323195e-07, 
    2.327644e-07, 2.310807e-07, 2.318333e-07, 2.297671e-07, 2.302702e-07, 
    2.300388e-07, 2.297849e-07, 2.305684e-07, 2.314028e-07, 2.314206e-07, 
    2.31688e-07, 2.324412e-07, 2.311461e-07, 2.351515e-07, 2.326792e-07, 
    2.289808e-07, 2.29741e-07, 2.298496e-07, 2.295552e-07, 2.315519e-07, 
    2.308288e-07, 2.327757e-07, 2.322498e-07, 2.331115e-07, 2.326833e-07, 
    2.326204e-07, 2.320703e-07, 2.317277e-07, 2.308619e-07, 2.301571e-07, 
    2.295979e-07, 2.297279e-07, 2.303421e-07, 2.314538e-07, 2.325047e-07, 
    2.322745e-07, 2.33046e-07, 2.310032e-07, 2.318601e-07, 2.31529e-07, 
    2.323923e-07, 2.305e-07, 2.321114e-07, 2.300878e-07, 2.302653e-07, 
    2.308144e-07, 2.319182e-07, 2.321623e-07, 2.324229e-07, 2.322621e-07, 
    2.31482e-07, 2.313542e-07, 2.308011e-07, 2.306483e-07, 2.302267e-07, 
    2.298775e-07, 2.301965e-07, 2.305315e-07, 2.314823e-07, 2.323387e-07, 
    2.332717e-07, 2.335e-07, 2.345892e-07, 2.337026e-07, 2.351652e-07, 
    2.339217e-07, 2.360737e-07, 2.322048e-07, 2.338852e-07, 2.308394e-07, 
    2.311678e-07, 2.317617e-07, 2.331229e-07, 2.323882e-07, 2.332474e-07, 
    2.313492e-07, 2.303633e-07, 2.301081e-07, 2.296319e-07, 2.30119e-07, 
    2.300794e-07, 2.305454e-07, 2.303956e-07, 2.315139e-07, 2.309133e-07, 
    2.326188e-07, 2.332406e-07, 2.349952e-07, 2.360698e-07, 2.371627e-07, 
    2.376449e-07, 2.377917e-07, 2.37853e-07,
  2.166787e-07, 2.177053e-07, 2.175057e-07, 2.183336e-07, 2.178744e-07, 
    2.184165e-07, 2.168868e-07, 2.17746e-07, 2.171975e-07, 2.167711e-07, 
    2.1994e-07, 2.183705e-07, 2.215696e-07, 2.205691e-07, 2.230822e-07, 
    2.21414e-07, 2.234185e-07, 2.23034e-07, 2.24191e-07, 2.238595e-07, 
    2.253391e-07, 2.243439e-07, 2.261059e-07, 2.251014e-07, 2.252586e-07, 
    2.243111e-07, 2.186864e-07, 2.197446e-07, 2.186237e-07, 2.187746e-07, 
    2.187069e-07, 2.178839e-07, 2.174691e-07, 2.166002e-07, 2.167579e-07, 
    2.173961e-07, 2.188425e-07, 2.183515e-07, 2.195887e-07, 2.195608e-07, 
    2.209378e-07, 2.20317e-07, 2.22631e-07, 2.219734e-07, 2.238734e-07, 
    2.233956e-07, 2.238509e-07, 2.237129e-07, 2.238527e-07, 2.23152e-07, 
    2.234523e-07, 2.228356e-07, 2.204333e-07, 2.211394e-07, 2.190331e-07, 
    2.177662e-07, 2.169245e-07, 2.163272e-07, 2.164116e-07, 2.165726e-07, 
    2.173998e-07, 2.181774e-07, 2.1877e-07, 2.191663e-07, 2.195568e-07, 
    2.207386e-07, 2.213639e-07, 2.227639e-07, 2.225113e-07, 2.229393e-07, 
    2.233481e-07, 2.240344e-07, 2.239214e-07, 2.242238e-07, 2.22928e-07, 
    2.237892e-07, 2.223674e-07, 2.227563e-07, 2.19663e-07, 2.18484e-07, 
    2.179828e-07, 2.175441e-07, 2.164766e-07, 2.172138e-07, 2.169232e-07, 
    2.176145e-07, 2.180538e-07, 2.178365e-07, 2.191771e-07, 2.18656e-07, 
    2.21401e-07, 2.202188e-07, 2.233004e-07, 2.225632e-07, 2.234771e-07, 
    2.230108e-07, 2.238098e-07, 2.230907e-07, 2.243363e-07, 2.246075e-07, 
    2.244222e-07, 2.25134e-07, 2.230508e-07, 2.238509e-07, 2.178304e-07, 
    2.178659e-07, 2.180309e-07, 2.173053e-07, 2.172609e-07, 2.165959e-07, 
    2.171876e-07, 2.174396e-07, 2.180792e-07, 2.184575e-07, 2.188171e-07, 
    2.196076e-07, 2.204904e-07, 2.217245e-07, 2.22611e-07, 2.232051e-07, 
    2.228408e-07, 2.231624e-07, 2.228029e-07, 2.226343e-07, 2.245059e-07, 
    2.234551e-07, 2.250316e-07, 2.249444e-07, 2.24231e-07, 2.249542e-07, 
    2.178907e-07, 2.176868e-07, 2.169789e-07, 2.175329e-07, 2.165234e-07, 
    2.170885e-07, 2.174134e-07, 2.186669e-07, 2.189422e-07, 2.191975e-07, 
    2.197018e-07, 2.203488e-07, 2.214836e-07, 2.224708e-07, 2.233719e-07, 
    2.233059e-07, 2.233291e-07, 2.235304e-07, 2.230318e-07, 2.236122e-07, 
    2.237096e-07, 2.234549e-07, 2.249327e-07, 2.245106e-07, 2.249426e-07, 
    2.246677e-07, 2.177531e-07, 2.180962e-07, 2.179108e-07, 2.182594e-07, 
    2.180138e-07, 2.191058e-07, 2.194331e-07, 2.209645e-07, 2.20336e-07, 
    2.213362e-07, 2.204376e-07, 2.205969e-07, 2.213688e-07, 2.204862e-07, 
    2.224164e-07, 2.211079e-07, 2.235382e-07, 2.222318e-07, 2.2362e-07, 
    2.23368e-07, 2.237853e-07, 2.241591e-07, 2.246292e-07, 2.254966e-07, 
    2.252958e-07, 2.260211e-07, 2.186076e-07, 2.190525e-07, 2.190133e-07, 
    2.194789e-07, 2.198232e-07, 2.205693e-07, 2.217658e-07, 2.213159e-07, 
    2.221418e-07, 2.223076e-07, 2.210528e-07, 2.218233e-07, 2.193503e-07, 
    2.197499e-07, 2.195119e-07, 2.186427e-07, 2.214196e-07, 2.199947e-07, 
    2.226256e-07, 2.218539e-07, 2.241058e-07, 2.22986e-07, 2.251852e-07, 
    2.261251e-07, 2.270095e-07, 2.280428e-07, 2.192953e-07, 2.18993e-07, 
    2.195343e-07, 2.20283e-07, 2.209776e-07, 2.21901e-07, 2.219954e-07, 
    2.221684e-07, 2.226164e-07, 2.22993e-07, 2.222231e-07, 2.230874e-07, 
    2.198426e-07, 2.215433e-07, 2.188787e-07, 2.196812e-07, 2.202389e-07, 
    2.199943e-07, 2.212645e-07, 2.215638e-07, 2.227801e-07, 2.221514e-07, 
    2.258932e-07, 2.24238e-07, 2.288294e-07, 2.275468e-07, 2.188874e-07, 
    2.192943e-07, 2.207101e-07, 2.200365e-07, 2.219626e-07, 2.224366e-07, 
    2.228219e-07, 2.233144e-07, 2.233676e-07, 2.236593e-07, 2.231812e-07, 
    2.236405e-07, 2.219029e-07, 2.226795e-07, 2.205483e-07, 2.210671e-07, 
    2.208284e-07, 2.205666e-07, 2.213745e-07, 2.222352e-07, 2.222536e-07, 
    2.225295e-07, 2.233071e-07, 2.219704e-07, 2.261068e-07, 2.235527e-07, 
    2.197379e-07, 2.205215e-07, 2.206334e-07, 2.203298e-07, 2.223891e-07, 
    2.21643e-07, 2.236522e-07, 2.231093e-07, 2.239989e-07, 2.235568e-07, 
    2.234918e-07, 2.22924e-07, 2.225705e-07, 2.216773e-07, 2.209504e-07, 
    2.203739e-07, 2.205079e-07, 2.211412e-07, 2.222878e-07, 2.233724e-07, 
    2.231348e-07, 2.239313e-07, 2.21823e-07, 2.227071e-07, 2.223654e-07, 
    2.232564e-07, 2.21304e-07, 2.229666e-07, 2.208789e-07, 2.21062e-07, 
    2.216282e-07, 2.227671e-07, 2.23019e-07, 2.23288e-07, 2.23122e-07, 
    2.223169e-07, 2.22185e-07, 2.216145e-07, 2.214569e-07, 2.210221e-07, 
    2.206621e-07, 2.20991e-07, 2.213364e-07, 2.223173e-07, 2.23201e-07, 
    2.241644e-07, 2.244001e-07, 2.255255e-07, 2.246094e-07, 2.26121e-07, 
    2.248359e-07, 2.270602e-07, 2.230629e-07, 2.247981e-07, 2.21654e-07, 
    2.219928e-07, 2.226056e-07, 2.240107e-07, 2.232522e-07, 2.241393e-07, 
    2.221799e-07, 2.21163e-07, 2.208999e-07, 2.204089e-07, 2.209111e-07, 
    2.208702e-07, 2.213507e-07, 2.211963e-07, 2.223498e-07, 2.217303e-07, 
    2.234902e-07, 2.241323e-07, 2.259451e-07, 2.270561e-07, 2.281868e-07, 
    2.286858e-07, 2.288377e-07, 2.289012e-07,
  2.081591e-07, 2.091279e-07, 2.089395e-07, 2.097213e-07, 2.092875e-07, 
    2.097996e-07, 2.083554e-07, 2.091664e-07, 2.086486e-07, 2.082462e-07, 
    2.112399e-07, 2.097562e-07, 2.127824e-07, 2.11835e-07, 2.142161e-07, 
    2.12635e-07, 2.145351e-07, 2.141704e-07, 2.152682e-07, 2.149536e-07, 
    2.163589e-07, 2.154134e-07, 2.170879e-07, 2.16133e-07, 2.162824e-07, 
    2.153823e-07, 2.100546e-07, 2.110551e-07, 2.099953e-07, 2.10138e-07, 
    2.10074e-07, 2.092965e-07, 2.08905e-07, 2.08085e-07, 2.082338e-07, 
    2.08836e-07, 2.102021e-07, 2.097382e-07, 2.109075e-07, 2.108811e-07, 
    2.12184e-07, 2.115964e-07, 2.137882e-07, 2.131649e-07, 2.149667e-07, 
    2.145134e-07, 2.149454e-07, 2.148144e-07, 2.149471e-07, 2.142823e-07, 
    2.145671e-07, 2.139822e-07, 2.117065e-07, 2.123749e-07, 2.103822e-07, 
    2.091855e-07, 2.08391e-07, 2.078275e-07, 2.079071e-07, 2.08059e-07, 
    2.088396e-07, 2.095738e-07, 2.101335e-07, 2.105081e-07, 2.108773e-07, 
    2.119955e-07, 2.125876e-07, 2.139143e-07, 2.136747e-07, 2.140805e-07, 
    2.144683e-07, 2.151196e-07, 2.150123e-07, 2.152994e-07, 2.140698e-07, 
    2.148869e-07, 2.135382e-07, 2.13907e-07, 2.109779e-07, 2.098633e-07, 
    2.0939e-07, 2.089757e-07, 2.079684e-07, 2.08664e-07, 2.083897e-07, 
    2.090422e-07, 2.09457e-07, 2.092518e-07, 2.105184e-07, 2.100258e-07, 
    2.126227e-07, 2.115035e-07, 2.14423e-07, 2.137239e-07, 2.145907e-07, 
    2.141483e-07, 2.149064e-07, 2.142241e-07, 2.154062e-07, 2.156638e-07, 
    2.154878e-07, 2.16164e-07, 2.141863e-07, 2.149455e-07, 2.092461e-07, 
    2.092795e-07, 2.094354e-07, 2.087504e-07, 2.087085e-07, 2.080809e-07, 
    2.086393e-07, 2.088771e-07, 2.09481e-07, 2.098383e-07, 2.101781e-07, 
    2.109254e-07, 2.117605e-07, 2.129291e-07, 2.137692e-07, 2.143326e-07, 
    2.139871e-07, 2.142921e-07, 2.139511e-07, 2.137913e-07, 2.155673e-07, 
    2.145698e-07, 2.160667e-07, 2.159838e-07, 2.153062e-07, 2.159931e-07, 
    2.09303e-07, 2.091105e-07, 2.084423e-07, 2.089652e-07, 2.080126e-07, 
    2.085458e-07, 2.088524e-07, 2.100362e-07, 2.102963e-07, 2.105377e-07, 
    2.110144e-07, 2.116265e-07, 2.127009e-07, 2.136363e-07, 2.144908e-07, 
    2.144282e-07, 2.144502e-07, 2.146412e-07, 2.141682e-07, 2.147189e-07, 
    2.148113e-07, 2.145696e-07, 2.159727e-07, 2.155717e-07, 2.15982e-07, 
    2.157209e-07, 2.091731e-07, 2.09497e-07, 2.09322e-07, 2.096512e-07, 
    2.094193e-07, 2.10451e-07, 2.107604e-07, 2.122093e-07, 2.116145e-07, 
    2.125613e-07, 2.117106e-07, 2.118613e-07, 2.125923e-07, 2.117565e-07, 
    2.135848e-07, 2.123451e-07, 2.146486e-07, 2.134098e-07, 2.147263e-07, 
    2.144871e-07, 2.148831e-07, 2.152379e-07, 2.156844e-07, 2.165086e-07, 
    2.163177e-07, 2.170073e-07, 2.099801e-07, 2.104006e-07, 2.103636e-07, 
    2.108037e-07, 2.111293e-07, 2.118352e-07, 2.129682e-07, 2.12542e-07, 
    2.133245e-07, 2.134816e-07, 2.122929e-07, 2.130227e-07, 2.106821e-07, 
    2.1106e-07, 2.108349e-07, 2.100133e-07, 2.126403e-07, 2.112915e-07, 
    2.137831e-07, 2.130516e-07, 2.151874e-07, 2.141249e-07, 2.162126e-07, 
    2.171063e-07, 2.179476e-07, 2.189318e-07, 2.106301e-07, 2.103443e-07, 
    2.10856e-07, 2.115643e-07, 2.122217e-07, 2.130962e-07, 2.131857e-07, 
    2.133497e-07, 2.137743e-07, 2.141314e-07, 2.134015e-07, 2.14221e-07, 
    2.111478e-07, 2.127574e-07, 2.102364e-07, 2.109951e-07, 2.115225e-07, 
    2.112911e-07, 2.124933e-07, 2.127768e-07, 2.139295e-07, 2.133335e-07, 
    2.168857e-07, 2.15313e-07, 2.196815e-07, 2.184593e-07, 2.102445e-07, 
    2.106291e-07, 2.119685e-07, 2.11331e-07, 2.131546e-07, 2.136039e-07, 
    2.139692e-07, 2.144363e-07, 2.144867e-07, 2.147636e-07, 2.143099e-07, 
    2.147457e-07, 2.130981e-07, 2.138341e-07, 2.118152e-07, 2.123064e-07, 
    2.120804e-07, 2.118326e-07, 2.125975e-07, 2.13413e-07, 2.134304e-07, 
    2.13692e-07, 2.144296e-07, 2.13162e-07, 2.17089e-07, 2.146626e-07, 
    2.110486e-07, 2.1179e-07, 2.118958e-07, 2.116086e-07, 2.135588e-07, 
    2.128519e-07, 2.147569e-07, 2.142417e-07, 2.150858e-07, 2.146663e-07, 
    2.146046e-07, 2.14066e-07, 2.137308e-07, 2.128843e-07, 2.121959e-07, 
    2.116502e-07, 2.117771e-07, 2.123766e-07, 2.134629e-07, 2.144913e-07, 
    2.14266e-07, 2.150217e-07, 2.130223e-07, 2.138604e-07, 2.135364e-07, 
    2.143812e-07, 2.125307e-07, 2.141066e-07, 2.121282e-07, 2.123015e-07, 
    2.128378e-07, 2.139173e-07, 2.141561e-07, 2.144113e-07, 2.142538e-07, 
    2.134905e-07, 2.133654e-07, 2.128248e-07, 2.126756e-07, 2.122638e-07, 
    2.11923e-07, 2.122344e-07, 2.125615e-07, 2.134908e-07, 2.143288e-07, 
    2.15243e-07, 2.154668e-07, 2.165361e-07, 2.156657e-07, 2.171025e-07, 
    2.15881e-07, 2.179961e-07, 2.141979e-07, 2.158449e-07, 2.128622e-07, 
    2.131832e-07, 2.137641e-07, 2.150972e-07, 2.143773e-07, 2.152192e-07, 
    2.133605e-07, 2.123973e-07, 2.121481e-07, 2.116834e-07, 2.121587e-07, 
    2.1212e-07, 2.12575e-07, 2.124288e-07, 2.135216e-07, 2.129345e-07, 
    2.146031e-07, 2.152125e-07, 2.16935e-07, 2.179921e-07, 2.190689e-07, 
    2.195446e-07, 2.196894e-07, 2.1975e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.359163e-08, 6.387121e-08, 6.381686e-08, 6.404235e-08, 6.391726e-08, 
    6.406492e-08, 6.364831e-08, 6.388231e-08, 6.373293e-08, 6.36168e-08, 
    6.447997e-08, 6.405241e-08, 6.492405e-08, 6.465138e-08, 6.533632e-08, 
    6.488163e-08, 6.542801e-08, 6.53232e-08, 6.563863e-08, 6.554826e-08, 
    6.595173e-08, 6.568033e-08, 6.616087e-08, 6.588692e-08, 6.592978e-08, 
    6.567138e-08, 6.413845e-08, 6.442674e-08, 6.412137e-08, 6.416248e-08, 
    6.414403e-08, 6.391985e-08, 6.380688e-08, 6.357025e-08, 6.361321e-08, 
    6.3787e-08, 6.418097e-08, 6.404723e-08, 6.438426e-08, 6.437665e-08, 
    6.475187e-08, 6.458269e-08, 6.521333e-08, 6.503409e-08, 6.555204e-08, 
    6.542178e-08, 6.554592e-08, 6.550827e-08, 6.554641e-08, 6.535537e-08, 
    6.543722e-08, 6.526912e-08, 6.461438e-08, 6.480681e-08, 6.423289e-08, 
    6.38878e-08, 6.365858e-08, 6.349591e-08, 6.351891e-08, 6.356274e-08, 
    6.378801e-08, 6.399981e-08, 6.416121e-08, 6.426918e-08, 6.437556e-08, 
    6.469757e-08, 6.486799e-08, 6.524958e-08, 6.518071e-08, 6.529738e-08, 
    6.540882e-08, 6.559594e-08, 6.556514e-08, 6.564758e-08, 6.529429e-08, 
    6.552909e-08, 6.514148e-08, 6.52475e-08, 6.44045e-08, 6.40833e-08, 
    6.394681e-08, 6.38273e-08, 6.353659e-08, 6.373735e-08, 6.365821e-08, 
    6.384649e-08, 6.396612e-08, 6.390695e-08, 6.427213e-08, 6.413016e-08, 
    6.487809e-08, 6.455593e-08, 6.539582e-08, 6.519484e-08, 6.544399e-08, 
    6.531685e-08, 6.55347e-08, 6.533864e-08, 6.567826e-08, 6.575221e-08, 
    6.570168e-08, 6.58958e-08, 6.532778e-08, 6.554592e-08, 6.39053e-08, 
    6.391495e-08, 6.39599e-08, 6.376228e-08, 6.375019e-08, 6.356908e-08, 
    6.373023e-08, 6.379886e-08, 6.397305e-08, 6.40761e-08, 6.417405e-08, 
    6.438941e-08, 6.462994e-08, 6.496626e-08, 6.520787e-08, 6.536983e-08, 
    6.527052e-08, 6.53582e-08, 6.526018e-08, 6.521424e-08, 6.572451e-08, 
    6.543799e-08, 6.586788e-08, 6.584409e-08, 6.564954e-08, 6.584677e-08, 
    6.392172e-08, 6.386619e-08, 6.367338e-08, 6.382427e-08, 6.354936e-08, 
    6.370324e-08, 6.379173e-08, 6.413313e-08, 6.420814e-08, 6.427769e-08, 
    6.441505e-08, 6.459135e-08, 6.49006e-08, 6.516968e-08, 6.54153e-08, 
    6.539731e-08, 6.540364e-08, 6.545852e-08, 6.53226e-08, 6.548083e-08, 
    6.550739e-08, 6.543795e-08, 6.58409e-08, 6.572579e-08, 6.584358e-08, 
    6.576862e-08, 6.388424e-08, 6.397768e-08, 6.392719e-08, 6.402214e-08, 
    6.395525e-08, 6.425269e-08, 6.434187e-08, 6.475913e-08, 6.458788e-08, 
    6.486043e-08, 6.461556e-08, 6.465896e-08, 6.486933e-08, 6.462879e-08, 
    6.515485e-08, 6.479821e-08, 6.546065e-08, 6.510453e-08, 6.548296e-08, 
    6.541424e-08, 6.552803e-08, 6.562993e-08, 6.575814e-08, 6.59947e-08, 
    6.593991e-08, 6.613774e-08, 6.411698e-08, 6.423819e-08, 6.422751e-08, 
    6.435434e-08, 6.444814e-08, 6.465145e-08, 6.497752e-08, 6.485489e-08, 
    6.508e-08, 6.512519e-08, 6.47832e-08, 6.499319e-08, 6.431929e-08, 
    6.442818e-08, 6.436335e-08, 6.412655e-08, 6.488316e-08, 6.449487e-08, 
    6.521186e-08, 6.500152e-08, 6.56154e-08, 6.531011e-08, 6.590976e-08, 
    6.616612e-08, 6.640736e-08, 6.668932e-08, 6.430432e-08, 6.422197e-08, 
    6.436942e-08, 6.457343e-08, 6.476271e-08, 6.501435e-08, 6.504009e-08, 
    6.508724e-08, 6.520934e-08, 6.531201e-08, 6.510215e-08, 6.533775e-08, 
    6.445345e-08, 6.491686e-08, 6.419084e-08, 6.440948e-08, 6.456141e-08, 
    6.449476e-08, 6.484088e-08, 6.492246e-08, 6.525397e-08, 6.50826e-08, 
    6.610285e-08, 6.565147e-08, 6.690398e-08, 6.655396e-08, 6.41932e-08, 
    6.430404e-08, 6.46898e-08, 6.450625e-08, 6.503114e-08, 6.516034e-08, 
    6.526538e-08, 6.539964e-08, 6.541413e-08, 6.549368e-08, 6.536332e-08, 
    6.548853e-08, 6.501489e-08, 6.522654e-08, 6.46457e-08, 6.478708e-08, 
    6.472204e-08, 6.46507e-08, 6.487087e-08, 6.510545e-08, 6.511046e-08, 
    6.518567e-08, 6.539766e-08, 6.503327e-08, 6.616113e-08, 6.546461e-08, 
    6.44249e-08, 6.463841e-08, 6.466889e-08, 6.458619e-08, 6.514739e-08, 
    6.494405e-08, 6.549174e-08, 6.534372e-08, 6.558625e-08, 6.546573e-08, 
    6.5448e-08, 6.529321e-08, 6.519684e-08, 6.495338e-08, 6.475528e-08, 
    6.459818e-08, 6.463471e-08, 6.480727e-08, 6.51198e-08, 6.541545e-08, 
    6.535068e-08, 6.556781e-08, 6.499309e-08, 6.523408e-08, 6.514095e-08, 
    6.538381e-08, 6.485164e-08, 6.530484e-08, 6.47358e-08, 6.47857e-08, 
    6.494002e-08, 6.525044e-08, 6.53191e-08, 6.539243e-08, 6.534718e-08, 
    6.512773e-08, 6.509178e-08, 6.493626e-08, 6.489333e-08, 6.477483e-08, 
    6.467673e-08, 6.476636e-08, 6.486049e-08, 6.512782e-08, 6.536873e-08, 
    6.563138e-08, 6.569566e-08, 6.600256e-08, 6.575274e-08, 6.616501e-08, 
    6.581453e-08, 6.642122e-08, 6.533109e-08, 6.58042e-08, 6.494704e-08, 
    6.503938e-08, 6.520641e-08, 6.558949e-08, 6.538266e-08, 6.562454e-08, 
    6.509037e-08, 6.481324e-08, 6.474151e-08, 6.460773e-08, 6.474458e-08, 
    6.473344e-08, 6.486439e-08, 6.482231e-08, 6.51367e-08, 6.496782e-08, 
    6.544756e-08, 6.562262e-08, 6.611701e-08, 6.642009e-08, 6.672858e-08, 
    6.686479e-08, 6.690624e-08, 6.692357e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10 ;

 LEAFN =
  0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09 ;

 LITHR =
  9.042218e-13, 9.066582e-13, 9.06185e-13, 9.081482e-13, 9.070596e-13, 
    9.083447e-13, 9.047163e-13, 9.067546e-13, 9.054538e-13, 9.044417e-13, 
    9.119526e-13, 9.082358e-13, 9.158099e-13, 9.134437e-13, 9.193833e-13, 
    9.154413e-13, 9.201776e-13, 9.192704e-13, 9.220014e-13, 9.212194e-13, 
    9.247071e-13, 9.223622e-13, 9.265142e-13, 9.241478e-13, 9.245178e-13, 
    9.222847e-13, 9.08985e-13, 9.1149e-13, 9.088363e-13, 9.091937e-13, 
    9.090335e-13, 9.070819e-13, 9.060972e-13, 9.04036e-13, 9.044105e-13, 
    9.059246e-13, 9.093545e-13, 9.081912e-13, 9.111232e-13, 9.11057e-13, 
    9.143163e-13, 9.128474e-13, 9.183185e-13, 9.167654e-13, 9.212521e-13, 
    9.201243e-13, 9.21199e-13, 9.208733e-13, 9.212032e-13, 9.195491e-13, 
    9.202579e-13, 9.18802e-13, 9.131223e-13, 9.14793e-13, 9.098064e-13, 
    9.068017e-13, 9.048056e-13, 9.033876e-13, 9.035881e-13, 9.039702e-13, 
    9.059335e-13, 9.077785e-13, 9.091833e-13, 9.101225e-13, 9.110475e-13, 
    9.138434e-13, 9.153234e-13, 9.186321e-13, 9.180359e-13, 9.190463e-13, 
    9.200121e-13, 9.216318e-13, 9.213653e-13, 9.220785e-13, 9.190202e-13, 
    9.210529e-13, 9.17696e-13, 9.186147e-13, 9.112964e-13, 9.085052e-13, 
    9.073157e-13, 9.062758e-13, 9.037423e-13, 9.05492e-13, 9.048023e-13, 
    9.064434e-13, 9.074851e-13, 9.0697e-13, 9.101482e-13, 9.08913e-13, 
    9.154111e-13, 9.126145e-13, 9.198995e-13, 9.181583e-13, 9.203168e-13, 
    9.192158e-13, 9.211016e-13, 9.194044e-13, 9.22344e-13, 9.229834e-13, 
    9.225464e-13, 9.242251e-13, 9.193102e-13, 9.211988e-13, 9.069555e-13, 
    9.070395e-13, 9.074311e-13, 9.057092e-13, 9.05604e-13, 9.040256e-13, 
    9.054304e-13, 9.060281e-13, 9.075457e-13, 9.084425e-13, 9.092948e-13, 
    9.111677e-13, 9.132571e-13, 9.161764e-13, 9.182712e-13, 9.196746e-13, 
    9.188143e-13, 9.195738e-13, 9.187247e-13, 9.183267e-13, 9.227437e-13, 
    9.202643e-13, 9.239838e-13, 9.237782e-13, 9.220953e-13, 9.238014e-13, 
    9.070985e-13, 9.06615e-13, 9.049348e-13, 9.062498e-13, 9.038537e-13, 
    9.051949e-13, 9.059656e-13, 9.089383e-13, 9.095915e-13, 9.101963e-13, 
    9.113908e-13, 9.129225e-13, 9.156069e-13, 9.1794e-13, 9.200684e-13, 
    9.199126e-13, 9.199674e-13, 9.204423e-13, 9.192653e-13, 9.206355e-13, 
    9.208652e-13, 9.202643e-13, 9.237507e-13, 9.227553e-13, 9.237739e-13, 
    9.231258e-13, 9.067723e-13, 9.075858e-13, 9.071462e-13, 9.079726e-13, 
    9.073903e-13, 9.099781e-13, 9.107536e-13, 9.143787e-13, 9.128923e-13, 
    9.152582e-13, 9.131329e-13, 9.135095e-13, 9.153342e-13, 9.13248e-13, 
    9.178109e-13, 9.147175e-13, 9.204609e-13, 9.173745e-13, 9.206541e-13, 
    9.200592e-13, 9.210443e-13, 9.219259e-13, 9.23035e-13, 9.250792e-13, 
    9.246061e-13, 9.26315e-13, 9.087983e-13, 9.098524e-13, 9.0976e-13, 
    9.10863e-13, 9.116782e-13, 9.134447e-13, 9.162744e-13, 9.152108e-13, 
    9.171635e-13, 9.175547e-13, 9.145887e-13, 9.164101e-13, 9.105579e-13, 
    9.115039e-13, 9.10941e-13, 9.088812e-13, 9.154553e-13, 9.120836e-13, 
    9.183058e-13, 9.164827e-13, 9.218002e-13, 9.191566e-13, 9.243456e-13, 
    9.265587e-13, 9.28642e-13, 9.310713e-13, 9.10428e-13, 9.097119e-13, 
    9.109943e-13, 9.127663e-13, 9.144105e-13, 9.165938e-13, 9.168174e-13, 
    9.17226e-13, 9.182842e-13, 9.191737e-13, 9.173547e-13, 9.193967e-13, 
    9.117223e-13, 9.157479e-13, 9.094407e-13, 9.113412e-13, 9.12662e-13, 
    9.120832e-13, 9.150894e-13, 9.157972e-13, 9.186703e-13, 9.17186e-13, 
    9.260123e-13, 9.221113e-13, 9.329207e-13, 9.299051e-13, 9.094616e-13, 
    9.104257e-13, 9.137772e-13, 9.121832e-13, 9.167398e-13, 9.178593e-13, 
    9.187697e-13, 9.199323e-13, 9.200581e-13, 9.207467e-13, 9.196182e-13, 
    9.207023e-13, 9.165985e-13, 9.184332e-13, 9.133949e-13, 9.14622e-13, 
    9.140578e-13, 9.134383e-13, 9.153496e-13, 9.173828e-13, 9.174271e-13, 
    9.180785e-13, 9.199124e-13, 9.167583e-13, 9.265139e-13, 9.204924e-13, 
    9.114765e-13, 9.133304e-13, 9.13596e-13, 9.12878e-13, 9.17747e-13, 
    9.159842e-13, 9.2073e-13, 9.194484e-13, 9.215481e-13, 9.205049e-13, 
    9.203514e-13, 9.190109e-13, 9.181757e-13, 9.16065e-13, 9.143459e-13, 
    9.129821e-13, 9.132994e-13, 9.147972e-13, 9.175073e-13, 9.200693e-13, 
    9.195082e-13, 9.213886e-13, 9.164097e-13, 9.184981e-13, 9.176907e-13, 
    9.197955e-13, 9.151824e-13, 9.19109e-13, 9.141773e-13, 9.146103e-13, 
    9.159492e-13, 9.186392e-13, 9.192352e-13, 9.1987e-13, 9.194785e-13, 
    9.175762e-13, 9.172653e-13, 9.159169e-13, 9.15544e-13, 9.145161e-13, 
    9.136643e-13, 9.144423e-13, 9.15259e-13, 9.175773e-13, 9.196646e-13, 
    9.219383e-13, 9.224947e-13, 9.251457e-13, 9.229868e-13, 9.265471e-13, 
    9.23519e-13, 9.287591e-13, 9.193374e-13, 9.234315e-13, 9.160103e-13, 
    9.168112e-13, 9.182579e-13, 9.21575e-13, 9.197856e-13, 9.218786e-13, 
    9.172531e-13, 9.148484e-13, 9.142268e-13, 9.13065e-13, 9.142534e-13, 
    9.141568e-13, 9.152933e-13, 9.149282e-13, 9.176543e-13, 9.161906e-13, 
    9.203472e-13, 9.218622e-13, 9.261357e-13, 9.287508e-13, 9.314109e-13, 
    9.325837e-13, 9.329406e-13, 9.330898e-13 ;

 LITR1C =
  3.186869e-05, 3.186857e-05, 3.186859e-05, 3.186849e-05, 3.186855e-05, 
    3.186848e-05, 3.186867e-05, 3.186856e-05, 3.186863e-05, 3.186868e-05, 
    3.186829e-05, 3.186848e-05, 3.186809e-05, 3.186821e-05, 3.186791e-05, 
    3.186811e-05, 3.186786e-05, 3.186791e-05, 3.186777e-05, 3.186781e-05, 
    3.186763e-05, 3.186775e-05, 3.186754e-05, 3.186766e-05, 3.186764e-05, 
    3.186776e-05, 3.186845e-05, 3.186832e-05, 3.186845e-05, 3.186844e-05, 
    3.186844e-05, 3.186855e-05, 3.18686e-05, 3.18687e-05, 3.186868e-05, 
    3.18686e-05, 3.186843e-05, 3.186849e-05, 3.186833e-05, 3.186834e-05, 
    3.186817e-05, 3.186825e-05, 3.186796e-05, 3.186804e-05, 3.186781e-05, 
    3.186787e-05, 3.186781e-05, 3.186783e-05, 3.186781e-05, 3.18679e-05, 
    3.186786e-05, 3.186794e-05, 3.186823e-05, 3.186815e-05, 3.18684e-05, 
    3.186856e-05, 3.186866e-05, 3.186873e-05, 3.186872e-05, 3.186871e-05, 
    3.18686e-05, 3.186851e-05, 3.186844e-05, 3.186839e-05, 3.186834e-05, 
    3.18682e-05, 3.186812e-05, 3.186794e-05, 3.186798e-05, 3.186793e-05, 
    3.186788e-05, 3.186779e-05, 3.186781e-05, 3.186777e-05, 3.186793e-05, 
    3.186782e-05, 3.1868e-05, 3.186795e-05, 3.186833e-05, 3.186847e-05, 
    3.186853e-05, 3.186859e-05, 3.186872e-05, 3.186863e-05, 3.186866e-05, 
    3.186858e-05, 3.186852e-05, 3.186855e-05, 3.186839e-05, 3.186845e-05, 
    3.186811e-05, 3.186826e-05, 3.186788e-05, 3.186797e-05, 3.186786e-05, 
    3.186792e-05, 3.186782e-05, 3.18679e-05, 3.186776e-05, 3.186772e-05, 
    3.186774e-05, 3.186766e-05, 3.186791e-05, 3.186781e-05, 3.186855e-05, 
    3.186855e-05, 3.186853e-05, 3.186861e-05, 3.186862e-05, 3.18687e-05, 
    3.186863e-05, 3.18686e-05, 3.186852e-05, 3.186847e-05, 3.186843e-05, 
    3.186833e-05, 3.186823e-05, 3.186807e-05, 3.186797e-05, 3.186789e-05, 
    3.186794e-05, 3.18679e-05, 3.186794e-05, 3.186796e-05, 3.186773e-05, 
    3.186786e-05, 3.186767e-05, 3.186768e-05, 3.186777e-05, 3.186768e-05, 
    3.186854e-05, 3.186857e-05, 3.186865e-05, 3.186859e-05, 3.186871e-05, 
    3.186864e-05, 3.18686e-05, 3.186845e-05, 3.186841e-05, 3.186838e-05, 
    3.186832e-05, 3.186824e-05, 3.18681e-05, 3.186798e-05, 3.186787e-05, 
    3.186788e-05, 3.186788e-05, 3.186785e-05, 3.186791e-05, 3.186784e-05, 
    3.186783e-05, 3.186786e-05, 3.186768e-05, 3.186773e-05, 3.186768e-05, 
    3.186772e-05, 3.186856e-05, 3.186852e-05, 3.186854e-05, 3.18685e-05, 
    3.186853e-05, 3.186839e-05, 3.186835e-05, 3.186817e-05, 3.186824e-05, 
    3.186812e-05, 3.186823e-05, 3.186821e-05, 3.186812e-05, 3.186823e-05, 
    3.186799e-05, 3.186815e-05, 3.186785e-05, 3.186801e-05, 3.186784e-05, 
    3.186787e-05, 3.186782e-05, 3.186778e-05, 3.186772e-05, 3.186761e-05, 
    3.186764e-05, 3.186755e-05, 3.186845e-05, 3.18684e-05, 3.186841e-05, 
    3.186835e-05, 3.186831e-05, 3.186821e-05, 3.186807e-05, 3.186812e-05, 
    3.186802e-05, 3.1868e-05, 3.186816e-05, 3.186806e-05, 3.186836e-05, 
    3.186832e-05, 3.186835e-05, 3.186845e-05, 3.186811e-05, 3.186829e-05, 
    3.186796e-05, 3.186806e-05, 3.186778e-05, 3.186792e-05, 3.186765e-05, 
    3.186754e-05, 3.186743e-05, 3.18673e-05, 3.186837e-05, 3.186841e-05, 
    3.186834e-05, 3.186825e-05, 3.186816e-05, 3.186805e-05, 3.186804e-05, 
    3.186802e-05, 3.186796e-05, 3.186792e-05, 3.186801e-05, 3.186791e-05, 
    3.186831e-05, 3.186809e-05, 3.186842e-05, 3.186832e-05, 3.186825e-05, 
    3.186829e-05, 3.186813e-05, 3.186809e-05, 3.186794e-05, 3.186802e-05, 
    3.186757e-05, 3.186777e-05, 3.186721e-05, 3.186736e-05, 3.186842e-05, 
    3.186837e-05, 3.18682e-05, 3.186828e-05, 3.186804e-05, 3.186798e-05, 
    3.186794e-05, 3.186788e-05, 3.186787e-05, 3.186784e-05, 3.186789e-05, 
    3.186784e-05, 3.186805e-05, 3.186796e-05, 3.186822e-05, 3.186815e-05, 
    3.186818e-05, 3.186821e-05, 3.186812e-05, 3.186801e-05, 3.186801e-05, 
    3.186797e-05, 3.186788e-05, 3.186804e-05, 3.186754e-05, 3.186785e-05, 
    3.186832e-05, 3.186822e-05, 3.186821e-05, 3.186824e-05, 3.186799e-05, 
    3.186808e-05, 3.186784e-05, 3.18679e-05, 3.18678e-05, 3.186785e-05, 
    3.186786e-05, 3.186793e-05, 3.186797e-05, 3.186808e-05, 3.186817e-05, 
    3.186824e-05, 3.186822e-05, 3.186815e-05, 3.1868e-05, 3.186787e-05, 
    3.18679e-05, 3.18678e-05, 3.186806e-05, 3.186795e-05, 3.1868e-05, 
    3.186789e-05, 3.186812e-05, 3.186792e-05, 3.186818e-05, 3.186816e-05, 
    3.186809e-05, 3.186794e-05, 3.186792e-05, 3.186788e-05, 3.18679e-05, 
    3.1868e-05, 3.186802e-05, 3.186809e-05, 3.18681e-05, 3.186816e-05, 
    3.18682e-05, 3.186816e-05, 3.186812e-05, 3.1868e-05, 3.186789e-05, 
    3.186777e-05, 3.186775e-05, 3.186761e-05, 3.186772e-05, 3.186754e-05, 
    3.186769e-05, 3.186742e-05, 3.186791e-05, 3.18677e-05, 3.186808e-05, 
    3.186804e-05, 3.186797e-05, 3.18678e-05, 3.186789e-05, 3.186778e-05, 
    3.186802e-05, 3.186814e-05, 3.186817e-05, 3.186824e-05, 3.186817e-05, 
    3.186818e-05, 3.186812e-05, 3.186814e-05, 3.1868e-05, 3.186807e-05, 
    3.186786e-05, 3.186778e-05, 3.186756e-05, 3.186742e-05, 3.186729e-05, 
    3.186722e-05, 3.186721e-05, 3.18672e-05 ;

 LITR1C_TO_SOIL1C =
  6.022506e-13, 6.03873e-13, 6.035578e-13, 6.048652e-13, 6.041403e-13, 
    6.04996e-13, 6.025798e-13, 6.039371e-13, 6.030709e-13, 6.02397e-13, 
    6.073986e-13, 6.049235e-13, 6.099672e-13, 6.083915e-13, 6.123468e-13, 
    6.097218e-13, 6.128757e-13, 6.122716e-13, 6.140902e-13, 6.135695e-13, 
    6.15892e-13, 6.143305e-13, 6.170954e-13, 6.155196e-13, 6.15766e-13, 
    6.142789e-13, 6.054224e-13, 6.070905e-13, 6.053234e-13, 6.055614e-13, 
    6.054548e-13, 6.041551e-13, 6.034994e-13, 6.021268e-13, 6.023762e-13, 
    6.033844e-13, 6.056685e-13, 6.048938e-13, 6.068463e-13, 6.068022e-13, 
    6.089726e-13, 6.079944e-13, 6.116377e-13, 6.106035e-13, 6.135913e-13, 
    6.128402e-13, 6.135559e-13, 6.13339e-13, 6.135587e-13, 6.124572e-13, 
    6.129292e-13, 6.119597e-13, 6.081776e-13, 6.0929e-13, 6.059694e-13, 
    6.039685e-13, 6.026393e-13, 6.01695e-13, 6.018285e-13, 6.020829e-13, 
    6.033903e-13, 6.046189e-13, 6.055545e-13, 6.061799e-13, 6.067959e-13, 
    6.086577e-13, 6.096432e-13, 6.118466e-13, 6.114496e-13, 6.121224e-13, 
    6.127655e-13, 6.138441e-13, 6.136667e-13, 6.141416e-13, 6.12105e-13, 
    6.134587e-13, 6.112233e-13, 6.11835e-13, 6.069616e-13, 6.051029e-13, 
    6.043108e-13, 6.036183e-13, 6.019312e-13, 6.030964e-13, 6.026371e-13, 
    6.037299e-13, 6.044236e-13, 6.040806e-13, 6.06197e-13, 6.053745e-13, 
    6.097017e-13, 6.078394e-13, 6.126906e-13, 6.115311e-13, 6.129684e-13, 
    6.122352e-13, 6.134911e-13, 6.123609e-13, 6.143184e-13, 6.147441e-13, 
    6.144532e-13, 6.155711e-13, 6.122981e-13, 6.135557e-13, 6.040709e-13, 
    6.041269e-13, 6.043876e-13, 6.03241e-13, 6.031709e-13, 6.021199e-13, 
    6.030553e-13, 6.034533e-13, 6.04464e-13, 6.050611e-13, 6.056287e-13, 
    6.068759e-13, 6.082673e-13, 6.102113e-13, 6.116063e-13, 6.125408e-13, 
    6.119679e-13, 6.124737e-13, 6.119082e-13, 6.116432e-13, 6.145845e-13, 
    6.129335e-13, 6.154103e-13, 6.152734e-13, 6.141528e-13, 6.152889e-13, 
    6.041662e-13, 6.038442e-13, 6.027253e-13, 6.03601e-13, 6.020054e-13, 
    6.028985e-13, 6.034117e-13, 6.053913e-13, 6.058263e-13, 6.06229e-13, 
    6.070245e-13, 6.080445e-13, 6.098321e-13, 6.113857e-13, 6.12803e-13, 
    6.126992e-13, 6.127358e-13, 6.13052e-13, 6.122682e-13, 6.131807e-13, 
    6.133337e-13, 6.129335e-13, 6.152551e-13, 6.145922e-13, 6.152705e-13, 
    6.14839e-13, 6.039489e-13, 6.044907e-13, 6.041979e-13, 6.047483e-13, 
    6.043604e-13, 6.060838e-13, 6.066001e-13, 6.090141e-13, 6.080243e-13, 
    6.095998e-13, 6.081846e-13, 6.084353e-13, 6.096505e-13, 6.082612e-13, 
    6.112997e-13, 6.092398e-13, 6.130643e-13, 6.110091e-13, 6.13193e-13, 
    6.127969e-13, 6.134529e-13, 6.1404e-13, 6.147785e-13, 6.161398e-13, 
    6.158247e-13, 6.169627e-13, 6.052981e-13, 6.06e-13, 6.059385e-13, 
    6.06673e-13, 6.072158e-13, 6.083921e-13, 6.102765e-13, 6.095683e-13, 
    6.108686e-13, 6.11129e-13, 6.09154e-13, 6.103668e-13, 6.064698e-13, 
    6.070998e-13, 6.06725e-13, 6.053533e-13, 6.097311e-13, 6.074858e-13, 
    6.116292e-13, 6.104153e-13, 6.139562e-13, 6.121958e-13, 6.156512e-13, 
    6.171251e-13, 6.185123e-13, 6.2013e-13, 6.063833e-13, 6.059065e-13, 
    6.067604e-13, 6.079404e-13, 6.090353e-13, 6.104893e-13, 6.106382e-13, 
    6.109102e-13, 6.116149e-13, 6.122073e-13, 6.10996e-13, 6.123558e-13, 
    6.072453e-13, 6.09926e-13, 6.057259e-13, 6.069915e-13, 6.07871e-13, 
    6.074856e-13, 6.094874e-13, 6.099588e-13, 6.11872e-13, 6.108836e-13, 
    6.167611e-13, 6.141635e-13, 6.213615e-13, 6.193534e-13, 6.057398e-13, 
    6.063818e-13, 6.086136e-13, 6.075521e-13, 6.105865e-13, 6.113319e-13, 
    6.119382e-13, 6.127124e-13, 6.127962e-13, 6.132547e-13, 6.125032e-13, 
    6.132251e-13, 6.104924e-13, 6.117141e-13, 6.08359e-13, 6.091762e-13, 
    6.088004e-13, 6.083879e-13, 6.096607e-13, 6.110147e-13, 6.110441e-13, 
    6.11478e-13, 6.126991e-13, 6.105988e-13, 6.170951e-13, 6.130854e-13, 
    6.070815e-13, 6.083161e-13, 6.084929e-13, 6.080148e-13, 6.112572e-13, 
    6.100833e-13, 6.132436e-13, 6.123901e-13, 6.137884e-13, 6.130937e-13, 
    6.129914e-13, 6.120988e-13, 6.115427e-13, 6.10137e-13, 6.089923e-13, 
    6.080842e-13, 6.082954e-13, 6.092928e-13, 6.110975e-13, 6.128035e-13, 
    6.124299e-13, 6.136822e-13, 6.103666e-13, 6.117573e-13, 6.112197e-13, 
    6.126213e-13, 6.095494e-13, 6.121641e-13, 6.0888e-13, 6.091684e-13, 
    6.1006e-13, 6.118513e-13, 6.122482e-13, 6.126709e-13, 6.124101e-13, 
    6.111435e-13, 6.109364e-13, 6.100384e-13, 6.097902e-13, 6.091056e-13, 
    6.085384e-13, 6.090565e-13, 6.096004e-13, 6.111442e-13, 6.125341e-13, 
    6.140483e-13, 6.144187e-13, 6.161841e-13, 6.147465e-13, 6.171173e-13, 
    6.151008e-13, 6.185902e-13, 6.123162e-13, 6.150425e-13, 6.101007e-13, 
    6.10634e-13, 6.115974e-13, 6.138063e-13, 6.126147e-13, 6.140084e-13, 
    6.109283e-13, 6.09327e-13, 6.08913e-13, 6.081393e-13, 6.089307e-13, 
    6.088664e-13, 6.096232e-13, 6.093801e-13, 6.111954e-13, 6.102207e-13, 
    6.129887e-13, 6.139975e-13, 6.168433e-13, 6.185848e-13, 6.203561e-13, 
    6.211371e-13, 6.213748e-13, 6.214741e-13 ;

 LITR1C_vr =
  0.001819735, 0.001819728, 0.001819729, 0.001819724, 0.001819727, 
    0.001819723, 0.001819734, 0.001819728, 0.001819732, 0.001819735, 
    0.001819712, 0.001819723, 0.001819701, 0.001819708, 0.00181969, 
    0.001819702, 0.001819688, 0.001819691, 0.001819683, 0.001819685, 
    0.001819675, 0.001819682, 0.001819669, 0.001819676, 0.001819675, 
    0.001819682, 0.001819721, 0.001819714, 0.001819722, 0.001819721, 
    0.001819721, 0.001819727, 0.00181973, 0.001819736, 0.001819735, 
    0.00181973, 0.00181972, 0.001819724, 0.001819715, 0.001819715, 
    0.001819705, 0.00181971, 0.001819694, 0.001819698, 0.001819685, 
    0.001819688, 0.001819685, 0.001819686, 0.001819685, 0.00181969, 
    0.001819688, 0.001819692, 0.001819709, 0.001819704, 0.001819719, 
    0.001819728, 0.001819734, 0.001819738, 0.001819737, 0.001819736, 
    0.00181973, 0.001819725, 0.001819721, 0.001819718, 0.001819715, 
    0.001819707, 0.001819702, 0.001819693, 0.001819694, 0.001819692, 
    0.001819689, 0.001819684, 0.001819685, 0.001819683, 0.001819692, 
    0.001819686, 0.001819695, 0.001819693, 0.001819714, 0.001819723, 
    0.001819726, 0.001819729, 0.001819737, 0.001819731, 0.001819734, 
    0.001819729, 0.001819726, 0.001819727, 0.001819718, 0.001819721, 
    0.001819702, 0.00181971, 0.001819689, 0.001819694, 0.001819688, 
    0.001819691, 0.001819685, 0.00181969, 0.001819682, 0.00181968, 
    0.001819681, 0.001819676, 0.001819691, 0.001819685, 0.001819727, 
    0.001819727, 0.001819726, 0.001819731, 0.001819731, 0.001819736, 
    0.001819732, 0.00181973, 0.001819725, 0.001819723, 0.00181972, 
    0.001819715, 0.001819709, 0.0018197, 0.001819694, 0.00181969, 
    0.001819692, 0.00181969, 0.001819692, 0.001819694, 0.001819681, 
    0.001819688, 0.001819677, 0.001819678, 0.001819682, 0.001819677, 
    0.001819727, 0.001819728, 0.001819733, 0.001819729, 0.001819736, 
    0.001819732, 0.00181973, 0.001819721, 0.001819719, 0.001819718, 
    0.001819714, 0.00181971, 0.001819702, 0.001819695, 0.001819688, 
    0.001819689, 0.001819689, 0.001819687, 0.001819691, 0.001819687, 
    0.001819686, 0.001819688, 0.001819678, 0.001819681, 0.001819678, 
    0.001819679, 0.001819728, 0.001819725, 0.001819727, 0.001819724, 
    0.001819726, 0.001819718, 0.001819716, 0.001819705, 0.00181971, 
    0.001819703, 0.001819709, 0.001819708, 0.001819702, 0.001819709, 
    0.001819695, 0.001819704, 0.001819687, 0.001819696, 0.001819687, 
    0.001819688, 0.001819686, 0.001819683, 0.00181968, 0.001819674, 
    0.001819675, 0.00181967, 0.001819722, 0.001819719, 0.001819719, 
    0.001819716, 0.001819713, 0.001819708, 0.0018197, 0.001819703, 
    0.001819697, 0.001819696, 0.001819705, 0.001819699, 0.001819717, 
    0.001819714, 0.001819715, 0.001819721, 0.001819702, 0.001819712, 
    0.001819694, 0.001819699, 0.001819683, 0.001819691, 0.001819676, 
    0.001819669, 0.001819663, 0.001819656, 0.001819717, 0.001819719, 
    0.001819715, 0.00181971, 0.001819705, 0.001819699, 0.001819698, 
    0.001819697, 0.001819694, 0.001819691, 0.001819697, 0.00181969, 
    0.001819713, 0.001819701, 0.00181972, 0.001819714, 0.00181971, 
    0.001819712, 0.001819703, 0.001819701, 0.001819693, 0.001819697, 
    0.001819671, 0.001819682, 0.001819651, 0.001819659, 0.00181972, 
    0.001819717, 0.001819707, 0.001819712, 0.001819698, 0.001819695, 
    0.001819692, 0.001819689, 0.001819688, 0.001819686, 0.00181969, 
    0.001819687, 0.001819699, 0.001819693, 0.001819708, 0.001819705, 
    0.001819706, 0.001819708, 0.001819702, 0.001819696, 0.001819696, 
    0.001819694, 0.001819689, 0.001819698, 0.001819669, 0.001819687, 
    0.001819714, 0.001819708, 0.001819708, 0.00181971, 0.001819695, 
    0.0018197, 0.001819686, 0.00181969, 0.001819684, 0.001819687, 
    0.001819688, 0.001819692, 0.001819694, 0.0018197, 0.001819705, 
    0.001819709, 0.001819708, 0.001819704, 0.001819696, 0.001819688, 
    0.00181969, 0.001819685, 0.001819699, 0.001819693, 0.001819695, 
    0.001819689, 0.001819703, 0.001819691, 0.001819706, 0.001819705, 
    0.001819701, 0.001819693, 0.001819691, 0.001819689, 0.00181969, 
    0.001819696, 0.001819697, 0.001819701, 0.001819702, 0.001819705, 
    0.001819707, 0.001819705, 0.001819703, 0.001819696, 0.00181969, 
    0.001819683, 0.001819681, 0.001819673, 0.00181968, 0.001819669, 
    0.001819678, 0.001819663, 0.001819691, 0.001819678, 0.0018197, 
    0.001819698, 0.001819694, 0.001819684, 0.001819689, 0.001819683, 
    0.001819697, 0.001819704, 0.001819706, 0.001819709, 0.001819706, 
    0.001819706, 0.001819703, 0.001819704, 0.001819696, 0.0018197, 
    0.001819688, 0.001819683, 0.001819671, 0.001819663, 0.001819655, 
    0.001819651, 0.00181965, 0.00181965,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  1.011395e-06, 1.011391e-06, 1.011392e-06, 1.011388e-06, 1.01139e-06, 
    1.011388e-06, 1.011394e-06, 1.011391e-06, 1.011393e-06, 1.011394e-06, 
    1.011382e-06, 1.011388e-06, 1.011376e-06, 1.01138e-06, 1.01137e-06, 
    1.011376e-06, 1.011369e-06, 1.01137e-06, 1.011365e-06, 1.011367e-06, 
    1.011361e-06, 1.011365e-06, 1.011358e-06, 1.011362e-06, 1.011361e-06, 
    1.011365e-06, 1.011387e-06, 1.011383e-06, 1.011387e-06, 1.011387e-06, 
    1.011387e-06, 1.01139e-06, 1.011392e-06, 1.011395e-06, 1.011394e-06, 
    1.011392e-06, 1.011386e-06, 1.011388e-06, 1.011383e-06, 1.011383e-06, 
    1.011378e-06, 1.011381e-06, 1.011372e-06, 1.011374e-06, 1.011367e-06, 
    1.011369e-06, 1.011367e-06, 1.011367e-06, 1.011367e-06, 1.01137e-06, 
    1.011368e-06, 1.011371e-06, 1.01138e-06, 1.011377e-06, 1.011386e-06, 
    1.011391e-06, 1.011394e-06, 1.011396e-06, 1.011396e-06, 1.011395e-06, 
    1.011392e-06, 1.011389e-06, 1.011387e-06, 1.011385e-06, 1.011383e-06, 
    1.011379e-06, 1.011377e-06, 1.011371e-06, 1.011372e-06, 1.01137e-06, 
    1.011369e-06, 1.011366e-06, 1.011367e-06, 1.011365e-06, 1.01137e-06, 
    1.011367e-06, 1.011373e-06, 1.011371e-06, 1.011383e-06, 1.011388e-06, 
    1.01139e-06, 1.011391e-06, 1.011396e-06, 1.011393e-06, 1.011394e-06, 
    1.011391e-06, 1.011389e-06, 1.01139e-06, 1.011385e-06, 1.011387e-06, 
    1.011376e-06, 1.011381e-06, 1.011369e-06, 1.011372e-06, 1.011368e-06, 
    1.01137e-06, 1.011367e-06, 1.01137e-06, 1.011365e-06, 1.011364e-06, 
    1.011365e-06, 1.011362e-06, 1.01137e-06, 1.011367e-06, 1.01139e-06, 
    1.01139e-06, 1.011389e-06, 1.011392e-06, 1.011392e-06, 1.011395e-06, 
    1.011393e-06, 1.011392e-06, 1.011389e-06, 1.011388e-06, 1.011386e-06, 
    1.011383e-06, 1.01138e-06, 1.011375e-06, 1.011372e-06, 1.011369e-06, 
    1.011371e-06, 1.011369e-06, 1.011371e-06, 1.011372e-06, 1.011364e-06, 
    1.011368e-06, 1.011362e-06, 1.011363e-06, 1.011365e-06, 1.011363e-06, 
    1.01139e-06, 1.011391e-06, 1.011394e-06, 1.011391e-06, 1.011395e-06, 
    1.011393e-06, 1.011392e-06, 1.011387e-06, 1.011386e-06, 1.011385e-06, 
    1.011383e-06, 1.01138e-06, 1.011376e-06, 1.011372e-06, 1.011369e-06, 
    1.011369e-06, 1.011369e-06, 1.011368e-06, 1.01137e-06, 1.011368e-06, 
    1.011367e-06, 1.011368e-06, 1.011363e-06, 1.011364e-06, 1.011363e-06, 
    1.011364e-06, 1.011391e-06, 1.011389e-06, 1.01139e-06, 1.011389e-06, 
    1.011389e-06, 1.011385e-06, 1.011384e-06, 1.011378e-06, 1.011381e-06, 
    1.011377e-06, 1.01138e-06, 1.011379e-06, 1.011376e-06, 1.01138e-06, 
    1.011372e-06, 1.011377e-06, 1.011368e-06, 1.011373e-06, 1.011368e-06, 
    1.011369e-06, 1.011367e-06, 1.011366e-06, 1.011364e-06, 1.01136e-06, 
    1.011361e-06, 1.011358e-06, 1.011387e-06, 1.011386e-06, 1.011386e-06, 
    1.011384e-06, 1.011382e-06, 1.01138e-06, 1.011375e-06, 1.011377e-06, 
    1.011373e-06, 1.011373e-06, 1.011378e-06, 1.011375e-06, 1.011384e-06, 
    1.011383e-06, 1.011384e-06, 1.011387e-06, 1.011376e-06, 1.011382e-06, 
    1.011372e-06, 1.011375e-06, 1.011366e-06, 1.01137e-06, 1.011362e-06, 
    1.011358e-06, 1.011355e-06, 1.011351e-06, 1.011384e-06, 1.011386e-06, 
    1.011384e-06, 1.011381e-06, 1.011378e-06, 1.011374e-06, 1.011374e-06, 
    1.011373e-06, 1.011372e-06, 1.01137e-06, 1.011373e-06, 1.01137e-06, 
    1.011382e-06, 1.011376e-06, 1.011386e-06, 1.011383e-06, 1.011381e-06, 
    1.011382e-06, 1.011377e-06, 1.011376e-06, 1.011371e-06, 1.011373e-06, 
    1.011359e-06, 1.011365e-06, 1.011348e-06, 1.011353e-06, 1.011386e-06, 
    1.011384e-06, 1.011379e-06, 1.011382e-06, 1.011374e-06, 1.011372e-06, 
    1.011371e-06, 1.011369e-06, 1.011369e-06, 1.011368e-06, 1.011369e-06, 
    1.011368e-06, 1.011374e-06, 1.011371e-06, 1.01138e-06, 1.011378e-06, 
    1.011379e-06, 1.01138e-06, 1.011376e-06, 1.011373e-06, 1.011373e-06, 
    1.011372e-06, 1.011369e-06, 1.011374e-06, 1.011358e-06, 1.011368e-06, 
    1.011383e-06, 1.01138e-06, 1.011379e-06, 1.011381e-06, 1.011373e-06, 
    1.011375e-06, 1.011368e-06, 1.01137e-06, 1.011366e-06, 1.011368e-06, 
    1.011368e-06, 1.01137e-06, 1.011372e-06, 1.011375e-06, 1.011378e-06, 
    1.01138e-06, 1.01138e-06, 1.011377e-06, 1.011373e-06, 1.011369e-06, 
    1.01137e-06, 1.011367e-06, 1.011375e-06, 1.011371e-06, 1.011373e-06, 
    1.011369e-06, 1.011377e-06, 1.01137e-06, 1.011378e-06, 1.011378e-06, 
    1.011376e-06, 1.011371e-06, 1.01137e-06, 1.011369e-06, 1.01137e-06, 
    1.011373e-06, 1.011373e-06, 1.011376e-06, 1.011376e-06, 1.011378e-06, 
    1.011379e-06, 1.011378e-06, 1.011377e-06, 1.011373e-06, 1.011369e-06, 
    1.011366e-06, 1.011365e-06, 1.01136e-06, 1.011364e-06, 1.011358e-06, 
    1.011363e-06, 1.011354e-06, 1.01137e-06, 1.011363e-06, 1.011375e-06, 
    1.011374e-06, 1.011372e-06, 1.011366e-06, 1.011369e-06, 1.011366e-06, 
    1.011373e-06, 1.011377e-06, 1.011378e-06, 1.01138e-06, 1.011378e-06, 
    1.011378e-06, 1.011377e-06, 1.011377e-06, 1.011373e-06, 1.011375e-06, 
    1.011368e-06, 1.011366e-06, 1.011359e-06, 1.011354e-06, 1.01135e-06, 
    1.011348e-06, 1.011348e-06, 1.011347e-06 ;

 LITR1N_TNDNCY_VERT_TRANS =
  -3.921449e-25, -2.058761e-25, 6.176282e-25, 1.176435e-25, -5.784137e-25, 
    -4.215557e-25, -9.803622e-27, -1.56858e-25, 1.862688e-25, -1.225453e-24, 
    2.843051e-25, 6.862535e-26, -4.41163e-25, -2.843051e-25, -3.431268e-25, 
    4.901811e-26, 4.509666e-25, 1.56858e-25, -3.529304e-25, 3.921449e-25, 
    6.176282e-25, -2.745014e-25, 1.176435e-25, 2.941087e-25, 2.843051e-25, 
    -9.117368e-25, 3.333231e-25, -2.745014e-25, 3.921449e-26, 3.823413e-25, 
    4.509666e-25, 4.901811e-25, -2.156797e-25, -9.803622e-27, 1.470543e-25, 
    2.254833e-25, 9.901658e-25, 3.333231e-25, -3.137159e-25, -2.450906e-25, 
    -1.372507e-25, 2.941087e-25, 5.882173e-25, 3.823413e-25, -6.862535e-26, 
    9.803622e-26, -9.803622e-26, 2.843051e-25, -2.156797e-25, -8.333079e-25, 
    3.529304e-25, 3.137159e-25, 5.293956e-25, -3.529304e-25, 2.058761e-25, 
    5.588064e-25, 2.646978e-25, -4.41163e-25, 5.882173e-25, 5.882173e-26, 
    -3.823413e-25, 1.019577e-24, 1.764652e-25, 4.705739e-25, 2.156797e-25, 
    2.941087e-26, -3.235195e-25, -8.137007e-25, -2.843051e-25, -3.333231e-25, 
    -5.19592e-25, 2.548942e-25, 7.058608e-25, 2.941087e-25, 6.47039e-25, 
    5.882173e-26, -2.254833e-25, 2.548942e-25, 2.156797e-25, -1.274471e-25, 
    4.999847e-25, 3.235195e-25, 3.137159e-25, -3.333231e-25, 9.803622e-26, 
    3.823413e-25, 3.62734e-25, 4.803775e-25, 0, 4.313593e-25, -3.62734e-25, 
    -5.686101e-25, 7.842898e-26, 3.921449e-25, 5.882173e-26, 4.999847e-25, 
    5.98021e-25, 7.842898e-26, -5.490028e-25, 2.941087e-25, -4.999847e-25, 
    -4.803775e-25, -3.62734e-25, -3.137159e-25, -1.088202e-24, 4.313593e-25, 
    -7.842898e-25, 1.470543e-25, -6.862535e-25, 1.372507e-25, -7.842898e-26, 
    5.882173e-25, -3.039123e-25, 3.921449e-25, -4.901811e-26, -5.490028e-25, 
    7.25468e-25, -2.254833e-25, 0, 4.509666e-25, -1.960724e-26, 9.803622e-26, 
    -3.235195e-25, 3.725376e-25, -6.47039e-25, 1.107809e-24, -2.646978e-25, 
    -8.82326e-26, 6.47039e-25, 8.137007e-25, -2.843051e-25, -1.764652e-25, 
    -4.509666e-25, 5.784137e-25, 2.254833e-25, 4.509666e-25, -6.862535e-26, 
    1.862688e-25, 1.372507e-25, 4.313593e-25, 4.705739e-25, -2.843051e-25, 
    -2.352869e-25, -9.803622e-26, -9.803622e-27, 2.646978e-25, 2.843051e-25, 
    2.058761e-25, 8.725224e-25, -3.921449e-25, 5.097883e-25, 1.960724e-26, 
    3.529304e-25, -2.156797e-25, -2.254833e-25, -1.960724e-26, -5.882173e-26, 
    -5.097883e-25, 4.509666e-25, 5.097883e-25, 4.117521e-25, -1.098006e-24, 
    1.215649e-24, -5.882173e-26, 2.941087e-25, 9.803622e-26, 1.960724e-26, 
    1.56858e-25, 1.078398e-25, 7.450753e-25, -4.607703e-25, -5.097883e-25, 
    6.862535e-26, -3.823413e-25, -3.823413e-25, 3.137159e-25, -9.803622e-26, 
    5.882173e-26, 6.764499e-25, 2.058761e-25, 1.470543e-25, -3.333231e-25, 
    5.293956e-25, -2.745014e-25, 7.842898e-26, -2.941087e-26, 2.254833e-25, 
    3.039123e-25, 1.078398e-25, 9.313441e-25, -1.960724e-25, 9.803622e-26, 
    1.470543e-25, -2.941087e-26, 8.03897e-25, -5.293956e-25, 3.235195e-25, 
    3.333231e-25, -1.078398e-25, -5.293956e-25, -7.646825e-25, 3.921449e-26, 
    3.921449e-25, -1.862688e-25, -3.921449e-26, 7.352717e-25, -1.960724e-25, 
    -1.960724e-25, -7.156644e-25, 3.333231e-25, -4.999847e-25, 3.137159e-25, 
    -5.097883e-25, -3.62734e-25, 7.842898e-26, -2.548942e-25, -2.450906e-25, 
    6.568427e-25, 1.078398e-25, -3.235195e-25, 2.941087e-25, -2.745014e-25, 
    1.274471e-25, -1.078398e-25, -1.862688e-25, -3.333231e-25, 5.98021e-25, 
    2.941087e-25, 8.529151e-25, -1.176435e-25, 7.842898e-25, -7.842898e-26, 
    -4.117521e-25, -1.960724e-26, -5.391992e-25, -2.843051e-25, 2.548942e-25, 
    3.137159e-25, 4.215557e-25, -8.137007e-25, -4.999847e-25, -1.960724e-26, 
    -3.333231e-25, -3.333231e-25, -9.019333e-25, -3.921449e-26, -8.82326e-25, 
    -4.705739e-25, 1.215649e-24, 1.078398e-25, 3.137159e-25, 4.607703e-25, 
    4.41163e-25, -1.088202e-24, 4.901811e-25, 2.058761e-25, -9.803622e-26, 
    -7.842898e-26, 7.352717e-25, -6.764499e-25, -7.352717e-25, -2.646978e-25, 
    4.607703e-25, 7.156644e-25, -2.745014e-25, -6.274318e-25, 3.921449e-26, 
    -8.82326e-26, -1.56858e-25, -2.843051e-25, 1.960724e-25, -9.803622e-26, 
    -7.450753e-25, 4.509666e-25, 1.372507e-25, -1.039184e-24, 3.62734e-25, 
    -5.097883e-25, -6.078246e-25, -4.117521e-25, -4.901811e-26, 
    -3.137159e-25, -2.352869e-25, -2.745014e-25, 1.960724e-25, 2.352869e-25, 
    -4.999847e-25, -5.882173e-25, -3.823413e-25, -1.176435e-25, 4.901811e-26, 
    4.901811e-26, -5.490028e-25, -5.882173e-26, 2.450906e-25, 8.137007e-25, 
    -2.450906e-25, 4.999847e-25, 1.960724e-25, 6.862535e-25, -2.745014e-25, 
    -5.588064e-25, 1.058791e-24, 5.19592e-25, 7.156644e-25, -5.98021e-25, 
    1.372507e-25, 7.842898e-25, -1.274471e-25, -1.862688e-25, -2.941087e-25, 
    2.548942e-25, -9.509513e-25, 3.039123e-25, 9.313441e-25, -5.391992e-25, 
    1.960724e-26, 8.725224e-25, -4.901811e-25, -4.901811e-26, 4.901811e-26, 
    -4.509666e-25, -7.842898e-26, -4.803775e-25, -3.529304e-25, 3.431268e-25, 
    6.176282e-25, 8.235043e-25, -2.646978e-25, -2.450906e-25, -6.078246e-25, 
    1.401918e-24, 1.225453e-24, -7.842898e-26, -4.019485e-25, -3.235195e-25, 
    -2.156797e-25, 2.941087e-26,
  9.819556e-32, 9.819516e-32, 9.819524e-32, 9.819491e-32, 9.819509e-32, 
    9.819488e-32, 9.819548e-32, 9.819514e-32, 9.819536e-32, 9.819553e-32, 
    9.819429e-32, 9.81949e-32, 9.819365e-32, 9.819404e-32, 9.819306e-32, 
    9.819371e-32, 9.819293e-32, 9.819308e-32, 9.819263e-32, 9.819276e-32, 
    9.819218e-32, 9.819257e-32, 9.819188e-32, 9.819228e-32, 9.819221e-32, 
    9.819258e-32, 9.819477e-32, 9.819436e-32, 9.81948e-32, 9.819474e-32, 
    9.819477e-32, 9.819509e-32, 9.819525e-32, 9.819559e-32, 9.819553e-32, 
    9.819528e-32, 9.819471e-32, 9.81949e-32, 9.819442e-32, 9.819443e-32, 
    9.81939e-32, 9.819414e-32, 9.819323e-32, 9.819349e-32, 9.819275e-32, 
    9.819294e-32, 9.819276e-32, 9.819282e-32, 9.819276e-32, 9.819303e-32, 
    9.819292e-32, 9.819316e-32, 9.819409e-32, 9.819382e-32, 9.819464e-32, 
    9.819513e-32, 9.819546e-32, 9.81957e-32, 9.819567e-32, 9.81956e-32, 
    9.819528e-32, 9.819497e-32, 9.819474e-32, 9.819459e-32, 9.819443e-32, 
    9.819397e-32, 9.819373e-32, 9.819318e-32, 9.819328e-32, 9.819312e-32, 
    9.819296e-32, 9.819269e-32, 9.819273e-32, 9.819262e-32, 9.819312e-32, 
    9.819279e-32, 9.819334e-32, 9.819319e-32, 9.819439e-32, 9.819486e-32, 
    9.819505e-32, 9.819522e-32, 9.819564e-32, 9.819535e-32, 9.819546e-32, 
    9.819519e-32, 9.819502e-32, 9.819511e-32, 9.819458e-32, 9.819479e-32, 
    9.819372e-32, 9.819417e-32, 9.819298e-32, 9.819326e-32, 9.81929e-32, 
    9.819309e-32, 9.819278e-32, 9.819306e-32, 9.819257e-32, 9.819246e-32, 
    9.819254e-32, 9.819226e-32, 9.819307e-32, 9.819276e-32, 9.819511e-32, 
    9.81951e-32, 9.819503e-32, 9.819531e-32, 9.819533e-32, 9.819559e-32, 
    9.819536e-32, 9.819526e-32, 9.819501e-32, 9.819486e-32, 9.819472e-32, 
    9.819442e-32, 9.819407e-32, 9.819359e-32, 9.819325e-32, 9.819301e-32, 
    9.819315e-32, 9.819303e-32, 9.819317e-32, 9.819323e-32, 9.81925e-32, 
    9.819292e-32, 9.81923e-32, 9.819233e-32, 9.819261e-32, 9.819233e-32, 
    9.819509e-32, 9.819517e-32, 9.819544e-32, 9.819523e-32, 9.819562e-32, 
    9.81954e-32, 9.819527e-32, 9.819478e-32, 9.819467e-32, 9.819457e-32, 
    9.819438e-32, 9.819413e-32, 9.819368e-32, 9.81933e-32, 9.819295e-32, 
    9.819298e-32, 9.819296e-32, 9.819289e-32, 9.819308e-32, 9.819285e-32, 
    9.819282e-32, 9.819292e-32, 9.819234e-32, 9.81925e-32, 9.819233e-32, 
    9.819244e-32, 9.819514e-32, 9.8195e-32, 9.819508e-32, 9.819494e-32, 
    9.819504e-32, 9.819461e-32, 9.819448e-32, 9.819389e-32, 9.819413e-32, 
    9.819374e-32, 9.819409e-32, 9.819403e-32, 9.819373e-32, 9.819407e-32, 
    9.819332e-32, 9.819383e-32, 9.819288e-32, 9.819339e-32, 9.819285e-32, 
    9.819295e-32, 9.819279e-32, 9.819264e-32, 9.819246e-32, 9.819212e-32, 
    9.81922e-32, 9.819192e-32, 9.81948e-32, 9.819463e-32, 9.819464e-32, 
    9.819446e-32, 9.819433e-32, 9.819404e-32, 9.819357e-32, 9.819375e-32, 
    9.819343e-32, 9.819336e-32, 9.819385e-32, 9.819355e-32, 9.819452e-32, 
    9.819436e-32, 9.819445e-32, 9.819479e-32, 9.819371e-32, 9.819426e-32, 
    9.819324e-32, 9.819354e-32, 9.819266e-32, 9.81931e-32, 9.819224e-32, 
    9.819188e-32, 9.819154e-32, 9.819114e-32, 9.819454e-32, 9.819466e-32, 
    9.819444e-32, 9.819415e-32, 9.819388e-32, 9.819352e-32, 9.819348e-32, 
    9.819342e-32, 9.819324e-32, 9.819309e-32, 9.819339e-32, 9.819306e-32, 
    9.819432e-32, 9.819366e-32, 9.81947e-32, 9.819439e-32, 9.819417e-32, 
    9.819426e-32, 9.819377e-32, 9.819365e-32, 9.819317e-32, 9.819342e-32, 
    9.819196e-32, 9.819261e-32, 9.819083e-32, 9.819132e-32, 9.81947e-32, 
    9.819454e-32, 9.819399e-32, 9.819424e-32, 9.81935e-32, 9.819331e-32, 
    9.819316e-32, 9.819297e-32, 9.819295e-32, 9.819283e-32, 9.819302e-32, 
    9.819284e-32, 9.819352e-32, 9.819322e-32, 9.819404e-32, 9.819385e-32, 
    9.819394e-32, 9.819404e-32, 9.819373e-32, 9.819339e-32, 9.819338e-32, 
    9.819327e-32, 9.819298e-32, 9.819349e-32, 9.819188e-32, 9.819288e-32, 
    9.819436e-32, 9.819406e-32, 9.819402e-32, 9.819413e-32, 9.819333e-32, 
    9.819362e-32, 9.819284e-32, 9.819305e-32, 9.81927e-32, 9.819288e-32, 
    9.81929e-32, 9.819312e-32, 9.819326e-32, 9.819361e-32, 9.819389e-32, 
    9.819412e-32, 9.819406e-32, 9.819382e-32, 9.819337e-32, 9.819295e-32, 
    9.819304e-32, 9.819273e-32, 9.819355e-32, 9.81932e-32, 9.819334e-32, 
    9.819299e-32, 9.819375e-32, 9.81931e-32, 9.819392e-32, 9.819385e-32, 
    9.819363e-32, 9.819318e-32, 9.819309e-32, 9.819298e-32, 9.819305e-32, 
    9.819336e-32, 9.819341e-32, 9.819363e-32, 9.819369e-32, 9.819386e-32, 
    9.8194e-32, 9.819387e-32, 9.819374e-32, 9.819336e-32, 9.819302e-32, 
    9.819264e-32, 9.819255e-32, 9.819211e-32, 9.819246e-32, 9.819188e-32, 
    9.819238e-32, 9.819151e-32, 9.819307e-32, 9.819239e-32, 9.819362e-32, 
    9.819349e-32, 9.819325e-32, 9.81927e-32, 9.819299e-32, 9.819265e-32, 
    9.819341e-32, 9.819381e-32, 9.819391e-32, 9.81941e-32, 9.81939e-32, 
    9.819392e-32, 9.819373e-32, 9.819379e-32, 9.819335e-32, 9.819359e-32, 
    9.81929e-32, 9.819265e-32, 9.819195e-32, 9.819152e-32, 9.819108e-32, 
    9.819088e-32, 9.819082e-32, 9.81908e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.247364e-14, 4.258806e-14, 4.256583e-14, 4.265804e-14, 4.260691e-14, 
    4.266727e-14, 4.249686e-14, 4.259259e-14, 4.25315e-14, 4.248397e-14, 
    4.283671e-14, 4.266215e-14, 4.301786e-14, 4.290674e-14, 4.318568e-14, 
    4.300055e-14, 4.322298e-14, 4.318038e-14, 4.330864e-14, 4.327191e-14, 
    4.343571e-14, 4.332558e-14, 4.352057e-14, 4.340944e-14, 4.342682e-14, 
    4.332194e-14, 4.269734e-14, 4.281498e-14, 4.269036e-14, 4.270714e-14, 
    4.269962e-14, 4.260796e-14, 4.256172e-14, 4.246492e-14, 4.24825e-14, 
    4.255361e-14, 4.271469e-14, 4.266006e-14, 4.279776e-14, 4.279465e-14, 
    4.294771e-14, 4.287873e-14, 4.313567e-14, 4.306273e-14, 4.327344e-14, 
    4.322048e-14, 4.327095e-14, 4.325565e-14, 4.327115e-14, 4.319346e-14, 
    4.322675e-14, 4.315838e-14, 4.289164e-14, 4.29701e-14, 4.273592e-14, 
    4.25948e-14, 4.250106e-14, 4.243446e-14, 4.244388e-14, 4.246182e-14, 
    4.255402e-14, 4.264068e-14, 4.270665e-14, 4.275076e-14, 4.27942e-14, 
    4.292551e-14, 4.299501e-14, 4.31504e-14, 4.31224e-14, 4.316985e-14, 
    4.321521e-14, 4.329127e-14, 4.327876e-14, 4.331225e-14, 4.316862e-14, 
    4.326409e-14, 4.310644e-14, 4.314958e-14, 4.280589e-14, 4.26748e-14, 
    4.261894e-14, 4.25701e-14, 4.245112e-14, 4.25333e-14, 4.25009e-14, 
    4.257797e-14, 4.26269e-14, 4.260271e-14, 4.275196e-14, 4.269395e-14, 
    4.299913e-14, 4.286779e-14, 4.320992e-14, 4.312815e-14, 4.322952e-14, 
    4.317781e-14, 4.326638e-14, 4.318667e-14, 4.332473e-14, 4.335475e-14, 
    4.333423e-14, 4.341307e-14, 4.318225e-14, 4.327094e-14, 4.260202e-14, 
    4.260597e-14, 4.262436e-14, 4.254349e-14, 4.253855e-14, 4.246443e-14, 
    4.25304e-14, 4.255847e-14, 4.262974e-14, 4.267186e-14, 4.271189e-14, 
    4.279985e-14, 4.289797e-14, 4.303507e-14, 4.313345e-14, 4.319936e-14, 
    4.315896e-14, 4.319463e-14, 4.315475e-14, 4.313606e-14, 4.334349e-14, 
    4.322706e-14, 4.340173e-14, 4.339208e-14, 4.331305e-14, 4.339317e-14, 
    4.260874e-14, 4.258603e-14, 4.250713e-14, 4.256888e-14, 4.245635e-14, 
    4.251934e-14, 4.255553e-14, 4.269514e-14, 4.272582e-14, 4.275422e-14, 
    4.281032e-14, 4.288226e-14, 4.300833e-14, 4.311789e-14, 4.321785e-14, 
    4.321054e-14, 4.321311e-14, 4.323542e-14, 4.318014e-14, 4.324449e-14, 
    4.325528e-14, 4.322706e-14, 4.339078e-14, 4.334404e-14, 4.339187e-14, 
    4.336144e-14, 4.259342e-14, 4.263163e-14, 4.261098e-14, 4.264979e-14, 
    4.262244e-14, 4.274398e-14, 4.27804e-14, 4.295065e-14, 4.288084e-14, 
    4.299195e-14, 4.289214e-14, 4.290982e-14, 4.299552e-14, 4.289754e-14, 
    4.311183e-14, 4.296656e-14, 4.323629e-14, 4.309134e-14, 4.324536e-14, 
    4.321742e-14, 4.326369e-14, 4.330509e-14, 4.335717e-14, 4.345318e-14, 
    4.343096e-14, 4.351122e-14, 4.268857e-14, 4.273807e-14, 4.273374e-14, 
    4.278553e-14, 4.282382e-14, 4.290678e-14, 4.303968e-14, 4.298972e-14, 
    4.308143e-14, 4.30998e-14, 4.296051e-14, 4.304604e-14, 4.27712e-14, 
    4.281564e-14, 4.27892e-14, 4.269246e-14, 4.300121e-14, 4.284286e-14, 
    4.313507e-14, 4.304946e-14, 4.329918e-14, 4.317503e-14, 4.341872e-14, 
    4.352266e-14, 4.36205e-14, 4.373459e-14, 4.27651e-14, 4.273148e-14, 
    4.27917e-14, 4.287492e-14, 4.295214e-14, 4.305468e-14, 4.306518e-14, 
    4.308437e-14, 4.313406e-14, 4.317584e-14, 4.309041e-14, 4.318631e-14, 
    4.282589e-14, 4.301495e-14, 4.271874e-14, 4.280799e-14, 4.287002e-14, 
    4.284284e-14, 4.298402e-14, 4.301726e-14, 4.31522e-14, 4.308249e-14, 
    4.3497e-14, 4.33138e-14, 4.382144e-14, 4.367982e-14, 4.271972e-14, 
    4.2765e-14, 4.29224e-14, 4.284754e-14, 4.306153e-14, 4.311411e-14, 
    4.315687e-14, 4.321146e-14, 4.321737e-14, 4.324971e-14, 4.319671e-14, 
    4.324763e-14, 4.305489e-14, 4.314106e-14, 4.290444e-14, 4.296207e-14, 
    4.293557e-14, 4.290648e-14, 4.299624e-14, 4.309173e-14, 4.30938e-14, 
    4.312441e-14, 4.321053e-14, 4.30624e-14, 4.352056e-14, 4.323777e-14, 
    4.281434e-14, 4.290141e-14, 4.291388e-14, 4.288016e-14, 4.310883e-14, 
    4.302604e-14, 4.324893e-14, 4.318874e-14, 4.328735e-14, 4.323835e-14, 
    4.323114e-14, 4.316819e-14, 4.312897e-14, 4.302984e-14, 4.29491e-14, 
    4.288506e-14, 4.289996e-14, 4.29703e-14, 4.309758e-14, 4.321789e-14, 
    4.319154e-14, 4.327986e-14, 4.304603e-14, 4.314411e-14, 4.310619e-14, 
    4.320504e-14, 4.298839e-14, 4.317279e-14, 4.294119e-14, 4.296152e-14, 
    4.30244e-14, 4.315073e-14, 4.317872e-14, 4.320853e-14, 4.319015e-14, 
    4.310081e-14, 4.308621e-14, 4.302288e-14, 4.300537e-14, 4.29571e-14, 
    4.29171e-14, 4.295363e-14, 4.299199e-14, 4.310086e-14, 4.319889e-14, 
    4.330567e-14, 4.33318e-14, 4.34563e-14, 4.335491e-14, 4.352212e-14, 
    4.33799e-14, 4.3626e-14, 4.318352e-14, 4.337579e-14, 4.302727e-14, 
    4.306489e-14, 4.313283e-14, 4.328861e-14, 4.320457e-14, 4.330286e-14, 
    4.308564e-14, 4.297271e-14, 4.294351e-14, 4.288895e-14, 4.294476e-14, 
    4.294022e-14, 4.29936e-14, 4.297645e-14, 4.310448e-14, 4.303574e-14, 
    4.323095e-14, 4.33021e-14, 4.35028e-14, 4.362561e-14, 4.375053e-14, 
    4.380561e-14, 4.382238e-14, 4.382938e-14 ;

 LITR1N_vr =
  5.775168e-05, 5.775145e-05, 5.77515e-05, 5.775131e-05, 5.775141e-05, 
    5.775129e-05, 5.775164e-05, 5.775144e-05, 5.775157e-05, 5.775166e-05, 
    5.775096e-05, 5.775131e-05, 5.77506e-05, 5.775082e-05, 5.775026e-05, 
    5.775063e-05, 5.775019e-05, 5.775027e-05, 5.775002e-05, 5.775009e-05, 
    5.774976e-05, 5.774998e-05, 5.774959e-05, 5.774981e-05, 5.774978e-05, 
    5.774999e-05, 5.775124e-05, 5.7751e-05, 5.775125e-05, 5.775121e-05, 
    5.775123e-05, 5.775141e-05, 5.775151e-05, 5.77517e-05, 5.775167e-05, 
    5.775152e-05, 5.77512e-05, 5.775131e-05, 5.775104e-05, 5.775104e-05, 
    5.775074e-05, 5.775087e-05, 5.775036e-05, 5.775051e-05, 5.775009e-05, 
    5.775019e-05, 5.775009e-05, 5.775012e-05, 5.775009e-05, 5.775025e-05, 
    5.775018e-05, 5.775032e-05, 5.775085e-05, 5.775069e-05, 5.775116e-05, 
    5.775144e-05, 5.775163e-05, 5.775176e-05, 5.775174e-05, 5.775171e-05, 
    5.775152e-05, 5.775135e-05, 5.775122e-05, 5.775113e-05, 5.775104e-05, 
    5.775078e-05, 5.775064e-05, 5.775033e-05, 5.775039e-05, 5.775029e-05, 
    5.77502e-05, 5.775005e-05, 5.775008e-05, 5.775001e-05, 5.775029e-05, 
    5.775011e-05, 5.775042e-05, 5.775033e-05, 5.775102e-05, 5.775128e-05, 
    5.775139e-05, 5.775149e-05, 5.775173e-05, 5.775156e-05, 5.775163e-05, 
    5.775147e-05, 5.775138e-05, 5.775143e-05, 5.775113e-05, 5.775124e-05, 
    5.775063e-05, 5.775089e-05, 5.775021e-05, 5.775038e-05, 5.775017e-05, 
    5.775028e-05, 5.77501e-05, 5.775026e-05, 5.774998e-05, 5.774992e-05, 
    5.774997e-05, 5.774981e-05, 5.775027e-05, 5.775009e-05, 5.775143e-05, 
    5.775142e-05, 5.775138e-05, 5.775154e-05, 5.775155e-05, 5.77517e-05, 
    5.775157e-05, 5.775151e-05, 5.775137e-05, 5.775129e-05, 5.775121e-05, 
    5.775103e-05, 5.775084e-05, 5.775056e-05, 5.775037e-05, 5.775024e-05, 
    5.775032e-05, 5.775024e-05, 5.775032e-05, 5.775036e-05, 5.774994e-05, 
    5.775018e-05, 5.774983e-05, 5.774985e-05, 5.775001e-05, 5.774985e-05, 
    5.775141e-05, 5.775146e-05, 5.775161e-05, 5.775149e-05, 5.775172e-05, 
    5.775159e-05, 5.775152e-05, 5.775124e-05, 5.775118e-05, 5.775112e-05, 
    5.775101e-05, 5.775087e-05, 5.775061e-05, 5.77504e-05, 5.77502e-05, 
    5.775021e-05, 5.775021e-05, 5.775016e-05, 5.775027e-05, 5.775015e-05, 
    5.775012e-05, 5.775018e-05, 5.774985e-05, 5.774994e-05, 5.774985e-05, 
    5.774991e-05, 5.775144e-05, 5.775137e-05, 5.775141e-05, 5.775133e-05, 
    5.775139e-05, 5.775114e-05, 5.775107e-05, 5.775073e-05, 5.775087e-05, 
    5.775065e-05, 5.775085e-05, 5.775081e-05, 5.775064e-05, 5.775084e-05, 
    5.775041e-05, 5.77507e-05, 5.775016e-05, 5.775045e-05, 5.775014e-05, 
    5.77502e-05, 5.775011e-05, 5.775003e-05, 5.774992e-05, 5.774973e-05, 
    5.774977e-05, 5.774961e-05, 5.775125e-05, 5.775116e-05, 5.775116e-05, 
    5.775106e-05, 5.775099e-05, 5.775082e-05, 5.775055e-05, 5.775065e-05, 
    5.775047e-05, 5.775043e-05, 5.775071e-05, 5.775054e-05, 5.775109e-05, 
    5.7751e-05, 5.775105e-05, 5.775125e-05, 5.775063e-05, 5.775095e-05, 
    5.775036e-05, 5.775053e-05, 5.775004e-05, 5.775028e-05, 5.77498e-05, 
    5.774959e-05, 5.77494e-05, 5.774917e-05, 5.77511e-05, 5.775117e-05, 
    5.775105e-05, 5.775088e-05, 5.775073e-05, 5.775052e-05, 5.77505e-05, 
    5.775047e-05, 5.775036e-05, 5.775028e-05, 5.775045e-05, 5.775026e-05, 
    5.775098e-05, 5.77506e-05, 5.775119e-05, 5.775101e-05, 5.775089e-05, 
    5.775095e-05, 5.775067e-05, 5.77506e-05, 5.775033e-05, 5.775047e-05, 
    5.774964e-05, 5.775001e-05, 5.774899e-05, 5.774928e-05, 5.775119e-05, 
    5.77511e-05, 5.775079e-05, 5.775093e-05, 5.775051e-05, 5.77504e-05, 
    5.775032e-05, 5.775021e-05, 5.77502e-05, 5.775013e-05, 5.775024e-05, 
    5.775014e-05, 5.775052e-05, 5.775035e-05, 5.775082e-05, 5.775071e-05, 
    5.775076e-05, 5.775082e-05, 5.775064e-05, 5.775045e-05, 5.775044e-05, 
    5.775039e-05, 5.775021e-05, 5.775051e-05, 5.774959e-05, 5.775016e-05, 
    5.7751e-05, 5.775083e-05, 5.77508e-05, 5.775087e-05, 5.775041e-05, 
    5.775058e-05, 5.775013e-05, 5.775025e-05, 5.775006e-05, 5.775016e-05, 
    5.775017e-05, 5.77503e-05, 5.775037e-05, 5.775057e-05, 5.775073e-05, 
    5.775086e-05, 5.775083e-05, 5.775069e-05, 5.775044e-05, 5.77502e-05, 
    5.775025e-05, 5.775007e-05, 5.775054e-05, 5.775035e-05, 5.775042e-05, 
    5.775022e-05, 5.775065e-05, 5.775029e-05, 5.775075e-05, 5.775071e-05, 
    5.775058e-05, 5.775033e-05, 5.775028e-05, 5.775021e-05, 5.775025e-05, 
    5.775043e-05, 5.775046e-05, 5.775059e-05, 5.775062e-05, 5.775072e-05, 
    5.77508e-05, 5.775072e-05, 5.775065e-05, 5.775043e-05, 5.775024e-05, 
    5.775002e-05, 5.774997e-05, 5.774972e-05, 5.774992e-05, 5.774959e-05, 
    5.774987e-05, 5.774938e-05, 5.775027e-05, 5.774988e-05, 5.775058e-05, 
    5.77505e-05, 5.775037e-05, 5.775006e-05, 5.775023e-05, 5.775003e-05, 
    5.775046e-05, 5.775069e-05, 5.775075e-05, 5.775085e-05, 5.775074e-05, 
    5.775075e-05, 5.775064e-05, 5.775068e-05, 5.775043e-05, 5.775056e-05, 
    5.775017e-05, 5.775003e-05, 5.774963e-05, 5.774938e-05, 5.774913e-05, 
    5.774902e-05, 5.774899e-05, 5.774898e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  7.36084e-13, 7.380669e-13, 7.376818e-13, 7.392797e-13, 7.383937e-13, 
    7.394395e-13, 7.364864e-13, 7.381454e-13, 7.370867e-13, 7.362629e-13, 
    7.42376e-13, 7.39351e-13, 7.455155e-13, 7.435897e-13, 7.484239e-13, 
    7.452155e-13, 7.490703e-13, 7.48332e-13, 7.505547e-13, 7.499182e-13, 
    7.52757e-13, 7.508484e-13, 7.542277e-13, 7.523016e-13, 7.526029e-13, 
    7.507853e-13, 7.399607e-13, 7.419995e-13, 7.398397e-13, 7.401306e-13, 
    7.400002e-13, 7.384118e-13, 7.376104e-13, 7.359327e-13, 7.362375e-13, 
    7.374699e-13, 7.402614e-13, 7.393147e-13, 7.41701e-13, 7.416471e-13, 
    7.442999e-13, 7.431043e-13, 7.475572e-13, 7.462931e-13, 7.499449e-13, 
    7.49027e-13, 7.499017e-13, 7.496365e-13, 7.499051e-13, 7.485588e-13, 
    7.491357e-13, 7.479507e-13, 7.433281e-13, 7.446878e-13, 7.406293e-13, 
    7.381837e-13, 7.365591e-13, 7.35405e-13, 7.355682e-13, 7.358792e-13, 
    7.374771e-13, 7.389787e-13, 7.401221e-13, 7.408865e-13, 7.416394e-13, 
    7.43915e-13, 7.451196e-13, 7.478125e-13, 7.473272e-13, 7.481496e-13, 
    7.489356e-13, 7.502539e-13, 7.500371e-13, 7.506175e-13, 7.481283e-13, 
    7.497828e-13, 7.470506e-13, 7.477983e-13, 7.41842e-13, 7.395702e-13, 
    7.386021e-13, 7.377557e-13, 7.356936e-13, 7.371178e-13, 7.365565e-13, 
    7.378921e-13, 7.3874e-13, 7.383208e-13, 7.409074e-13, 7.399021e-13, 
    7.451909e-13, 7.429147e-13, 7.48844e-13, 7.474269e-13, 7.491836e-13, 
    7.482875e-13, 7.498225e-13, 7.484411e-13, 7.508336e-13, 7.513539e-13, 
    7.509983e-13, 7.523646e-13, 7.483644e-13, 7.499014e-13, 7.383089e-13, 
    7.383773e-13, 7.38696e-13, 7.372946e-13, 7.372089e-13, 7.359243e-13, 
    7.370676e-13, 7.375541e-13, 7.387893e-13, 7.395192e-13, 7.402128e-13, 
    7.417372e-13, 7.434378e-13, 7.458138e-13, 7.475187e-13, 7.48661e-13, 
    7.479608e-13, 7.485789e-13, 7.478878e-13, 7.475639e-13, 7.511588e-13, 
    7.491409e-13, 7.521681e-13, 7.520008e-13, 7.506312e-13, 7.520197e-13, 
    7.384253e-13, 7.380318e-13, 7.366643e-13, 7.377346e-13, 7.357844e-13, 
    7.36876e-13, 7.375032e-13, 7.399227e-13, 7.404544e-13, 7.409466e-13, 
    7.419188e-13, 7.431655e-13, 7.453503e-13, 7.472492e-13, 7.489815e-13, 
    7.488546e-13, 7.488993e-13, 7.492858e-13, 7.483278e-13, 7.494431e-13, 
    7.4963e-13, 7.491409e-13, 7.519784e-13, 7.511683e-13, 7.519973e-13, 
    7.514699e-13, 7.381598e-13, 7.388219e-13, 7.384641e-13, 7.391368e-13, 
    7.386628e-13, 7.407691e-13, 7.414001e-13, 7.443507e-13, 7.431408e-13, 
    7.450664e-13, 7.433367e-13, 7.436432e-13, 7.451284e-13, 7.434303e-13, 
    7.471441e-13, 7.446264e-13, 7.493009e-13, 7.467889e-13, 7.494582e-13, 
    7.48974e-13, 7.497757e-13, 7.504933e-13, 7.51396e-13, 7.530597e-13, 
    7.526747e-13, 7.540655e-13, 7.398088e-13, 7.406667e-13, 7.405916e-13, 
    7.414892e-13, 7.421527e-13, 7.435904e-13, 7.458935e-13, 7.450279e-13, 
    7.466172e-13, 7.469355e-13, 7.445216e-13, 7.46004e-13, 7.412409e-13, 
    7.420109e-13, 7.415528e-13, 7.398763e-13, 7.452269e-13, 7.424827e-13, 
    7.475469e-13, 7.460631e-13, 7.50391e-13, 7.482393e-13, 7.524626e-13, 
    7.542639e-13, 7.559595e-13, 7.579366e-13, 7.411351e-13, 7.405524e-13, 
    7.41596e-13, 7.430383e-13, 7.443765e-13, 7.461536e-13, 7.463355e-13, 
    7.466681e-13, 7.475293e-13, 7.482533e-13, 7.467729e-13, 7.484348e-13, 
    7.421886e-13, 7.454651e-13, 7.403316e-13, 7.418785e-13, 7.429534e-13, 
    7.424824e-13, 7.449291e-13, 7.455051e-13, 7.478436e-13, 7.466355e-13, 
    7.538192e-13, 7.506442e-13, 7.594419e-13, 7.569875e-13, 7.403486e-13, 
    7.411333e-13, 7.43861e-13, 7.425638e-13, 7.462723e-13, 7.471835e-13, 
    7.479245e-13, 7.488707e-13, 7.489731e-13, 7.495335e-13, 7.486151e-13, 
    7.494974e-13, 7.461574e-13, 7.476505e-13, 7.435499e-13, 7.445487e-13, 
    7.440894e-13, 7.435852e-13, 7.451408e-13, 7.467957e-13, 7.468316e-13, 
    7.47362e-13, 7.488544e-13, 7.462874e-13, 7.542274e-13, 7.493266e-13, 
    7.419885e-13, 7.434974e-13, 7.437136e-13, 7.431291e-13, 7.470921e-13, 
    7.456573e-13, 7.4952e-13, 7.484769e-13, 7.501858e-13, 7.493367e-13, 
    7.492118e-13, 7.481207e-13, 7.47441e-13, 7.45723e-13, 7.443239e-13, 
    7.43214e-13, 7.434722e-13, 7.446913e-13, 7.46897e-13, 7.489821e-13, 
    7.485255e-13, 7.50056e-13, 7.460037e-13, 7.477034e-13, 7.470463e-13, 
    7.487593e-13, 7.450048e-13, 7.482005e-13, 7.441867e-13, 7.445391e-13, 
    7.456289e-13, 7.478183e-13, 7.483033e-13, 7.4882e-13, 7.485013e-13, 
    7.469531e-13, 7.467e-13, 7.456025e-13, 7.452991e-13, 7.444624e-13, 
    7.437692e-13, 7.444024e-13, 7.450671e-13, 7.46954e-13, 7.486528e-13, 
    7.505034e-13, 7.509562e-13, 7.531139e-13, 7.513568e-13, 7.542545e-13, 
    7.517899e-13, 7.560548e-13, 7.483865e-13, 7.517186e-13, 7.456786e-13, 
    7.463305e-13, 7.475078e-13, 7.502077e-13, 7.487513e-13, 7.504547e-13, 
    7.466901e-13, 7.447329e-13, 7.44227e-13, 7.432814e-13, 7.442486e-13, 
    7.4417e-13, 7.450951e-13, 7.447979e-13, 7.470167e-13, 7.458254e-13, 
    7.492084e-13, 7.504414e-13, 7.539196e-13, 7.56048e-13, 7.58213e-13, 
    7.591676e-13, 7.594581e-13, 7.595795e-13 ;

 LITR2C =
  2.015622e-05, 2.01562e-05, 2.015621e-05, 2.015619e-05, 2.01562e-05, 
    2.015619e-05, 2.015622e-05, 2.01562e-05, 2.015621e-05, 2.015622e-05, 
    2.015615e-05, 2.015619e-05, 2.015612e-05, 2.015614e-05, 2.015609e-05, 
    2.015613e-05, 2.015608e-05, 2.015609e-05, 2.015607e-05, 2.015607e-05, 
    2.015605e-05, 2.015607e-05, 2.015603e-05, 2.015605e-05, 2.015605e-05, 
    2.015607e-05, 2.015618e-05, 2.015616e-05, 2.015618e-05, 2.015618e-05, 
    2.015618e-05, 2.01562e-05, 2.015621e-05, 2.015622e-05, 2.015622e-05, 
    2.015621e-05, 2.015618e-05, 2.015619e-05, 2.015616e-05, 2.015616e-05, 
    2.015613e-05, 2.015615e-05, 2.01561e-05, 2.015611e-05, 2.015607e-05, 
    2.015609e-05, 2.015607e-05, 2.015608e-05, 2.015607e-05, 2.015609e-05, 
    2.015608e-05, 2.01561e-05, 2.015615e-05, 2.015613e-05, 2.015617e-05, 
    2.01562e-05, 2.015622e-05, 2.015623e-05, 2.015623e-05, 2.015622e-05, 
    2.015621e-05, 2.015619e-05, 2.015618e-05, 2.015617e-05, 2.015616e-05, 
    2.015614e-05, 2.015613e-05, 2.01561e-05, 2.01561e-05, 2.015609e-05, 
    2.015609e-05, 2.015607e-05, 2.015607e-05, 2.015607e-05, 2.015609e-05, 
    2.015608e-05, 2.015611e-05, 2.01561e-05, 2.015616e-05, 2.015619e-05, 
    2.015619e-05, 2.01562e-05, 2.015623e-05, 2.015621e-05, 2.015622e-05, 
    2.01562e-05, 2.015619e-05, 2.01562e-05, 2.015617e-05, 2.015618e-05, 
    2.015613e-05, 2.015615e-05, 2.015609e-05, 2.01561e-05, 2.015608e-05, 
    2.015609e-05, 2.015608e-05, 2.015609e-05, 2.015607e-05, 2.015606e-05, 
    2.015606e-05, 2.015605e-05, 2.015609e-05, 2.015607e-05, 2.01562e-05, 
    2.01562e-05, 2.015619e-05, 2.015621e-05, 2.015621e-05, 2.015622e-05, 
    2.015621e-05, 2.015621e-05, 2.015619e-05, 2.015619e-05, 2.015618e-05, 
    2.015616e-05, 2.015614e-05, 2.015612e-05, 2.01561e-05, 2.015609e-05, 
    2.01561e-05, 2.015609e-05, 2.01561e-05, 2.01561e-05, 2.015606e-05, 
    2.015608e-05, 2.015605e-05, 2.015605e-05, 2.015607e-05, 2.015605e-05, 
    2.01562e-05, 2.01562e-05, 2.015622e-05, 2.015621e-05, 2.015623e-05, 
    2.015621e-05, 2.015621e-05, 2.015618e-05, 2.015618e-05, 2.015617e-05, 
    2.015616e-05, 2.015615e-05, 2.015612e-05, 2.01561e-05, 2.015609e-05, 
    2.015609e-05, 2.015609e-05, 2.015608e-05, 2.015609e-05, 2.015608e-05, 
    2.015608e-05, 2.015608e-05, 2.015605e-05, 2.015606e-05, 2.015605e-05, 
    2.015606e-05, 2.01562e-05, 2.015619e-05, 2.01562e-05, 2.015619e-05, 
    2.015619e-05, 2.015617e-05, 2.015617e-05, 2.015613e-05, 2.015615e-05, 
    2.015613e-05, 2.015615e-05, 2.015614e-05, 2.015613e-05, 2.015614e-05, 
    2.015611e-05, 2.015613e-05, 2.015608e-05, 2.015611e-05, 2.015608e-05, 
    2.015609e-05, 2.015608e-05, 2.015607e-05, 2.015606e-05, 2.015604e-05, 
    2.015605e-05, 2.015603e-05, 2.015618e-05, 2.015617e-05, 2.015617e-05, 
    2.015617e-05, 2.015616e-05, 2.015614e-05, 2.015612e-05, 2.015613e-05, 
    2.015611e-05, 2.015611e-05, 2.015613e-05, 2.015612e-05, 2.015617e-05, 
    2.015616e-05, 2.015616e-05, 2.015618e-05, 2.015613e-05, 2.015615e-05, 
    2.01561e-05, 2.015612e-05, 2.015607e-05, 2.015609e-05, 2.015605e-05, 
    2.015603e-05, 2.015601e-05, 2.015599e-05, 2.015617e-05, 2.015617e-05, 
    2.015616e-05, 2.015615e-05, 2.015613e-05, 2.015611e-05, 2.015611e-05, 
    2.015611e-05, 2.01561e-05, 2.015609e-05, 2.015611e-05, 2.015609e-05, 
    2.015616e-05, 2.015612e-05, 2.015618e-05, 2.015616e-05, 2.015615e-05, 
    2.015615e-05, 2.015613e-05, 2.015612e-05, 2.01561e-05, 2.015611e-05, 
    2.015603e-05, 2.015607e-05, 2.015597e-05, 2.0156e-05, 2.015618e-05, 
    2.015617e-05, 2.015614e-05, 2.015615e-05, 2.015611e-05, 2.01561e-05, 
    2.01561e-05, 2.015609e-05, 2.015609e-05, 2.015608e-05, 2.015609e-05, 
    2.015608e-05, 2.015611e-05, 2.01561e-05, 2.015614e-05, 2.015613e-05, 
    2.015614e-05, 2.015614e-05, 2.015613e-05, 2.015611e-05, 2.015611e-05, 
    2.01561e-05, 2.015609e-05, 2.015611e-05, 2.015603e-05, 2.015608e-05, 
    2.015616e-05, 2.015614e-05, 2.015614e-05, 2.015615e-05, 2.015611e-05, 
    2.015612e-05, 2.015608e-05, 2.015609e-05, 2.015607e-05, 2.015608e-05, 
    2.015608e-05, 2.015609e-05, 2.01561e-05, 2.015612e-05, 2.015613e-05, 
    2.015615e-05, 2.015614e-05, 2.015613e-05, 2.015611e-05, 2.015609e-05, 
    2.015609e-05, 2.015607e-05, 2.015612e-05, 2.01561e-05, 2.015611e-05, 
    2.015609e-05, 2.015613e-05, 2.015609e-05, 2.015614e-05, 2.015613e-05, 
    2.015612e-05, 2.01561e-05, 2.015609e-05, 2.015609e-05, 2.015609e-05, 
    2.015611e-05, 2.015611e-05, 2.015612e-05, 2.015612e-05, 2.015613e-05, 
    2.015614e-05, 2.015613e-05, 2.015613e-05, 2.015611e-05, 2.015609e-05, 
    2.015607e-05, 2.015606e-05, 2.015604e-05, 2.015606e-05, 2.015603e-05, 
    2.015605e-05, 2.015601e-05, 2.015609e-05, 2.015606e-05, 2.015612e-05, 
    2.015611e-05, 2.01561e-05, 2.015607e-05, 2.015609e-05, 2.015607e-05, 
    2.015611e-05, 2.015613e-05, 2.015614e-05, 2.015615e-05, 2.015613e-05, 
    2.015614e-05, 2.015613e-05, 2.015613e-05, 2.015611e-05, 2.015612e-05, 
    2.015608e-05, 2.015607e-05, 2.015603e-05, 2.015601e-05, 2.015599e-05, 
    2.015598e-05, 2.015597e-05, 2.015597e-05 ;

 LITR2C_TO_SOIL1C =
  1.120919e-13, 1.123942e-13, 1.123355e-13, 1.12579e-13, 1.12444e-13, 
    1.126034e-13, 1.121533e-13, 1.124061e-13, 1.122448e-13, 1.121192e-13, 
    1.13051e-13, 1.125899e-13, 1.135296e-13, 1.13236e-13, 1.13973e-13, 
    1.134839e-13, 1.140715e-13, 1.13959e-13, 1.142978e-13, 1.142008e-13, 
    1.146335e-13, 1.143426e-13, 1.148577e-13, 1.145641e-13, 1.1461e-13, 
    1.143329e-13, 1.126829e-13, 1.129936e-13, 1.126644e-13, 1.127088e-13, 
    1.126889e-13, 1.124467e-13, 1.123246e-13, 1.120689e-13, 1.121153e-13, 
    1.123032e-13, 1.127287e-13, 1.125844e-13, 1.129481e-13, 1.129399e-13, 
    1.133443e-13, 1.13162e-13, 1.138408e-13, 1.136482e-13, 1.142048e-13, 
    1.140649e-13, 1.141982e-13, 1.141578e-13, 1.141988e-13, 1.139935e-13, 
    1.140815e-13, 1.139008e-13, 1.131962e-13, 1.134034e-13, 1.127848e-13, 
    1.12412e-13, 1.121643e-13, 1.119884e-13, 1.120133e-13, 1.120607e-13, 
    1.123043e-13, 1.125332e-13, 1.127075e-13, 1.12824e-13, 1.129388e-13, 
    1.132856e-13, 1.134693e-13, 1.138798e-13, 1.138058e-13, 1.139312e-13, 
    1.14051e-13, 1.142519e-13, 1.142189e-13, 1.143074e-13, 1.139279e-13, 
    1.141801e-13, 1.137636e-13, 1.138776e-13, 1.129696e-13, 1.126233e-13, 
    1.124758e-13, 1.123467e-13, 1.120324e-13, 1.122495e-13, 1.121639e-13, 
    1.123675e-13, 1.124968e-13, 1.124329e-13, 1.128272e-13, 1.126739e-13, 
    1.134801e-13, 1.131332e-13, 1.14037e-13, 1.13821e-13, 1.140888e-13, 
    1.139522e-13, 1.141862e-13, 1.139756e-13, 1.143403e-13, 1.144196e-13, 
    1.143654e-13, 1.145737e-13, 1.139639e-13, 1.141982e-13, 1.124311e-13, 
    1.124415e-13, 1.124901e-13, 1.122764e-13, 1.122634e-13, 1.120676e-13, 
    1.122418e-13, 1.12316e-13, 1.125043e-13, 1.126156e-13, 1.127213e-13, 
    1.129537e-13, 1.132129e-13, 1.135751e-13, 1.13835e-13, 1.140091e-13, 
    1.139024e-13, 1.139966e-13, 1.138913e-13, 1.138419e-13, 1.143899e-13, 
    1.140823e-13, 1.145438e-13, 1.145182e-13, 1.143095e-13, 1.145211e-13, 
    1.124488e-13, 1.123888e-13, 1.121804e-13, 1.123435e-13, 1.120462e-13, 
    1.122126e-13, 1.123083e-13, 1.126771e-13, 1.127581e-13, 1.128331e-13, 
    1.129813e-13, 1.131714e-13, 1.135044e-13, 1.137939e-13, 1.14058e-13, 
    1.140386e-13, 1.140454e-13, 1.141044e-13, 1.139583e-13, 1.141283e-13, 
    1.141568e-13, 1.140823e-13, 1.145148e-13, 1.143913e-13, 1.145177e-13, 
    1.144373e-13, 1.124083e-13, 1.125093e-13, 1.124547e-13, 1.125573e-13, 
    1.12485e-13, 1.128061e-13, 1.129023e-13, 1.13352e-13, 1.131676e-13, 
    1.134612e-13, 1.131975e-13, 1.132442e-13, 1.134706e-13, 1.132118e-13, 
    1.137779e-13, 1.133941e-13, 1.141067e-13, 1.137237e-13, 1.141306e-13, 
    1.140568e-13, 1.14179e-13, 1.142884e-13, 1.14426e-13, 1.146797e-13, 
    1.14621e-13, 1.14833e-13, 1.126597e-13, 1.127905e-13, 1.12779e-13, 
    1.129159e-13, 1.13017e-13, 1.132362e-13, 1.135872e-13, 1.134553e-13, 
    1.136976e-13, 1.137461e-13, 1.133781e-13, 1.136041e-13, 1.12878e-13, 
    1.129954e-13, 1.129255e-13, 1.1267e-13, 1.134856e-13, 1.130673e-13, 
    1.138393e-13, 1.136131e-13, 1.142728e-13, 1.139448e-13, 1.145886e-13, 
    1.148632e-13, 1.151217e-13, 1.154231e-13, 1.128619e-13, 1.12773e-13, 
    1.129321e-13, 1.13152e-13, 1.13356e-13, 1.136269e-13, 1.136546e-13, 
    1.137053e-13, 1.138366e-13, 1.13947e-13, 1.137213e-13, 1.139746e-13, 
    1.130225e-13, 1.135219e-13, 1.127394e-13, 1.129752e-13, 1.131391e-13, 
    1.130673e-13, 1.134402e-13, 1.13528e-13, 1.138845e-13, 1.137003e-13, 
    1.147954e-13, 1.143114e-13, 1.156526e-13, 1.152784e-13, 1.12742e-13, 
    1.128616e-13, 1.132774e-13, 1.130797e-13, 1.13645e-13, 1.137839e-13, 
    1.138968e-13, 1.140411e-13, 1.140567e-13, 1.141421e-13, 1.140021e-13, 
    1.141366e-13, 1.136275e-13, 1.138551e-13, 1.1323e-13, 1.133822e-13, 
    1.133122e-13, 1.132354e-13, 1.134725e-13, 1.137248e-13, 1.137302e-13, 
    1.138111e-13, 1.140386e-13, 1.136473e-13, 1.148577e-13, 1.141106e-13, 
    1.12992e-13, 1.13222e-13, 1.132549e-13, 1.131658e-13, 1.1377e-13, 
    1.135512e-13, 1.1414e-13, 1.13981e-13, 1.142416e-13, 1.141121e-13, 
    1.140931e-13, 1.139268e-13, 1.138231e-13, 1.135613e-13, 1.13348e-13, 
    1.131788e-13, 1.132181e-13, 1.13404e-13, 1.137402e-13, 1.140581e-13, 
    1.139884e-13, 1.142218e-13, 1.13604e-13, 1.138631e-13, 1.13763e-13, 
    1.140241e-13, 1.134518e-13, 1.139389e-13, 1.133271e-13, 1.133808e-13, 
    1.135469e-13, 1.138807e-13, 1.139546e-13, 1.140333e-13, 1.139848e-13, 
    1.137488e-13, 1.137102e-13, 1.135429e-13, 1.134966e-13, 1.133691e-13, 
    1.132634e-13, 1.133599e-13, 1.134613e-13, 1.137489e-13, 1.140079e-13, 
    1.1429e-13, 1.14359e-13, 1.146879e-13, 1.144201e-13, 1.148618e-13, 
    1.144861e-13, 1.151362e-13, 1.139673e-13, 1.144752e-13, 1.135545e-13, 
    1.136539e-13, 1.138333e-13, 1.142449e-13, 1.140229e-13, 1.142826e-13, 
    1.137087e-13, 1.134103e-13, 1.133332e-13, 1.131891e-13, 1.133365e-13, 
    1.133245e-13, 1.134655e-13, 1.134202e-13, 1.137584e-13, 1.135769e-13, 
    1.140926e-13, 1.142805e-13, 1.148107e-13, 1.151352e-13, 1.154652e-13, 
    1.156108e-13, 1.15655e-13, 1.156735e-13 ;

 LITR2C_vr =
  0.001150941, 0.00115094, 0.00115094, 0.001150939, 0.00115094, 0.001150939, 
    0.001150941, 0.00115094, 0.001150941, 0.001150941, 0.001150937, 
    0.001150939, 0.001150935, 0.001150937, 0.001150934, 0.001150936, 
    0.001150933, 0.001150934, 0.001150932, 0.001150933, 0.001150931, 
    0.001150932, 0.00115093, 0.001150931, 0.001150931, 0.001150932, 
    0.001150939, 0.001150938, 0.001150939, 0.001150939, 0.001150939, 
    0.00115094, 0.00115094, 0.001150941, 0.001150941, 0.00115094, 
    0.001150939, 0.001150939, 0.001150938, 0.001150938, 0.001150936, 
    0.001150937, 0.001150934, 0.001150935, 0.001150933, 0.001150933, 
    0.001150933, 0.001150933, 0.001150933, 0.001150934, 0.001150933, 
    0.001150934, 0.001150937, 0.001150936, 0.001150938, 0.00115094, 
    0.001150941, 0.001150941, 0.001150941, 0.001150941, 0.00115094, 
    0.001150939, 0.001150939, 0.001150938, 0.001150938, 0.001150936, 
    0.001150936, 0.001150934, 0.001150934, 0.001150934, 0.001150933, 
    0.001150933, 0.001150933, 0.001150932, 0.001150934, 0.001150933, 
    0.001150934, 0.001150934, 0.001150938, 0.001150939, 0.00115094, 
    0.00115094, 0.001150941, 0.00115094, 0.001150941, 0.00115094, 
    0.001150939, 0.00115094, 0.001150938, 0.001150939, 0.001150936, 
    0.001150937, 0.001150933, 0.001150934, 0.001150933, 0.001150934, 
    0.001150933, 0.001150934, 0.001150932, 0.001150932, 0.001150932, 
    0.001150931, 0.001150934, 0.001150933, 0.00115094, 0.00115094, 
    0.001150939, 0.00115094, 0.00115094, 0.001150941, 0.001150941, 
    0.00115094, 0.001150939, 0.001150939, 0.001150939, 0.001150938, 
    0.001150937, 0.001150935, 0.001150934, 0.001150933, 0.001150934, 
    0.001150934, 0.001150934, 0.001150934, 0.001150932, 0.001150933, 
    0.001150931, 0.001150931, 0.001150932, 0.001150931, 0.00115094, 
    0.00115094, 0.001150941, 0.00115094, 0.001150941, 0.001150941, 
    0.00115094, 0.001150939, 0.001150938, 0.001150938, 0.001150938, 
    0.001150937, 0.001150935, 0.001150934, 0.001150933, 0.001150933, 
    0.001150933, 0.001150933, 0.001150934, 0.001150933, 0.001150933, 
    0.001150933, 0.001150931, 0.001150932, 0.001150931, 0.001150932, 
    0.00115094, 0.001150939, 0.00115094, 0.001150939, 0.001150939, 
    0.001150938, 0.001150938, 0.001150936, 0.001150937, 0.001150936, 
    0.001150937, 0.001150936, 0.001150936, 0.001150937, 0.001150934, 
    0.001150936, 0.001150933, 0.001150935, 0.001150933, 0.001150933, 
    0.001150933, 0.001150932, 0.001150932, 0.001150931, 0.001150931, 
    0.00115093, 0.001150939, 0.001150938, 0.001150938, 0.001150938, 
    0.001150937, 0.001150937, 0.001150935, 0.001150936, 0.001150935, 
    0.001150934, 0.001150936, 0.001150935, 0.001150938, 0.001150938, 
    0.001150938, 0.001150939, 0.001150936, 0.001150937, 0.001150934, 
    0.001150935, 0.001150932, 0.001150934, 0.001150931, 0.00115093, 
    0.001150929, 0.001150928, 0.001150938, 0.001150938, 0.001150938, 
    0.001150937, 0.001150936, 0.001150935, 0.001150935, 0.001150935, 
    0.001150934, 0.001150934, 0.001150935, 0.001150934, 0.001150937, 
    0.001150935, 0.001150939, 0.001150938, 0.001150937, 0.001150937, 
    0.001150936, 0.001150935, 0.001150934, 0.001150935, 0.00115093, 
    0.001150932, 0.001150927, 0.001150928, 0.001150939, 0.001150938, 
    0.001150936, 0.001150937, 0.001150935, 0.001150934, 0.001150934, 
    0.001150933, 0.001150933, 0.001150933, 0.001150933, 0.001150933, 
    0.001150935, 0.001150934, 0.001150937, 0.001150936, 0.001150936, 
    0.001150937, 0.001150936, 0.001150935, 0.001150935, 0.001150934, 
    0.001150933, 0.001150935, 0.00115093, 0.001150933, 0.001150938, 
    0.001150937, 0.001150936, 0.001150937, 0.001150934, 0.001150935, 
    0.001150933, 0.001150934, 0.001150933, 0.001150933, 0.001150933, 
    0.001150934, 0.001150934, 0.001150935, 0.001150936, 0.001150937, 
    0.001150937, 0.001150936, 0.001150934, 0.001150933, 0.001150934, 
    0.001150933, 0.001150935, 0.001150934, 0.001150934, 0.001150933, 
    0.001150936, 0.001150934, 0.001150936, 0.001150936, 0.001150935, 
    0.001150934, 0.001150934, 0.001150933, 0.001150934, 0.001150934, 
    0.001150935, 0.001150935, 0.001150936, 0.001150936, 0.001150936, 
    0.001150936, 0.001150936, 0.001150934, 0.001150933, 0.001150932, 
    0.001150932, 0.001150931, 0.001150932, 0.00115093, 0.001150932, 
    0.001150929, 0.001150934, 0.001150932, 0.001150935, 0.001150935, 
    0.001150934, 0.001150933, 0.001150933, 0.001150932, 0.001150935, 
    0.001150936, 0.001150936, 0.001150937, 0.001150936, 0.001150936, 
    0.001150936, 0.001150936, 0.001150934, 0.001150935, 0.001150933, 
    0.001150932, 0.00115093, 0.001150929, 0.001150928, 0.001150927, 
    0.001150927, 0.001150927,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.789473e-07, 2.78947e-07, 2.789471e-07, 2.789468e-07, 2.789469e-07, 
    2.789468e-07, 2.789472e-07, 2.78947e-07, 2.789471e-07, 2.789473e-07, 
    2.789463e-07, 2.789468e-07, 2.789459e-07, 2.789462e-07, 2.789455e-07, 
    2.789459e-07, 2.789454e-07, 2.789455e-07, 2.789452e-07, 2.789452e-07, 
    2.789448e-07, 2.789451e-07, 2.789446e-07, 2.789449e-07, 2.789448e-07, 
    2.789451e-07, 2.789467e-07, 2.789464e-07, 2.789467e-07, 2.789467e-07, 
    2.789467e-07, 2.789469e-07, 2.789471e-07, 2.789473e-07, 2.789473e-07, 
    2.789471e-07, 2.789467e-07, 2.789468e-07, 2.789465e-07, 2.789465e-07, 
    2.789461e-07, 2.789463e-07, 2.789456e-07, 2.789458e-07, 2.789452e-07, 
    2.789454e-07, 2.789452e-07, 2.789453e-07, 2.789452e-07, 2.789454e-07, 
    2.789454e-07, 2.789455e-07, 2.789462e-07, 2.78946e-07, 2.789466e-07, 
    2.78947e-07, 2.789472e-07, 2.789474e-07, 2.789474e-07, 2.789473e-07, 
    2.789471e-07, 2.789469e-07, 2.789467e-07, 2.789466e-07, 2.789465e-07, 
    2.789461e-07, 2.789459e-07, 2.789455e-07, 2.789456e-07, 2.789455e-07, 
    2.789454e-07, 2.789452e-07, 2.789452e-07, 2.789452e-07, 2.789455e-07, 
    2.789453e-07, 2.789457e-07, 2.789455e-07, 2.789464e-07, 2.789468e-07, 
    2.789469e-07, 2.78947e-07, 2.789473e-07, 2.789471e-07, 2.789472e-07, 
    2.78947e-07, 2.789469e-07, 2.789469e-07, 2.789466e-07, 2.789467e-07, 
    2.789459e-07, 2.789463e-07, 2.789454e-07, 2.789456e-07, 2.789454e-07, 
    2.789455e-07, 2.789453e-07, 2.789455e-07, 2.789451e-07, 2.78945e-07, 
    2.789451e-07, 2.789449e-07, 2.789455e-07, 2.789452e-07, 2.789469e-07, 
    2.789469e-07, 2.789469e-07, 2.789471e-07, 2.789471e-07, 2.789473e-07, 
    2.789471e-07, 2.789471e-07, 2.789469e-07, 2.789468e-07, 2.789467e-07, 
    2.789465e-07, 2.789462e-07, 2.789459e-07, 2.789456e-07, 2.789454e-07, 
    2.789455e-07, 2.789454e-07, 2.789455e-07, 2.789456e-07, 2.789451e-07, 
    2.789454e-07, 2.789449e-07, 2.789449e-07, 2.789452e-07, 2.789449e-07, 
    2.789469e-07, 2.78947e-07, 2.789472e-07, 2.78947e-07, 2.789473e-07, 
    2.789472e-07, 2.789471e-07, 2.789467e-07, 2.789466e-07, 2.789466e-07, 
    2.789464e-07, 2.789462e-07, 2.789459e-07, 2.789456e-07, 2.789454e-07, 
    2.789454e-07, 2.789454e-07, 2.789454e-07, 2.789455e-07, 2.789453e-07, 
    2.789453e-07, 2.789454e-07, 2.78945e-07, 2.789451e-07, 2.789449e-07, 
    2.78945e-07, 2.78947e-07, 2.789469e-07, 2.789469e-07, 2.789468e-07, 
    2.789469e-07, 2.789466e-07, 2.789465e-07, 2.789461e-07, 2.789462e-07, 
    2.789459e-07, 2.789462e-07, 2.789462e-07, 2.789459e-07, 2.789462e-07, 
    2.789457e-07, 2.78946e-07, 2.789453e-07, 2.789457e-07, 2.789453e-07, 
    2.789454e-07, 2.789453e-07, 2.789452e-07, 2.78945e-07, 2.789448e-07, 
    2.789448e-07, 2.789446e-07, 2.789467e-07, 2.789466e-07, 2.789466e-07, 
    2.789465e-07, 2.789464e-07, 2.789462e-07, 2.789458e-07, 2.78946e-07, 
    2.789457e-07, 2.789457e-07, 2.78946e-07, 2.789458e-07, 2.789465e-07, 
    2.789464e-07, 2.789465e-07, 2.789467e-07, 2.789459e-07, 2.789463e-07, 
    2.789456e-07, 2.789458e-07, 2.789452e-07, 2.789455e-07, 2.789449e-07, 
    2.789446e-07, 2.789444e-07, 2.789441e-07, 2.789465e-07, 2.789466e-07, 
    2.789465e-07, 2.789463e-07, 2.789461e-07, 2.789458e-07, 2.789458e-07, 
    2.789457e-07, 2.789456e-07, 2.789455e-07, 2.789457e-07, 2.789455e-07, 
    2.789464e-07, 2.789459e-07, 2.789467e-07, 2.789464e-07, 2.789463e-07, 
    2.789463e-07, 2.78946e-07, 2.789459e-07, 2.789455e-07, 2.789457e-07, 
    2.789447e-07, 2.789452e-07, 2.789438e-07, 2.789442e-07, 2.789467e-07, 
    2.789465e-07, 2.789461e-07, 2.789463e-07, 2.789458e-07, 2.789456e-07, 
    2.789455e-07, 2.789454e-07, 2.789454e-07, 2.789453e-07, 2.789454e-07, 
    2.789453e-07, 2.789458e-07, 2.789456e-07, 2.789462e-07, 2.78946e-07, 
    2.789461e-07, 2.789462e-07, 2.789459e-07, 2.789457e-07, 2.789457e-07, 
    2.789456e-07, 2.789454e-07, 2.789458e-07, 2.789446e-07, 2.789453e-07, 
    2.789464e-07, 2.789462e-07, 2.789461e-07, 2.789462e-07, 2.789457e-07, 
    2.789459e-07, 2.789453e-07, 2.789455e-07, 2.789452e-07, 2.789453e-07, 
    2.789454e-07, 2.789455e-07, 2.789456e-07, 2.789459e-07, 2.789461e-07, 
    2.789462e-07, 2.789462e-07, 2.78946e-07, 2.789457e-07, 2.789454e-07, 
    2.789454e-07, 2.789452e-07, 2.789458e-07, 2.789456e-07, 2.789457e-07, 
    2.789454e-07, 2.78946e-07, 2.789455e-07, 2.789461e-07, 2.78946e-07, 
    2.789459e-07, 2.789455e-07, 2.789455e-07, 2.789454e-07, 2.789455e-07, 
    2.789457e-07, 2.789457e-07, 2.789459e-07, 2.789459e-07, 2.789461e-07, 
    2.789461e-07, 2.789461e-07, 2.789459e-07, 2.789457e-07, 2.789454e-07, 
    2.789452e-07, 2.789451e-07, 2.789448e-07, 2.78945e-07, 2.789446e-07, 
    2.78945e-07, 2.789443e-07, 2.789455e-07, 2.78945e-07, 2.789459e-07, 
    2.789458e-07, 2.789456e-07, 2.789452e-07, 2.789454e-07, 2.789452e-07, 
    2.789457e-07, 2.78946e-07, 2.789461e-07, 2.789462e-07, 2.789461e-07, 
    2.789461e-07, 2.789459e-07, 2.78946e-07, 2.789457e-07, 2.789458e-07, 
    2.789454e-07, 2.789452e-07, 2.789447e-07, 2.789444e-07, 2.78944e-07, 
    2.789439e-07, 2.789438e-07, 2.789438e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  5.637083e-26, 1.053889e-25, 3.161668e-25, -1.004871e-25, 1.347998e-25, 
    9.803622e-26, -2.181306e-25, -2.475414e-25, -1.715634e-25, -6.617445e-26, 
    1.666616e-25, 1.715634e-26, -2.450905e-26, 8.087988e-26, 2.279342e-25, 
    2.450906e-27, 3.921449e-26, 3.186177e-26, 1.004871e-25, -4.166539e-26, 
    -1.176435e-25, -1.470543e-26, 7.352717e-26, -1.347998e-25, 7.107626e-26, 
    4.166539e-26, -2.695996e-26, 1.740143e-25, -8.087988e-26, 2.058761e-25, 
    -1.249962e-25, 1.249962e-25, 1.274471e-25, 6.127264e-26, 9.558531e-26, 
    -4.65672e-26, 7.352717e-26, 4.901811e-26, 3.431268e-25, 1.127417e-25, 
    1.470543e-26, -9.068351e-26, 8.333079e-26, 1.200944e-25, 4.901811e-26, 
    -1.715634e-25, -1.56858e-25, -1.470543e-25, 3.186177e-26, 7.352717e-26, 
    2.156797e-25, -2.499924e-25, -8.82326e-26, 1.715634e-26, -5.391992e-26, 
    -8.578169e-26, 1.29898e-25, 1.127417e-25, -9.068351e-26, -3.921449e-26, 
    9.068351e-26, 7.352717e-26, -3.186177e-26, 2.695996e-26, 6.617445e-26, 
    2.034252e-25, 2.205815e-26, 1.225453e-25, -3.186177e-26, 2.965596e-25, 
    1.960724e-26, -2.990105e-25, 4.901811e-26, -6.372354e-26, -2.941087e-26, 
    -4.901811e-26, -3.431268e-26, -2.499924e-25, 1.715634e-25, -1.666616e-25, 
    4.901811e-27, 1.004871e-25, 2.499924e-25, 1.81367e-25, 9.803622e-26, 
    -5.146902e-26, -1.470543e-26, 4.65672e-26, 7.352717e-27, 3.186177e-26, 
    1.225453e-26, 1.911706e-25, 2.769523e-25, -1.642107e-25, -6.372354e-26, 
    8.333079e-26, -2.695996e-26, 9.068351e-26, 9.803622e-27, 1.617598e-25, 
    -1.56858e-25, 5.882173e-26, 2.450905e-26, -7.352717e-26, -1.274471e-25, 
    -3.921449e-26, 7.597807e-26, -1.004871e-25, 2.892069e-25, 3.921449e-26, 
    5.882173e-26, -3.431268e-26, 1.225453e-26, -6.862535e-26, 3.039123e-25, 
    1.176435e-25, -6.617445e-26, 1.666616e-25, -4.166539e-26, 2.646978e-25, 
    -1.004871e-25, -7.352717e-26, -1.960724e-26, -4.901811e-26, 
    -3.676358e-26, -1.470543e-26, 2.450906e-27, -7.352717e-27, -3.38225e-25, 
    4.41163e-26, 7.842898e-26, 1.397016e-25, 2.450906e-27, 2.377378e-25, 
    5.637083e-26, -2.034252e-25, 1.530638e-41, -8.578169e-26, -1.985233e-25, 
    -2.034252e-25, 1.911706e-25, 1.225453e-25, 1.004871e-25, -2.622469e-25, 
    2.450905e-26, -1.715634e-25, 6.127264e-26, -3.431268e-26, -2.450905e-26, 
    9.558531e-26, 2.941087e-26, -1.960724e-26, -1.715634e-25, 7.352717e-27, 
    1.666616e-25, 1.004871e-25, 1.666616e-25, -1.936215e-25, 1.593089e-25, 
    1.127417e-25, -2.622469e-25, 5.146902e-26, 1.666616e-25, 7.352717e-26, 
    -6.372354e-26, 7.352717e-26, -4.65672e-26, 3.921449e-26, 2.058761e-25, 
    -3.431268e-26, -1.02938e-25, 8.087988e-26, -2.254833e-25, -1.81367e-25, 
    1.81367e-25, -1.151926e-25, -1.004871e-25, -4.901811e-27, -7.352717e-27, 
    -2.941087e-26, -3.431268e-26, 5.146902e-26, 9.803622e-26, 1.176435e-25, 
    2.450905e-26, -1.56858e-25, -2.205815e-26, -2.132288e-25, 1.887197e-25, 
    -3.676358e-26, 2.450905e-26, -2.156797e-25, -1.470543e-26, -4.901811e-26, 
    1.593089e-25, 1.495052e-25, -1.862688e-25, -7.352717e-26, -4.41163e-26, 
    1.56858e-25, 1.078398e-25, 1.347998e-25, -9.803622e-26, 1.81367e-25, 
    -2.990105e-25, 9.803622e-27, -5.882173e-26, 2.695996e-26, 1.127417e-25, 
    -1.249962e-25, -4.901811e-26, 2.450905e-26, 6.127264e-26, -7.352717e-27, 
    6.862535e-26, 1.985233e-25, -1.936215e-25, 1.249962e-25, 8.333079e-26, 
    5.637083e-26, 1.960724e-26, -9.313441e-26, -1.274471e-25, 8.82326e-26, 
    -3.676358e-26, -4.166539e-26, -9.313441e-26, 1.54407e-25, 1.078398e-25, 
    -4.901811e-27, 3.284213e-25, -3.284213e-25, 2.034252e-25, -1.470543e-25, 
    1.102908e-25, 1.715634e-26, 2.769523e-25, 0, -1.274471e-25, 
    -1.960724e-26, -2.499924e-25, -1.764652e-25, 1.446034e-25, 1.715634e-26, 
    3.431268e-26, -1.495052e-25, 6.127264e-26, -1.470543e-26, 1.176435e-25, 
    7.352717e-26, -6.372354e-26, -1.862688e-25, 5.637083e-26, -7.597807e-26, 
    -5.637083e-26, -1.960724e-25, -1.960724e-26, 8.82326e-26, -5.146902e-26, 
    -1.740143e-25, -1.691125e-25, -2.695996e-26, -4.65672e-26, 1.691125e-25, 
    -1.446034e-25, -1.078398e-25, -8.578169e-26, 4.166539e-26, 1.151926e-25, 
    -1.053889e-25, 1.81367e-25, -4.166539e-26, 5.391992e-26, -1.397016e-25, 
    2.450906e-27, -5.146902e-26, -8.087988e-26, 1.151926e-25, -4.901811e-26, 
    -9.803622e-27, 9.803622e-26, -1.81367e-25, -2.009742e-25, 1.102908e-25, 
    9.803622e-27, 7.352717e-27, 1.200944e-25, 4.65672e-26, -3.431268e-26, 
    1.347998e-25, 1.176435e-25, -3.749886e-25, 2.695996e-25, -1.691125e-25, 
    8.82326e-26, -4.65672e-26, 9.558531e-26, -1.053889e-25, 4.65672e-26, 
    4.166539e-26, 6.862535e-26, 4.41163e-26, 3.921449e-26, -1.225453e-26, 
    -1.470543e-26, -1.470543e-25, 4.901811e-26, -7.352717e-26, 1.274471e-25, 
    -9.313441e-26, -5.391992e-26, 1.372507e-25, -8.333079e-26, 8.578169e-26, 
    2.941087e-26, 2.450906e-27, 8.087988e-26, -1.519561e-25, -5.882173e-26, 
    -1.642107e-25, -2.205815e-26, -2.32836e-25, 1.642107e-25, 8.578169e-26, 
    3.431268e-26, -2.695996e-26, 1.323489e-25, -9.313441e-26, -6.617445e-26, 
    -9.068351e-26, -2.058761e-25, 5.146902e-26, -1.225453e-25, 2.132288e-25, 
    -1.02938e-25, 9.803622e-27, -2.401887e-25, 3.11265e-25,
  2.781948e-32, 2.781945e-32, 2.781945e-32, 2.781943e-32, 2.781944e-32, 
    2.781943e-32, 2.781947e-32, 2.781945e-32, 2.781946e-32, 2.781947e-32, 
    2.781938e-32, 2.781943e-32, 2.781934e-32, 2.781936e-32, 2.781929e-32, 
    2.781934e-32, 2.781928e-32, 2.78193e-32, 2.781926e-32, 2.781927e-32, 
    2.781923e-32, 2.781926e-32, 2.781921e-32, 2.781924e-32, 2.781923e-32, 
    2.781926e-32, 2.781942e-32, 2.781939e-32, 2.781942e-32, 2.781942e-32, 
    2.781942e-32, 2.781944e-32, 2.781946e-32, 2.781948e-32, 2.781948e-32, 
    2.781946e-32, 2.781941e-32, 2.781943e-32, 2.781939e-32, 2.781939e-32, 
    2.781936e-32, 2.781937e-32, 2.781931e-32, 2.781933e-32, 2.781927e-32, 
    2.781928e-32, 2.781927e-32, 2.781928e-32, 2.781927e-32, 2.781929e-32, 
    2.781928e-32, 2.78193e-32, 2.781937e-32, 2.781935e-32, 2.781941e-32, 
    2.781945e-32, 2.781947e-32, 2.781949e-32, 2.781948e-32, 2.781948e-32, 
    2.781946e-32, 2.781943e-32, 2.781942e-32, 2.781941e-32, 2.781939e-32, 
    2.781936e-32, 2.781934e-32, 2.78193e-32, 2.781931e-32, 2.78193e-32, 
    2.781929e-32, 2.781927e-32, 2.781927e-32, 2.781926e-32, 2.78193e-32, 
    2.781927e-32, 2.781931e-32, 2.78193e-32, 2.781939e-32, 2.781943e-32, 
    2.781944e-32, 2.781945e-32, 2.781948e-32, 2.781946e-32, 2.781947e-32, 
    2.781945e-32, 2.781944e-32, 2.781944e-32, 2.781941e-32, 2.781942e-32, 
    2.781934e-32, 2.781938e-32, 2.781929e-32, 2.781931e-32, 2.781928e-32, 
    2.78193e-32, 2.781927e-32, 2.781929e-32, 2.781926e-32, 2.781925e-32, 
    2.781926e-32, 2.781923e-32, 2.781929e-32, 2.781927e-32, 2.781944e-32, 
    2.781944e-32, 2.781944e-32, 2.781946e-32, 2.781946e-32, 2.781948e-32, 
    2.781946e-32, 2.781946e-32, 2.781944e-32, 2.781943e-32, 2.781941e-32, 
    2.781939e-32, 2.781937e-32, 2.781933e-32, 2.781931e-32, 2.781929e-32, 
    2.78193e-32, 2.781929e-32, 2.78193e-32, 2.781931e-32, 2.781925e-32, 
    2.781928e-32, 2.781924e-32, 2.781924e-32, 2.781926e-32, 2.781924e-32, 
    2.781944e-32, 2.781945e-32, 2.781947e-32, 2.781945e-32, 2.781948e-32, 
    2.781946e-32, 2.781946e-32, 2.781942e-32, 2.781941e-32, 2.781941e-32, 
    2.781939e-32, 2.781937e-32, 2.781934e-32, 2.781931e-32, 2.781928e-32, 
    2.781929e-32, 2.781929e-32, 2.781928e-32, 2.78193e-32, 2.781928e-32, 
    2.781928e-32, 2.781928e-32, 2.781924e-32, 2.781925e-32, 2.781924e-32, 
    2.781925e-32, 2.781945e-32, 2.781943e-32, 2.781944e-32, 2.781943e-32, 
    2.781944e-32, 2.781941e-32, 2.78194e-32, 2.781936e-32, 2.781937e-32, 
    2.781934e-32, 2.781937e-32, 2.781936e-32, 2.781934e-32, 2.781937e-32, 
    2.781931e-32, 2.781935e-32, 2.781928e-32, 2.781932e-32, 2.781928e-32, 
    2.781928e-32, 2.781927e-32, 2.781926e-32, 2.781925e-32, 2.781923e-32, 
    2.781923e-32, 2.781921e-32, 2.781942e-32, 2.781941e-32, 2.781941e-32, 
    2.78194e-32, 2.781939e-32, 2.781936e-32, 2.781933e-32, 2.781934e-32, 
    2.781932e-32, 2.781932e-32, 2.781935e-32, 2.781933e-32, 2.78194e-32, 
    2.781939e-32, 2.78194e-32, 2.781942e-32, 2.781934e-32, 2.781938e-32, 
    2.781931e-32, 2.781933e-32, 2.781926e-32, 2.78193e-32, 2.781923e-32, 
    2.781921e-32, 2.781918e-32, 2.781915e-32, 2.78194e-32, 2.781941e-32, 
    2.78194e-32, 2.781937e-32, 2.781936e-32, 2.781933e-32, 2.781933e-32, 
    2.781932e-32, 2.781931e-32, 2.78193e-32, 2.781932e-32, 2.781929e-32, 
    2.781939e-32, 2.781934e-32, 2.781941e-32, 2.781939e-32, 2.781938e-32, 
    2.781938e-32, 2.781935e-32, 2.781934e-32, 2.78193e-32, 2.781932e-32, 
    2.781921e-32, 2.781926e-32, 2.781913e-32, 2.781917e-32, 2.781941e-32, 
    2.78194e-32, 2.781936e-32, 2.781938e-32, 2.781933e-32, 2.781931e-32, 
    2.78193e-32, 2.781929e-32, 2.781928e-32, 2.781928e-32, 2.781929e-32, 
    2.781928e-32, 2.781933e-32, 2.781931e-32, 2.781937e-32, 2.781935e-32, 
    2.781936e-32, 2.781937e-32, 2.781934e-32, 2.781932e-32, 2.781932e-32, 
    2.781931e-32, 2.781929e-32, 2.781933e-32, 2.781921e-32, 2.781928e-32, 
    2.781939e-32, 2.781937e-32, 2.781936e-32, 2.781937e-32, 2.781931e-32, 
    2.781933e-32, 2.781928e-32, 2.781929e-32, 2.781927e-32, 2.781928e-32, 
    2.781928e-32, 2.78193e-32, 2.781931e-32, 2.781933e-32, 2.781936e-32, 
    2.781937e-32, 2.781937e-32, 2.781935e-32, 2.781932e-32, 2.781928e-32, 
    2.781929e-32, 2.781927e-32, 2.781933e-32, 2.781931e-32, 2.781931e-32, 
    2.781929e-32, 2.781934e-32, 2.78193e-32, 2.781936e-32, 2.781935e-32, 
    2.781933e-32, 2.78193e-32, 2.78193e-32, 2.781929e-32, 2.781929e-32, 
    2.781932e-32, 2.781932e-32, 2.781933e-32, 2.781934e-32, 2.781935e-32, 
    2.781936e-32, 2.781935e-32, 2.781934e-32, 2.781932e-32, 2.781929e-32, 
    2.781926e-32, 2.781926e-32, 2.781923e-32, 2.781925e-32, 2.781921e-32, 
    2.781924e-32, 2.781918e-32, 2.781929e-32, 2.781925e-32, 2.781933e-32, 
    2.781933e-32, 2.781931e-32, 2.781927e-32, 2.781929e-32, 2.781926e-32, 
    2.781932e-32, 2.781935e-32, 2.781936e-32, 2.781937e-32, 2.781936e-32, 
    2.781936e-32, 2.781934e-32, 2.781935e-32, 2.781931e-32, 2.781933e-32, 
    2.781928e-32, 2.781926e-32, 2.781921e-32, 2.781918e-32, 2.781915e-32, 
    2.781913e-32, 2.781913e-32, 2.781913e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.102539e-15, 3.110906e-15, 3.10928e-15, 3.116022e-15, 3.112284e-15, 
    3.116697e-15, 3.104237e-15, 3.111237e-15, 3.10677e-15, 3.103294e-15, 
    3.129087e-15, 3.116323e-15, 3.142333e-15, 3.134207e-15, 3.154604e-15, 
    3.141067e-15, 3.157332e-15, 3.154216e-15, 3.163595e-15, 3.160909e-15, 
    3.172887e-15, 3.164834e-15, 3.179092e-15, 3.170966e-15, 3.172237e-15, 
    3.164568e-15, 3.118896e-15, 3.127498e-15, 3.118385e-15, 3.119613e-15, 
    3.119063e-15, 3.112361e-15, 3.108979e-15, 3.101901e-15, 3.103187e-15, 
    3.108387e-15, 3.120165e-15, 3.11617e-15, 3.126239e-15, 3.126012e-15, 
    3.137204e-15, 3.132159e-15, 3.150947e-15, 3.145614e-15, 3.161022e-15, 
    3.157149e-15, 3.160839e-15, 3.159721e-15, 3.160854e-15, 3.155173e-15, 
    3.157608e-15, 3.152608e-15, 3.133104e-15, 3.138841e-15, 3.121717e-15, 
    3.111399e-15, 3.104544e-15, 3.099675e-15, 3.100363e-15, 3.101675e-15, 
    3.108417e-15, 3.114753e-15, 3.119577e-15, 3.122802e-15, 3.125979e-15, 
    3.13558e-15, 3.140662e-15, 3.152025e-15, 3.149977e-15, 3.153447e-15, 
    3.156763e-15, 3.162326e-15, 3.161411e-15, 3.16386e-15, 3.153357e-15, 
    3.160338e-15, 3.14881e-15, 3.151965e-15, 3.126834e-15, 3.117248e-15, 
    3.113164e-15, 3.109593e-15, 3.100892e-15, 3.106901e-15, 3.104533e-15, 
    3.110168e-15, 3.113745e-15, 3.111977e-15, 3.12289e-15, 3.118649e-15, 
    3.140963e-15, 3.13136e-15, 3.156377e-15, 3.150398e-15, 3.15781e-15, 
    3.154029e-15, 3.160505e-15, 3.154677e-15, 3.164772e-15, 3.166967e-15, 
    3.165467e-15, 3.171231e-15, 3.154353e-15, 3.160838e-15, 3.111927e-15, 
    3.112215e-15, 3.11356e-15, 3.107647e-15, 3.107286e-15, 3.101866e-15, 
    3.106689e-15, 3.108742e-15, 3.113953e-15, 3.117033e-15, 3.11996e-15, 
    3.126391e-15, 3.133567e-15, 3.143591e-15, 3.150785e-15, 3.155604e-15, 
    3.15265e-15, 3.155258e-15, 3.152342e-15, 3.150976e-15, 3.166144e-15, 
    3.15763e-15, 3.170402e-15, 3.169697e-15, 3.163918e-15, 3.169776e-15, 
    3.112418e-15, 3.110758e-15, 3.104988e-15, 3.109503e-15, 3.101275e-15, 
    3.105881e-15, 3.108527e-15, 3.118736e-15, 3.120979e-15, 3.123055e-15, 
    3.127158e-15, 3.132417e-15, 3.141636e-15, 3.149648e-15, 3.156957e-15, 
    3.156422e-15, 3.15661e-15, 3.158241e-15, 3.154199e-15, 3.158905e-15, 
    3.159693e-15, 3.15763e-15, 3.169602e-15, 3.166184e-15, 3.169682e-15, 
    3.167456e-15, 3.111297e-15, 3.114091e-15, 3.112582e-15, 3.11542e-15, 
    3.11342e-15, 3.122307e-15, 3.124969e-15, 3.137418e-15, 3.132313e-15, 
    3.140438e-15, 3.13314e-15, 3.134433e-15, 3.140699e-15, 3.133535e-15, 
    3.149204e-15, 3.138582e-15, 3.158304e-15, 3.147706e-15, 3.158968e-15, 
    3.156925e-15, 3.160308e-15, 3.163336e-15, 3.167144e-15, 3.174164e-15, 
    3.17254e-15, 3.178408e-15, 3.118255e-15, 3.121875e-15, 3.121557e-15, 
    3.125345e-15, 3.128144e-15, 3.13421e-15, 3.143928e-15, 3.140276e-15, 
    3.146981e-15, 3.148324e-15, 3.138139e-15, 3.144394e-15, 3.124297e-15, 
    3.127546e-15, 3.125613e-15, 3.11854e-15, 3.141115e-15, 3.129536e-15, 
    3.150904e-15, 3.144643e-15, 3.162904e-15, 3.153825e-15, 3.171645e-15, 
    3.179245e-15, 3.186399e-15, 3.194742e-15, 3.123851e-15, 3.121392e-15, 
    3.125796e-15, 3.131881e-15, 3.137527e-15, 3.145025e-15, 3.145793e-15, 
    3.147196e-15, 3.15083e-15, 3.153884e-15, 3.147638e-15, 3.15465e-15, 
    3.128296e-15, 3.14212e-15, 3.120461e-15, 3.126987e-15, 3.131523e-15, 
    3.129535e-15, 3.139859e-15, 3.142289e-15, 3.152156e-15, 3.147059e-15, 
    3.177369e-15, 3.163973e-15, 3.201093e-15, 3.190737e-15, 3.120532e-15, 
    3.123843e-15, 3.135352e-15, 3.129879e-15, 3.145526e-15, 3.149371e-15, 
    3.152497e-15, 3.156489e-15, 3.156921e-15, 3.159286e-15, 3.155411e-15, 
    3.159134e-15, 3.145041e-15, 3.151341e-15, 3.134039e-15, 3.138254e-15, 
    3.136316e-15, 3.134189e-15, 3.140752e-15, 3.147734e-15, 3.147886e-15, 
    3.150124e-15, 3.156421e-15, 3.14559e-15, 3.179091e-15, 3.158413e-15, 
    3.127452e-15, 3.133818e-15, 3.13473e-15, 3.132264e-15, 3.148985e-15, 
    3.142931e-15, 3.159229e-15, 3.154828e-15, 3.162038e-15, 3.158456e-15, 
    3.157928e-15, 3.153325e-15, 3.150457e-15, 3.143209e-15, 3.137305e-15, 
    3.132622e-15, 3.133712e-15, 3.138855e-15, 3.148162e-15, 3.15696e-15, 
    3.155033e-15, 3.161491e-15, 3.144393e-15, 3.151564e-15, 3.148792e-15, 
    3.15602e-15, 3.140178e-15, 3.153662e-15, 3.136726e-15, 3.138213e-15, 
    3.142811e-15, 3.152049e-15, 3.154095e-15, 3.156275e-15, 3.154931e-15, 
    3.148399e-15, 3.147331e-15, 3.1427e-15, 3.14142e-15, 3.13789e-15, 
    3.134965e-15, 3.137637e-15, 3.140441e-15, 3.148402e-15, 3.15557e-15, 
    3.163378e-15, 3.165289e-15, 3.174393e-15, 3.166979e-15, 3.179205e-15, 
    3.168806e-15, 3.186801e-15, 3.154446e-15, 3.168506e-15, 3.143021e-15, 
    3.145772e-15, 3.150739e-15, 3.16213e-15, 3.155986e-15, 3.163173e-15, 
    3.147289e-15, 3.139031e-15, 3.136896e-15, 3.132907e-15, 3.136988e-15, 
    3.136656e-15, 3.140559e-15, 3.139305e-15, 3.148667e-15, 3.14364e-15, 
    3.157914e-15, 3.163117e-15, 3.177792e-15, 3.186773e-15, 3.195908e-15, 
    3.199936e-15, 3.201161e-15, 3.201674e-15 ;

 LITR2N_vr =
  1.592818e-05, 1.592816e-05, 1.592816e-05, 1.592815e-05, 1.592816e-05, 
    1.592815e-05, 1.592818e-05, 1.592816e-05, 1.592817e-05, 1.592818e-05, 
    1.592812e-05, 1.592815e-05, 1.59281e-05, 1.592812e-05, 1.592807e-05, 
    1.59281e-05, 1.592807e-05, 1.592808e-05, 1.592806e-05, 1.592806e-05, 
    1.592804e-05, 1.592805e-05, 1.592803e-05, 1.592804e-05, 1.592804e-05, 
    1.592806e-05, 1.592815e-05, 1.592813e-05, 1.592815e-05, 1.592814e-05, 
    1.592814e-05, 1.592816e-05, 1.592816e-05, 1.592818e-05, 1.592818e-05, 
    1.592817e-05, 1.592814e-05, 1.592815e-05, 1.592813e-05, 1.592813e-05, 
    1.592811e-05, 1.592812e-05, 1.592808e-05, 1.592809e-05, 1.592806e-05, 
    1.592807e-05, 1.592806e-05, 1.592806e-05, 1.592806e-05, 1.592807e-05, 
    1.592807e-05, 1.592808e-05, 1.592812e-05, 1.592811e-05, 1.592814e-05, 
    1.592816e-05, 1.592817e-05, 1.592818e-05, 1.592818e-05, 1.592818e-05, 
    1.592817e-05, 1.592815e-05, 1.592814e-05, 1.592814e-05, 1.592813e-05, 
    1.592811e-05, 1.59281e-05, 1.592808e-05, 1.592808e-05, 1.592808e-05, 
    1.592807e-05, 1.592806e-05, 1.592806e-05, 1.592806e-05, 1.592808e-05, 
    1.592806e-05, 1.592809e-05, 1.592808e-05, 1.592813e-05, 1.592815e-05, 
    1.592816e-05, 1.592816e-05, 1.592818e-05, 1.592817e-05, 1.592817e-05, 
    1.592816e-05, 1.592816e-05, 1.592816e-05, 1.592814e-05, 1.592815e-05, 
    1.59281e-05, 1.592812e-05, 1.592807e-05, 1.592808e-05, 1.592807e-05, 
    1.592808e-05, 1.592806e-05, 1.592807e-05, 1.592805e-05, 1.592805e-05, 
    1.592805e-05, 1.592804e-05, 1.592808e-05, 1.592806e-05, 1.592816e-05, 
    1.592816e-05, 1.592816e-05, 1.592817e-05, 1.592817e-05, 1.592818e-05, 
    1.592817e-05, 1.592817e-05, 1.592816e-05, 1.592815e-05, 1.592814e-05, 
    1.592813e-05, 1.592812e-05, 1.59281e-05, 1.592808e-05, 1.592807e-05, 
    1.592808e-05, 1.592807e-05, 1.592808e-05, 1.592808e-05, 1.592805e-05, 
    1.592807e-05, 1.592804e-05, 1.592804e-05, 1.592806e-05, 1.592804e-05, 
    1.592816e-05, 1.592816e-05, 1.592817e-05, 1.592816e-05, 1.592818e-05, 
    1.592817e-05, 1.592817e-05, 1.592815e-05, 1.592814e-05, 1.592814e-05, 
    1.592813e-05, 1.592812e-05, 1.59281e-05, 1.592808e-05, 1.592807e-05, 
    1.592807e-05, 1.592807e-05, 1.592807e-05, 1.592808e-05, 1.592807e-05, 
    1.592806e-05, 1.592807e-05, 1.592804e-05, 1.592805e-05, 1.592804e-05, 
    1.592805e-05, 1.592816e-05, 1.592816e-05, 1.592816e-05, 1.592815e-05, 
    1.592816e-05, 1.592814e-05, 1.592813e-05, 1.592811e-05, 1.592812e-05, 
    1.59281e-05, 1.592812e-05, 1.592812e-05, 1.59281e-05, 1.592812e-05, 
    1.592808e-05, 1.592811e-05, 1.592807e-05, 1.592809e-05, 1.592807e-05, 
    1.592807e-05, 1.592806e-05, 1.592806e-05, 1.592805e-05, 1.592804e-05, 
    1.592804e-05, 1.592803e-05, 1.592815e-05, 1.592814e-05, 1.592814e-05, 
    1.592813e-05, 1.592813e-05, 1.592812e-05, 1.59281e-05, 1.59281e-05, 
    1.592809e-05, 1.592809e-05, 1.592811e-05, 1.59281e-05, 1.592814e-05, 
    1.592813e-05, 1.592813e-05, 1.592815e-05, 1.59281e-05, 1.592812e-05, 
    1.592808e-05, 1.592809e-05, 1.592806e-05, 1.592808e-05, 1.592804e-05, 
    1.592802e-05, 1.592801e-05, 1.592799e-05, 1.592814e-05, 1.592814e-05, 
    1.592813e-05, 1.592812e-05, 1.592811e-05, 1.592809e-05, 1.592809e-05, 
    1.592809e-05, 1.592808e-05, 1.592808e-05, 1.592809e-05, 1.592807e-05, 
    1.592813e-05, 1.59281e-05, 1.592814e-05, 1.592813e-05, 1.592812e-05, 
    1.592812e-05, 1.59281e-05, 1.59281e-05, 1.592808e-05, 1.592809e-05, 
    1.592803e-05, 1.592806e-05, 1.592798e-05, 1.5928e-05, 1.592814e-05, 
    1.592814e-05, 1.592811e-05, 1.592812e-05, 1.592809e-05, 1.592808e-05, 
    1.592808e-05, 1.592807e-05, 1.592807e-05, 1.592806e-05, 1.592807e-05, 
    1.592806e-05, 1.592809e-05, 1.592808e-05, 1.592812e-05, 1.592811e-05, 
    1.592811e-05, 1.592812e-05, 1.59281e-05, 1.592809e-05, 1.592809e-05, 
    1.592808e-05, 1.592807e-05, 1.592809e-05, 1.592803e-05, 1.592807e-05, 
    1.592813e-05, 1.592812e-05, 1.592811e-05, 1.592812e-05, 1.592809e-05, 
    1.59281e-05, 1.592806e-05, 1.592807e-05, 1.592806e-05, 1.592807e-05, 
    1.592807e-05, 1.592808e-05, 1.592808e-05, 1.59281e-05, 1.592811e-05, 
    1.592812e-05, 1.592812e-05, 1.592811e-05, 1.592809e-05, 1.592807e-05, 
    1.592807e-05, 1.592806e-05, 1.59281e-05, 1.592808e-05, 1.592809e-05, 
    1.592807e-05, 1.59281e-05, 1.592808e-05, 1.592811e-05, 1.592811e-05, 
    1.59281e-05, 1.592808e-05, 1.592808e-05, 1.592807e-05, 1.592807e-05, 
    1.592809e-05, 1.592809e-05, 1.59281e-05, 1.59281e-05, 1.592811e-05, 
    1.592811e-05, 1.592811e-05, 1.59281e-05, 1.592809e-05, 1.592807e-05, 
    1.592806e-05, 1.592805e-05, 1.592804e-05, 1.592805e-05, 1.592802e-05, 
    1.592805e-05, 1.592801e-05, 1.592808e-05, 1.592805e-05, 1.59281e-05, 
    1.592809e-05, 1.592808e-05, 1.592806e-05, 1.592807e-05, 1.592806e-05, 
    1.592809e-05, 1.592811e-05, 1.592811e-05, 1.592812e-05, 1.592811e-05, 
    1.592811e-05, 1.59281e-05, 1.59281e-05, 1.592809e-05, 1.59281e-05, 
    1.592807e-05, 1.592806e-05, 1.592803e-05, 1.592801e-05, 1.592799e-05, 
    1.592798e-05, 1.592798e-05, 1.592798e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.120919e-13, 1.123942e-13, 1.123355e-13, 1.12579e-13, 1.12444e-13, 
    1.126034e-13, 1.121533e-13, 1.124061e-13, 1.122448e-13, 1.121192e-13, 
    1.13051e-13, 1.125899e-13, 1.135296e-13, 1.13236e-13, 1.13973e-13, 
    1.134839e-13, 1.140715e-13, 1.13959e-13, 1.142978e-13, 1.142008e-13, 
    1.146335e-13, 1.143426e-13, 1.148577e-13, 1.145641e-13, 1.1461e-13, 
    1.143329e-13, 1.126829e-13, 1.129936e-13, 1.126644e-13, 1.127088e-13, 
    1.126889e-13, 1.124467e-13, 1.123246e-13, 1.120689e-13, 1.121153e-13, 
    1.123032e-13, 1.127287e-13, 1.125844e-13, 1.129481e-13, 1.129399e-13, 
    1.133443e-13, 1.13162e-13, 1.138408e-13, 1.136482e-13, 1.142048e-13, 
    1.140649e-13, 1.141982e-13, 1.141578e-13, 1.141988e-13, 1.139935e-13, 
    1.140815e-13, 1.139008e-13, 1.131962e-13, 1.134034e-13, 1.127848e-13, 
    1.12412e-13, 1.121643e-13, 1.119884e-13, 1.120133e-13, 1.120607e-13, 
    1.123043e-13, 1.125332e-13, 1.127075e-13, 1.12824e-13, 1.129388e-13, 
    1.132856e-13, 1.134693e-13, 1.138798e-13, 1.138058e-13, 1.139312e-13, 
    1.14051e-13, 1.142519e-13, 1.142189e-13, 1.143074e-13, 1.139279e-13, 
    1.141801e-13, 1.137636e-13, 1.138776e-13, 1.129696e-13, 1.126233e-13, 
    1.124758e-13, 1.123467e-13, 1.120324e-13, 1.122495e-13, 1.121639e-13, 
    1.123675e-13, 1.124968e-13, 1.124329e-13, 1.128272e-13, 1.126739e-13, 
    1.134801e-13, 1.131332e-13, 1.14037e-13, 1.13821e-13, 1.140888e-13, 
    1.139522e-13, 1.141862e-13, 1.139756e-13, 1.143403e-13, 1.144196e-13, 
    1.143654e-13, 1.145737e-13, 1.139639e-13, 1.141982e-13, 1.124311e-13, 
    1.124415e-13, 1.124901e-13, 1.122764e-13, 1.122634e-13, 1.120676e-13, 
    1.122418e-13, 1.12316e-13, 1.125043e-13, 1.126156e-13, 1.127213e-13, 
    1.129537e-13, 1.132129e-13, 1.135751e-13, 1.13835e-13, 1.140091e-13, 
    1.139024e-13, 1.139966e-13, 1.138913e-13, 1.138419e-13, 1.143899e-13, 
    1.140823e-13, 1.145438e-13, 1.145182e-13, 1.143095e-13, 1.145211e-13, 
    1.124488e-13, 1.123888e-13, 1.121804e-13, 1.123435e-13, 1.120462e-13, 
    1.122126e-13, 1.123083e-13, 1.126771e-13, 1.127581e-13, 1.128331e-13, 
    1.129813e-13, 1.131714e-13, 1.135044e-13, 1.137939e-13, 1.14058e-13, 
    1.140386e-13, 1.140454e-13, 1.141044e-13, 1.139583e-13, 1.141283e-13, 
    1.141568e-13, 1.140823e-13, 1.145148e-13, 1.143913e-13, 1.145177e-13, 
    1.144373e-13, 1.124083e-13, 1.125093e-13, 1.124547e-13, 1.125573e-13, 
    1.12485e-13, 1.128061e-13, 1.129023e-13, 1.13352e-13, 1.131676e-13, 
    1.134612e-13, 1.131975e-13, 1.132442e-13, 1.134706e-13, 1.132118e-13, 
    1.137779e-13, 1.133941e-13, 1.141067e-13, 1.137237e-13, 1.141306e-13, 
    1.140568e-13, 1.14179e-13, 1.142884e-13, 1.14426e-13, 1.146797e-13, 
    1.14621e-13, 1.14833e-13, 1.126597e-13, 1.127905e-13, 1.12779e-13, 
    1.129159e-13, 1.13017e-13, 1.132362e-13, 1.135872e-13, 1.134553e-13, 
    1.136976e-13, 1.137461e-13, 1.133781e-13, 1.136041e-13, 1.12878e-13, 
    1.129954e-13, 1.129255e-13, 1.1267e-13, 1.134856e-13, 1.130673e-13, 
    1.138393e-13, 1.136131e-13, 1.142728e-13, 1.139448e-13, 1.145886e-13, 
    1.148632e-13, 1.151217e-13, 1.154231e-13, 1.128619e-13, 1.12773e-13, 
    1.129321e-13, 1.13152e-13, 1.13356e-13, 1.136269e-13, 1.136546e-13, 
    1.137053e-13, 1.138366e-13, 1.13947e-13, 1.137213e-13, 1.139746e-13, 
    1.130225e-13, 1.135219e-13, 1.127394e-13, 1.129752e-13, 1.131391e-13, 
    1.130673e-13, 1.134402e-13, 1.13528e-13, 1.138845e-13, 1.137003e-13, 
    1.147954e-13, 1.143114e-13, 1.156526e-13, 1.152784e-13, 1.12742e-13, 
    1.128616e-13, 1.132774e-13, 1.130797e-13, 1.13645e-13, 1.137839e-13, 
    1.138968e-13, 1.140411e-13, 1.140567e-13, 1.141421e-13, 1.140021e-13, 
    1.141366e-13, 1.136275e-13, 1.138551e-13, 1.1323e-13, 1.133822e-13, 
    1.133122e-13, 1.132354e-13, 1.134725e-13, 1.137248e-13, 1.137302e-13, 
    1.138111e-13, 1.140386e-13, 1.136473e-13, 1.148577e-13, 1.141106e-13, 
    1.12992e-13, 1.13222e-13, 1.132549e-13, 1.131658e-13, 1.1377e-13, 
    1.135512e-13, 1.1414e-13, 1.13981e-13, 1.142416e-13, 1.141121e-13, 
    1.140931e-13, 1.139268e-13, 1.138231e-13, 1.135613e-13, 1.13348e-13, 
    1.131788e-13, 1.132181e-13, 1.13404e-13, 1.137402e-13, 1.140581e-13, 
    1.139884e-13, 1.142218e-13, 1.13604e-13, 1.138631e-13, 1.13763e-13, 
    1.140241e-13, 1.134518e-13, 1.139389e-13, 1.133271e-13, 1.133808e-13, 
    1.135469e-13, 1.138807e-13, 1.139546e-13, 1.140333e-13, 1.139848e-13, 
    1.137488e-13, 1.137102e-13, 1.135429e-13, 1.134966e-13, 1.133691e-13, 
    1.132634e-13, 1.133599e-13, 1.134613e-13, 1.137489e-13, 1.140079e-13, 
    1.1429e-13, 1.14359e-13, 1.146879e-13, 1.144201e-13, 1.148618e-13, 
    1.144861e-13, 1.151362e-13, 1.139673e-13, 1.144752e-13, 1.135545e-13, 
    1.136539e-13, 1.138333e-13, 1.142449e-13, 1.140229e-13, 1.142826e-13, 
    1.137087e-13, 1.134103e-13, 1.133332e-13, 1.131891e-13, 1.133365e-13, 
    1.133245e-13, 1.134655e-13, 1.134202e-13, 1.137584e-13, 1.135769e-13, 
    1.140926e-13, 1.142805e-13, 1.148107e-13, 1.151352e-13, 1.154652e-13, 
    1.156108e-13, 1.15655e-13, 1.156735e-13 ;

 LITR3C =
  1.007811e-05, 1.00781e-05, 1.00781e-05, 1.007809e-05, 1.00781e-05, 
    1.007809e-05, 1.007811e-05, 1.00781e-05, 1.00781e-05, 1.007811e-05, 
    1.007807e-05, 1.007809e-05, 1.007806e-05, 1.007807e-05, 1.007804e-05, 
    1.007806e-05, 1.007804e-05, 1.007804e-05, 1.007803e-05, 1.007803e-05, 
    1.007802e-05, 1.007803e-05, 1.007801e-05, 1.007802e-05, 1.007802e-05, 
    1.007803e-05, 1.007809e-05, 1.007808e-05, 1.007809e-05, 1.007809e-05, 
    1.007809e-05, 1.00781e-05, 1.00781e-05, 1.007811e-05, 1.007811e-05, 
    1.00781e-05, 1.007809e-05, 1.007809e-05, 1.007808e-05, 1.007808e-05, 
    1.007806e-05, 1.007807e-05, 1.007805e-05, 1.007805e-05, 1.007803e-05, 
    1.007804e-05, 1.007803e-05, 1.007804e-05, 1.007803e-05, 1.007804e-05, 
    1.007804e-05, 1.007804e-05, 1.007807e-05, 1.007806e-05, 1.007808e-05, 
    1.00781e-05, 1.007811e-05, 1.007811e-05, 1.007811e-05, 1.007811e-05, 
    1.00781e-05, 1.007809e-05, 1.007809e-05, 1.007808e-05, 1.007808e-05, 
    1.007807e-05, 1.007806e-05, 1.007805e-05, 1.007805e-05, 1.007804e-05, 
    1.007804e-05, 1.007803e-05, 1.007803e-05, 1.007803e-05, 1.007804e-05, 
    1.007804e-05, 1.007805e-05, 1.007805e-05, 1.007808e-05, 1.007809e-05, 
    1.007809e-05, 1.00781e-05, 1.007811e-05, 1.00781e-05, 1.007811e-05, 
    1.00781e-05, 1.007809e-05, 1.00781e-05, 1.007808e-05, 1.007809e-05, 
    1.007806e-05, 1.007807e-05, 1.007804e-05, 1.007805e-05, 1.007804e-05, 
    1.007804e-05, 1.007803e-05, 1.007804e-05, 1.007803e-05, 1.007803e-05, 
    1.007803e-05, 1.007802e-05, 1.007804e-05, 1.007803e-05, 1.00781e-05, 
    1.00781e-05, 1.007809e-05, 1.00781e-05, 1.00781e-05, 1.007811e-05, 
    1.00781e-05, 1.00781e-05, 1.007809e-05, 1.007809e-05, 1.007809e-05, 
    1.007808e-05, 1.007807e-05, 1.007806e-05, 1.007805e-05, 1.007804e-05, 
    1.007804e-05, 1.007804e-05, 1.007805e-05, 1.007805e-05, 1.007803e-05, 
    1.007804e-05, 1.007802e-05, 1.007802e-05, 1.007803e-05, 1.007802e-05, 
    1.00781e-05, 1.00781e-05, 1.00781e-05, 1.00781e-05, 1.007811e-05, 
    1.00781e-05, 1.00781e-05, 1.007809e-05, 1.007808e-05, 1.007808e-05, 
    1.007808e-05, 1.007807e-05, 1.007806e-05, 1.007805e-05, 1.007804e-05, 
    1.007804e-05, 1.007804e-05, 1.007804e-05, 1.007804e-05, 1.007804e-05, 
    1.007804e-05, 1.007804e-05, 1.007802e-05, 1.007803e-05, 1.007802e-05, 
    1.007803e-05, 1.00781e-05, 1.007809e-05, 1.00781e-05, 1.007809e-05, 
    1.007809e-05, 1.007808e-05, 1.007808e-05, 1.007806e-05, 1.007807e-05, 
    1.007806e-05, 1.007807e-05, 1.007807e-05, 1.007806e-05, 1.007807e-05, 
    1.007805e-05, 1.007806e-05, 1.007804e-05, 1.007805e-05, 1.007804e-05, 
    1.007804e-05, 1.007804e-05, 1.007803e-05, 1.007803e-05, 1.007802e-05, 
    1.007802e-05, 1.007801e-05, 1.007809e-05, 1.007808e-05, 1.007808e-05, 
    1.007808e-05, 1.007808e-05, 1.007807e-05, 1.007806e-05, 1.007806e-05, 
    1.007805e-05, 1.007805e-05, 1.007806e-05, 1.007806e-05, 1.007808e-05, 
    1.007808e-05, 1.007808e-05, 1.007809e-05, 1.007806e-05, 1.007807e-05, 
    1.007805e-05, 1.007805e-05, 1.007803e-05, 1.007804e-05, 1.007802e-05, 
    1.007801e-05, 1.0078e-05, 1.007799e-05, 1.007808e-05, 1.007808e-05, 
    1.007808e-05, 1.007807e-05, 1.007806e-05, 1.007805e-05, 1.007805e-05, 
    1.007805e-05, 1.007805e-05, 1.007804e-05, 1.007805e-05, 1.007804e-05, 
    1.007808e-05, 1.007806e-05, 1.007809e-05, 1.007808e-05, 1.007807e-05, 
    1.007807e-05, 1.007806e-05, 1.007806e-05, 1.007805e-05, 1.007805e-05, 
    1.007801e-05, 1.007803e-05, 1.007798e-05, 1.0078e-05, 1.007809e-05, 
    1.007808e-05, 1.007807e-05, 1.007807e-05, 1.007805e-05, 1.007805e-05, 
    1.007805e-05, 1.007804e-05, 1.007804e-05, 1.007804e-05, 1.007804e-05, 
    1.007804e-05, 1.007805e-05, 1.007805e-05, 1.007807e-05, 1.007806e-05, 
    1.007807e-05, 1.007807e-05, 1.007806e-05, 1.007805e-05, 1.007805e-05, 
    1.007805e-05, 1.007804e-05, 1.007805e-05, 1.007801e-05, 1.007804e-05, 
    1.007808e-05, 1.007807e-05, 1.007807e-05, 1.007807e-05, 1.007805e-05, 
    1.007806e-05, 1.007804e-05, 1.007804e-05, 1.007803e-05, 1.007804e-05, 
    1.007804e-05, 1.007804e-05, 1.007805e-05, 1.007806e-05, 1.007806e-05, 
    1.007807e-05, 1.007807e-05, 1.007806e-05, 1.007805e-05, 1.007804e-05, 
    1.007804e-05, 1.007803e-05, 1.007806e-05, 1.007805e-05, 1.007805e-05, 
    1.007804e-05, 1.007806e-05, 1.007804e-05, 1.007806e-05, 1.007806e-05, 
    1.007806e-05, 1.007805e-05, 1.007804e-05, 1.007804e-05, 1.007804e-05, 
    1.007805e-05, 1.007805e-05, 1.007806e-05, 1.007806e-05, 1.007806e-05, 
    1.007807e-05, 1.007806e-05, 1.007806e-05, 1.007805e-05, 1.007804e-05, 
    1.007803e-05, 1.007803e-05, 1.007802e-05, 1.007803e-05, 1.007801e-05, 
    1.007802e-05, 1.0078e-05, 1.007804e-05, 1.007802e-05, 1.007806e-05, 
    1.007805e-05, 1.007805e-05, 1.007803e-05, 1.007804e-05, 1.007803e-05, 
    1.007805e-05, 1.007806e-05, 1.007806e-05, 1.007807e-05, 1.007806e-05, 
    1.007806e-05, 1.007806e-05, 1.007806e-05, 1.007805e-05, 1.007806e-05, 
    1.007804e-05, 1.007803e-05, 1.007801e-05, 1.0078e-05, 1.007799e-05, 
    1.007799e-05, 1.007798e-05, 1.007798e-05 ;

 LITR3C_TO_SOIL2C =
  5.604594e-14, 5.619708e-14, 5.616772e-14, 5.628951e-14, 5.622197e-14, 
    5.630169e-14, 5.607661e-14, 5.620306e-14, 5.612236e-14, 5.605958e-14, 
    5.65255e-14, 5.629494e-14, 5.676479e-14, 5.6618e-14, 5.698647e-14, 
    5.674193e-14, 5.703574e-14, 5.697947e-14, 5.714888e-14, 5.710037e-14, 
    5.731673e-14, 5.717126e-14, 5.742883e-14, 5.728203e-14, 5.730499e-14, 
    5.716645e-14, 5.634141e-14, 5.649681e-14, 5.633219e-14, 5.635437e-14, 
    5.634442e-14, 5.622336e-14, 5.616228e-14, 5.603441e-14, 5.605764e-14, 
    5.615157e-14, 5.636433e-14, 5.629217e-14, 5.647405e-14, 5.646995e-14, 
    5.667214e-14, 5.658101e-14, 5.692041e-14, 5.682406e-14, 5.710239e-14, 
    5.703244e-14, 5.70991e-14, 5.707889e-14, 5.709937e-14, 5.699675e-14, 
    5.704072e-14, 5.69504e-14, 5.659807e-14, 5.670171e-14, 5.639237e-14, 
    5.620598e-14, 5.608215e-14, 5.599419e-14, 5.600663e-14, 5.603033e-14, 
    5.615211e-14, 5.626657e-14, 5.635372e-14, 5.641197e-14, 5.646936e-14, 
    5.66428e-14, 5.673461e-14, 5.693987e-14, 5.690288e-14, 5.696556e-14, 
    5.702548e-14, 5.712595e-14, 5.710942e-14, 5.715366e-14, 5.696393e-14, 
    5.709004e-14, 5.68818e-14, 5.693878e-14, 5.648481e-14, 5.631165e-14, 
    5.623786e-14, 5.617335e-14, 5.601619e-14, 5.612474e-14, 5.608195e-14, 
    5.618375e-14, 5.624837e-14, 5.621642e-14, 5.641357e-14, 5.633695e-14, 
    5.674005e-14, 5.656656e-14, 5.701849e-14, 5.691048e-14, 5.704437e-14, 
    5.697607e-14, 5.709306e-14, 5.698777e-14, 5.717014e-14, 5.720979e-14, 
    5.718269e-14, 5.728683e-14, 5.698193e-14, 5.709909e-14, 5.621552e-14, 
    5.622073e-14, 5.624502e-14, 5.613821e-14, 5.613168e-14, 5.603377e-14, 
    5.612091e-14, 5.615799e-14, 5.625213e-14, 5.630776e-14, 5.636063e-14, 
    5.647682e-14, 5.660643e-14, 5.678752e-14, 5.691748e-14, 5.700454e-14, 
    5.695117e-14, 5.699828e-14, 5.694561e-14, 5.692092e-14, 5.719492e-14, 
    5.704112e-14, 5.727185e-14, 5.72591e-14, 5.715471e-14, 5.726054e-14, 
    5.622439e-14, 5.61944e-14, 5.609017e-14, 5.617174e-14, 5.60231e-14, 
    5.61063e-14, 5.615411e-14, 5.633852e-14, 5.637904e-14, 5.641655e-14, 
    5.649065e-14, 5.658567e-14, 5.67522e-14, 5.689693e-14, 5.702897e-14, 
    5.70193e-14, 5.70227e-14, 5.705216e-14, 5.697915e-14, 5.706415e-14, 
    5.70784e-14, 5.704112e-14, 5.725739e-14, 5.719564e-14, 5.725883e-14, 
    5.721863e-14, 5.620415e-14, 5.625462e-14, 5.622735e-14, 5.627862e-14, 
    5.624249e-14, 5.640303e-14, 5.645112e-14, 5.667601e-14, 5.65838e-14, 
    5.673057e-14, 5.659872e-14, 5.662209e-14, 5.673528e-14, 5.660586e-14, 
    5.688892e-14, 5.669703e-14, 5.705331e-14, 5.686185e-14, 5.70653e-14, 
    5.70284e-14, 5.708951e-14, 5.71442e-14, 5.7213e-14, 5.733981e-14, 
    5.731047e-14, 5.741647e-14, 5.632984e-14, 5.639522e-14, 5.638949e-14, 
    5.645791e-14, 5.650848e-14, 5.661806e-14, 5.679361e-14, 5.672763e-14, 
    5.684876e-14, 5.687302e-14, 5.668904e-14, 5.680202e-14, 5.643898e-14, 
    5.649767e-14, 5.646276e-14, 5.633498e-14, 5.674279e-14, 5.653363e-14, 
    5.691962e-14, 5.680653e-14, 5.71364e-14, 5.69724e-14, 5.72943e-14, 
    5.74316e-14, 5.756084e-14, 5.771153e-14, 5.643092e-14, 5.638651e-14, 
    5.646605e-14, 5.657598e-14, 5.667798e-14, 5.681343e-14, 5.682729e-14, 
    5.685264e-14, 5.691828e-14, 5.697346e-14, 5.686062e-14, 5.69873e-14, 
    5.651122e-14, 5.676095e-14, 5.636968e-14, 5.648758e-14, 5.656952e-14, 
    5.653361e-14, 5.672009e-14, 5.6764e-14, 5.694224e-14, 5.685016e-14, 
    5.73977e-14, 5.71557e-14, 5.782627e-14, 5.763919e-14, 5.637098e-14, 
    5.643079e-14, 5.663869e-14, 5.653981e-14, 5.682248e-14, 5.689192e-14, 
    5.69484e-14, 5.702052e-14, 5.702833e-14, 5.707104e-14, 5.700104e-14, 
    5.706829e-14, 5.681371e-14, 5.692753e-14, 5.661498e-14, 5.66911e-14, 
    5.66561e-14, 5.661767e-14, 5.673624e-14, 5.686237e-14, 5.686511e-14, 
    5.690553e-14, 5.701928e-14, 5.682362e-14, 5.742881e-14, 5.705527e-14, 
    5.649597e-14, 5.661098e-14, 5.662745e-14, 5.658291e-14, 5.688496e-14, 
    5.67756e-14, 5.707001e-14, 5.69905e-14, 5.712076e-14, 5.705604e-14, 
    5.704652e-14, 5.696337e-14, 5.691155e-14, 5.678061e-14, 5.667397e-14, 
    5.658937e-14, 5.660905e-14, 5.670197e-14, 5.687009e-14, 5.702901e-14, 
    5.699421e-14, 5.711086e-14, 5.6802e-14, 5.693155e-14, 5.688147e-14, 
    5.701203e-14, 5.672586e-14, 5.696944e-14, 5.666351e-14, 5.669037e-14, 
    5.677343e-14, 5.694031e-14, 5.697728e-14, 5.701665e-14, 5.699237e-14, 
    5.687437e-14, 5.685507e-14, 5.677142e-14, 5.67483e-14, 5.668453e-14, 
    5.663169e-14, 5.667996e-14, 5.673061e-14, 5.687443e-14, 5.700391e-14, 
    5.714497e-14, 5.717948e-14, 5.734394e-14, 5.721001e-14, 5.743088e-14, 
    5.724302e-14, 5.756809e-14, 5.698362e-14, 5.723759e-14, 5.677722e-14, 
    5.682691e-14, 5.691665e-14, 5.712242e-14, 5.701142e-14, 5.714126e-14, 
    5.685432e-14, 5.670515e-14, 5.666659e-14, 5.659451e-14, 5.666823e-14, 
    5.666224e-14, 5.673275e-14, 5.67101e-14, 5.687921e-14, 5.678841e-14, 
    5.704627e-14, 5.714024e-14, 5.740535e-14, 5.756758e-14, 5.77326e-14, 
    5.780536e-14, 5.78275e-14, 5.783675e-14 ;

 LITR3C_vr =
  0.0005754704, 0.0005754697, 0.0005754699, 0.0005754694, 0.0005754697, 
    0.0005754693, 0.0005754703, 0.0005754697, 0.00057547, 0.0005754703, 
    0.0005754685, 0.0005754694, 0.0005754675, 0.0005754681, 0.0005754666, 
    0.0005754676, 0.0005754664, 0.0005754667, 0.000575466, 0.0005754662, 
    0.0005754653, 0.0005754659, 0.0005754649, 0.0005754654, 0.0005754654, 
    0.0005754659, 0.0005754692, 0.0005754686, 0.0005754692, 0.0005754692, 
    0.0005754692, 0.0005754697, 0.0005754699, 0.0005754704, 0.0005754703, 
    0.0005754699, 0.0005754691, 0.0005754694, 0.0005754686, 0.0005754687, 
    0.0005754679, 0.0005754682, 0.0005754669, 0.0005754672, 0.0005754661, 
    0.0005754664, 0.0005754662, 0.0005754663, 0.0005754662, 0.0005754666, 
    0.0005754664, 0.0005754668, 0.0005754682, 0.0005754678, 0.000575469, 
    0.0005754697, 0.0005754702, 0.0005754706, 0.0005754705, 0.0005754704, 
    0.0005754699, 0.0005754695, 0.0005754692, 0.0005754689, 0.0005754687, 
    0.000575468, 0.0005754677, 0.0005754668, 0.000575467, 0.0005754667, 
    0.0005754665, 0.0005754661, 0.0005754661, 0.000575466, 0.0005754667, 
    0.0005754662, 0.000575467, 0.0005754668, 0.0005754686, 0.0005754693, 
    0.0005754696, 0.0005754699, 0.0005754705, 0.00057547, 0.0005754702, 
    0.0005754698, 0.0005754696, 0.0005754697, 0.0005754689, 0.0005754692, 
    0.0005754676, 0.0005754683, 0.0005754665, 0.000575467, 0.0005754664, 
    0.0005754667, 0.0005754662, 0.0005754666, 0.0005754659, 0.0005754657, 
    0.0005754658, 0.0005754654, 0.0005754667, 0.0005754662, 0.0005754697, 
    0.0005754697, 0.0005754696, 0.00057547, 0.00057547, 0.0005754704, 
    0.0005754701, 0.0005754699, 0.0005754696, 0.0005754693, 0.0005754691, 
    0.0005754686, 0.0005754681, 0.0005754674, 0.0005754669, 0.0005754665, 
    0.0005754668, 0.0005754666, 0.0005754668, 0.0005754669, 0.0005754658, 
    0.0005754664, 0.0005754655, 0.0005754656, 0.000575466, 0.0005754656, 
    0.0005754696, 0.0005754698, 0.0005754702, 0.0005754699, 0.0005754704, 
    0.0005754702, 0.0005754699, 0.0005754692, 0.0005754691, 0.0005754689, 
    0.0005754686, 0.0005754682, 0.0005754675, 0.000575467, 0.0005754664, 
    0.0005754665, 0.0005754665, 0.0005754664, 0.0005754667, 0.0005754663, 
    0.0005754663, 0.0005754664, 0.0005754656, 0.0005754658, 0.0005754656, 
    0.0005754657, 0.0005754697, 0.0005754695, 0.0005754696, 0.0005754695, 
    0.0005754696, 0.0005754689, 0.0005754688, 0.0005754679, 0.0005754682, 
    0.0005754677, 0.0005754682, 0.0005754681, 0.0005754676, 0.0005754681, 
    0.000575467, 0.0005754678, 0.0005754664, 0.0005754671, 0.0005754663, 
    0.0005754664, 0.0005754662, 0.000575466, 0.0005754657, 0.0005754652, 
    0.0005754653, 0.0005754649, 0.0005754692, 0.000575469, 0.000575469, 
    0.0005754687, 0.0005754685, 0.0005754681, 0.0005754674, 0.0005754677, 
    0.0005754672, 0.0005754671, 0.0005754678, 0.0005754674, 0.0005754688, 
    0.0005754686, 0.0005754687, 0.0005754692, 0.0005754676, 0.0005754684, 
    0.0005754669, 0.0005754674, 0.000575466, 0.0005754667, 0.0005754654, 
    0.0005754649, 0.0005754643, 0.0005754638, 0.0005754688, 0.000575469, 
    0.0005754687, 0.0005754682, 0.0005754678, 0.0005754673, 0.0005754672, 
    0.0005754671, 0.0005754669, 0.0005754667, 0.0005754671, 0.0005754666, 
    0.0005754685, 0.0005754675, 0.0005754691, 0.0005754686, 0.0005754683, 
    0.0005754684, 0.0005754677, 0.0005754675, 0.0005754668, 0.0005754672, 
    0.000575465, 0.000575466, 0.0005754633, 0.000575464, 0.0005754691, 
    0.0005754688, 0.000575468, 0.0005754684, 0.0005754673, 0.000575467, 
    0.0005754668, 0.0005754665, 0.0005754664, 0.0005754663, 0.0005754665, 
    0.0005754663, 0.0005754673, 0.0005754668, 0.0005754681, 0.0005754678, 
    0.0005754679, 0.0005754681, 0.0005754676, 0.0005754671, 0.0005754671, 
    0.000575467, 0.0005754665, 0.0005754672, 0.0005754649, 0.0005754664, 
    0.0005754686, 0.0005754681, 0.0005754681, 0.0005754682, 0.000575467, 
    0.0005754675, 0.0005754663, 0.0005754666, 0.0005754661, 0.0005754664, 
    0.0005754664, 0.0005754667, 0.0005754669, 0.0005754674, 0.0005754679, 
    0.0005754682, 0.0005754681, 0.0005754678, 0.0005754671, 0.0005754664, 
    0.0005754666, 0.0005754661, 0.0005754674, 0.0005754668, 0.000575467, 
    0.0005754665, 0.0005754677, 0.0005754667, 0.0005754679, 0.0005754678, 
    0.0005754675, 0.0005754668, 0.0005754667, 0.0005754665, 0.0005754666, 
    0.0005754671, 0.0005754671, 0.0005754675, 0.0005754676, 0.0005754678, 
    0.0005754681, 0.0005754678, 0.0005754677, 0.0005754671, 0.0005754665, 
    0.000575466, 0.0005754658, 0.0005754652, 0.0005754657, 0.0005754649, 
    0.0005754656, 0.0005754643, 0.0005754667, 0.0005754656, 0.0005754675, 
    0.0005754672, 0.0005754669, 0.0005754661, 0.0005754665, 0.000575466, 
    0.0005754671, 0.0005754678, 0.0005754679, 0.0005754682, 0.0005754679, 
    0.0005754679, 0.0005754677, 0.0005754677, 0.0005754671, 0.0005754674, 
    0.0005754664, 0.000575466, 0.000575465, 0.0005754643, 0.0005754636, 
    0.0005754633, 0.0005754633, 0.0005754632,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.394736e-07, 1.394735e-07, 1.394735e-07, 1.394734e-07, 1.394735e-07, 
    1.394734e-07, 1.394736e-07, 1.394735e-07, 1.394736e-07, 1.394736e-07, 
    1.394732e-07, 1.394734e-07, 1.394729e-07, 1.394731e-07, 1.394727e-07, 
    1.39473e-07, 1.394727e-07, 1.394727e-07, 1.394726e-07, 1.394726e-07, 
    1.394724e-07, 1.394725e-07, 1.394723e-07, 1.394724e-07, 1.394724e-07, 
    1.394725e-07, 1.394733e-07, 1.394732e-07, 1.394734e-07, 1.394733e-07, 
    1.394733e-07, 1.394735e-07, 1.394735e-07, 1.394736e-07, 1.394736e-07, 
    1.394735e-07, 1.394733e-07, 1.394734e-07, 1.394732e-07, 1.394732e-07, 
    1.39473e-07, 1.394731e-07, 1.394728e-07, 1.394729e-07, 1.394726e-07, 
    1.394727e-07, 1.394726e-07, 1.394726e-07, 1.394726e-07, 1.394727e-07, 
    1.394727e-07, 1.394728e-07, 1.394731e-07, 1.39473e-07, 1.394733e-07, 
    1.394735e-07, 1.394736e-07, 1.394737e-07, 1.394737e-07, 1.394737e-07, 
    1.394735e-07, 1.394734e-07, 1.394733e-07, 1.394733e-07, 1.394732e-07, 
    1.394731e-07, 1.39473e-07, 1.394728e-07, 1.394728e-07, 1.394727e-07, 
    1.394727e-07, 1.394726e-07, 1.394726e-07, 1.394726e-07, 1.394727e-07, 
    1.394726e-07, 1.394728e-07, 1.394728e-07, 1.394732e-07, 1.394734e-07, 
    1.394734e-07, 1.394735e-07, 1.394737e-07, 1.394736e-07, 1.394736e-07, 
    1.394735e-07, 1.394734e-07, 1.394735e-07, 1.394733e-07, 1.394734e-07, 
    1.39473e-07, 1.394731e-07, 1.394727e-07, 1.394728e-07, 1.394727e-07, 
    1.394727e-07, 1.394726e-07, 1.394727e-07, 1.394725e-07, 1.394725e-07, 
    1.394725e-07, 1.394724e-07, 1.394727e-07, 1.394726e-07, 1.394735e-07, 
    1.394735e-07, 1.394734e-07, 1.394735e-07, 1.394736e-07, 1.394736e-07, 
    1.394736e-07, 1.394735e-07, 1.394734e-07, 1.394734e-07, 1.394733e-07, 
    1.394732e-07, 1.394731e-07, 1.394729e-07, 1.394728e-07, 1.394727e-07, 
    1.394728e-07, 1.394727e-07, 1.394728e-07, 1.394728e-07, 1.394725e-07, 
    1.394727e-07, 1.394724e-07, 1.394725e-07, 1.394726e-07, 1.394725e-07, 
    1.394735e-07, 1.394735e-07, 1.394736e-07, 1.394735e-07, 1.394737e-07, 
    1.394736e-07, 1.394735e-07, 1.394734e-07, 1.394733e-07, 1.394733e-07, 
    1.394732e-07, 1.394731e-07, 1.39473e-07, 1.394728e-07, 1.394727e-07, 
    1.394727e-07, 1.394727e-07, 1.394727e-07, 1.394727e-07, 1.394726e-07, 
    1.394726e-07, 1.394727e-07, 1.394725e-07, 1.394725e-07, 1.394725e-07, 
    1.394725e-07, 1.394735e-07, 1.394734e-07, 1.394735e-07, 1.394734e-07, 
    1.394734e-07, 1.394733e-07, 1.394732e-07, 1.39473e-07, 1.394731e-07, 
    1.39473e-07, 1.394731e-07, 1.394731e-07, 1.39473e-07, 1.394731e-07, 
    1.394728e-07, 1.39473e-07, 1.394727e-07, 1.394728e-07, 1.394726e-07, 
    1.394727e-07, 1.394726e-07, 1.394726e-07, 1.394725e-07, 1.394724e-07, 
    1.394724e-07, 1.394723e-07, 1.394734e-07, 1.394733e-07, 1.394733e-07, 
    1.394732e-07, 1.394732e-07, 1.394731e-07, 1.394729e-07, 1.39473e-07, 
    1.394729e-07, 1.394728e-07, 1.39473e-07, 1.394729e-07, 1.394733e-07, 
    1.394732e-07, 1.394732e-07, 1.394734e-07, 1.39473e-07, 1.394732e-07, 
    1.394728e-07, 1.394729e-07, 1.394726e-07, 1.394727e-07, 1.394724e-07, 
    1.394723e-07, 1.394722e-07, 1.39472e-07, 1.394733e-07, 1.394733e-07, 
    1.394732e-07, 1.394731e-07, 1.39473e-07, 1.394729e-07, 1.394729e-07, 
    1.394729e-07, 1.394728e-07, 1.394727e-07, 1.394728e-07, 1.394727e-07, 
    1.394732e-07, 1.394729e-07, 1.394733e-07, 1.394732e-07, 1.394731e-07, 
    1.394732e-07, 1.39473e-07, 1.394729e-07, 1.394728e-07, 1.394729e-07, 
    1.394723e-07, 1.394726e-07, 1.394719e-07, 1.394721e-07, 1.394733e-07, 
    1.394733e-07, 1.394731e-07, 1.394732e-07, 1.394729e-07, 1.394728e-07, 
    1.394728e-07, 1.394727e-07, 1.394727e-07, 1.394726e-07, 1.394727e-07, 
    1.394726e-07, 1.394729e-07, 1.394728e-07, 1.394731e-07, 1.39473e-07, 
    1.39473e-07, 1.394731e-07, 1.39473e-07, 1.394728e-07, 1.394728e-07, 
    1.394728e-07, 1.394727e-07, 1.394729e-07, 1.394723e-07, 1.394727e-07, 
    1.394732e-07, 1.394731e-07, 1.394731e-07, 1.394731e-07, 1.394728e-07, 
    1.394729e-07, 1.394726e-07, 1.394727e-07, 1.394726e-07, 1.394727e-07, 
    1.394727e-07, 1.394727e-07, 1.394728e-07, 1.394729e-07, 1.39473e-07, 
    1.394731e-07, 1.394731e-07, 1.39473e-07, 1.394728e-07, 1.394727e-07, 
    1.394727e-07, 1.394726e-07, 1.394729e-07, 1.394728e-07, 1.394728e-07, 
    1.394727e-07, 1.39473e-07, 1.394727e-07, 1.39473e-07, 1.39473e-07, 
    1.394729e-07, 1.394728e-07, 1.394727e-07, 1.394727e-07, 1.394727e-07, 
    1.394728e-07, 1.394729e-07, 1.394729e-07, 1.39473e-07, 1.39473e-07, 
    1.394731e-07, 1.39473e-07, 1.39473e-07, 1.394728e-07, 1.394727e-07, 
    1.394726e-07, 1.394725e-07, 1.394724e-07, 1.394725e-07, 1.394723e-07, 
    1.394725e-07, 1.394722e-07, 1.394727e-07, 1.394725e-07, 1.394729e-07, 
    1.394729e-07, 1.394728e-07, 1.394726e-07, 1.394727e-07, 1.394726e-07, 
    1.394729e-07, 1.39473e-07, 1.39473e-07, 1.394731e-07, 1.39473e-07, 
    1.39473e-07, 1.39473e-07, 1.39473e-07, 1.394728e-07, 1.394729e-07, 
    1.394727e-07, 1.394726e-07, 1.394723e-07, 1.394722e-07, 1.39472e-07, 
    1.394719e-07, 1.394719e-07, 1.394719e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  6.862535e-26, 6.372354e-26, 2.941087e-26, 3.798904e-26, -4.779266e-26, 
    4.534175e-26, 7.965443e-26, -1.372507e-25, 1.347998e-26, -9.803622e-27, 
    -9.681077e-26, 2.450905e-26, -5.269447e-26, -2.205815e-26, 0, 
    2.08327e-26, -4.166539e-26, 9.068351e-26, -1.838179e-26, -2.450906e-27, 
    -5.146902e-26, -7.842898e-26, -2.450905e-26, 3.308722e-26, 1.225453e-25, 
    2.450906e-27, 4.166539e-26, -4.901811e-27, 9.803622e-27, -4.043994e-26, 
    -7.597807e-26, -5.146902e-26, 4.901811e-26, -1.004871e-25, 8.578169e-27, 
    8.578169e-27, -4.65672e-26, -2.08327e-26, 2.450905e-26, 5.637083e-26, 
    -3.798904e-26, -1.715634e-26, -9.803622e-27, -2.941087e-26, 
    -5.146902e-26, -1.617598e-25, 5.514538e-26, 6.249809e-26, 1.838179e-26, 
    -4.901811e-27, 7.352717e-27, 8.700715e-26, 2.205815e-26, 3.308722e-26, 
    -6.4949e-26, 8.087988e-26, -5.514538e-26, 5.024356e-26, -7.107626e-26, 
    7.475262e-26, 4.901811e-26, -1.838179e-26, 5.514538e-26, 6.004719e-26, 
    3.921449e-26, 1.715634e-26, 6.372354e-26, 6.617445e-26, 1.666616e-25, 
    5.882173e-26, -7.842898e-26, 9.435986e-26, 3.676358e-26, 9.803622e-26, 
    9.313441e-26, -2.450905e-26, 1.470543e-26, -1.139671e-25, -2.450906e-27, 
    1.102908e-26, 8.700715e-26, 7.652491e-42, 1.470543e-26, -1.727888e-25, 
    -6.98508e-26, 0, -4.779266e-26, 1.286725e-25, -7.352717e-26, 
    1.666616e-25, 2.573451e-26, -2.818541e-26, -9.068351e-26, -1.29898e-25, 
    5.514538e-26, 4.534175e-26, -6.617445e-26, -3.921449e-26, -2.573451e-26, 
    -9.313441e-26, 7.107626e-26, 7.720352e-26, -1.225453e-26, -3.676358e-26, 
    1.311234e-25, -2.450906e-27, 8.210533e-26, 7.352717e-27, -7.475262e-26, 
    1.715634e-26, -2.695996e-26, -6.127264e-27, -1.470543e-26, -5.024356e-26, 
    5.759628e-26, 2.32836e-26, -1.960724e-26, -2.818541e-26, -1.715634e-26, 
    1.225453e-26, 1.053889e-25, 8.700715e-26, 2.08327e-26, 1.470543e-26, 
    -4.41163e-26, -1.593089e-26, 1.887197e-25, -4.65672e-26, 2.695996e-26, 
    1.102908e-26, 1.593089e-26, 1.838179e-26, -1.715634e-26, 1.188689e-25, 
    -3.308722e-26, 3.676358e-26, -5.514538e-26, 6.4949e-26, 1.372507e-25, 
    1.54407e-25, -3.676358e-26, 4.901811e-27, -9.803622e-26, -6.127264e-26, 
    -1.715634e-26, -7.107626e-26, 3.431268e-26, -4.901811e-27, -1.225453e-27, 
    1.066144e-25, 1.041635e-25, -1.237707e-25, 0, 1.470543e-25, 
    -8.210533e-26, -8.578169e-27, -2.08327e-26, 3.186177e-26, -3.676358e-26, 
    -4.901811e-27, -4.901811e-27, 2.695996e-26, 9.068351e-26, -3.063632e-26, 
    4.41163e-26, 8.455624e-26, 2.08327e-26, -2.450906e-27, 1.078398e-25, 
    4.166539e-26, 1.764652e-25, 9.313441e-26, 6.617445e-26, -1.139671e-25, 
    8.210533e-26, 9.803622e-26, 1.482798e-25, 3.308722e-26, 4.043994e-26, 
    3.063632e-26, 5.391992e-26, -1.347998e-26, 8.82326e-26, -7.965443e-26, 
    -6.862535e-26, -1.715634e-26, 1.482798e-25, 1.409271e-25, -1.470543e-26, 
    4.289085e-26, -1.102908e-26, -7.597807e-26, 1.347998e-25, 5.637083e-26, 
    6.4949e-26, 1.960724e-26, 6.372354e-26, -3.676358e-26, 4.289085e-26, 
    1.960724e-26, -1.102908e-26, 8.333079e-26, -1.115162e-25, -5.024356e-26, 
    4.901811e-26, 2.695996e-26, -5.024356e-26, 4.534175e-26, 6.862535e-26, 
    3.431268e-26, 0, -1.237707e-25, -6.98508e-26, 6.73999e-26, 1.67887e-25, 
    -6.004719e-26, 6.249809e-26, -1.470543e-26, 9.558531e-26, 4.779266e-26, 
    3.798904e-26, -4.289085e-26, 7.230172e-26, 5.269447e-26, -9.803622e-26, 
    -1.176435e-25, 1.617598e-25, -5.391992e-26, 1.54407e-25, 1.715634e-26, 
    5.146902e-26, -6.4949e-26, 1.16418e-25, -3.186177e-26, -9.068351e-26, 
    8.578169e-27, -5.269447e-26, 8.087988e-26, -2.08327e-26, 1.617598e-25, 
    -5.146902e-26, -8.087988e-26, 4.534175e-26, -3.921449e-26, -4.043994e-26, 
    4.289085e-26, -8.578169e-27, -2.573451e-26, 0, 2.695996e-26, 8.82326e-26, 
    3.798904e-26, -6.862535e-26, 6.617445e-26, 6.249809e-26, 3.676358e-26, 
    -2.573451e-26, 1.090653e-25, 4.166539e-26, 6.4949e-26, 7.842898e-26, 
    4.901811e-26, 5.146902e-26, -7.352717e-27, 7.965443e-26, 6.98508e-26, 
    -1.470543e-26, 1.470543e-26, 7.720352e-26, -8.578169e-26, 4.043994e-26, 
    -1.078398e-25, -7.107626e-26, 1.053889e-25, -7.965443e-26, 7.475262e-26, 
    -7.352717e-27, 6.004719e-26, -1.176435e-25, -1.56858e-25, -5.146902e-26, 
    1.347998e-26, -1.470543e-26, 1.838179e-26, -2.941087e-26, -4.779266e-26, 
    5.269447e-26, 7.107626e-26, 9.803622e-26, 7.475262e-26, -1.066144e-25, 
    -5.146902e-26, 4.901811e-26, -2.205815e-26, 6.862535e-26, 3.308722e-26, 
    -3.431268e-26, 7.720352e-26, 7.597807e-26, -7.842898e-26, -2.450906e-27, 
    -9.313441e-26, 5.637083e-26, -4.41163e-26, -3.798904e-26, -2.450906e-27, 
    0, -9.926167e-26, 1.470543e-26, -3.308722e-26, 2.573451e-26, 
    4.901811e-26, -1.360253e-25, 6.004719e-26, 6.4949e-26, 1.102908e-26, 
    -2.450905e-26, 6.617445e-26, 2.450906e-27, 3.186177e-26, 1.470543e-26, 
    3.553813e-26, 1.54407e-25, -1.225453e-26, 7.842898e-26, 1.715634e-26, 
    1.470543e-26, -4.166539e-26, 7.842898e-26, 1.715634e-26, 4.534175e-26, 
    8.210533e-26, -7.965443e-26, 3.798904e-26, 1.960724e-26, -1.347998e-26, 
    8.455624e-26, 3.553813e-26,
  1.390974e-32, 1.390972e-32, 1.390973e-32, 1.390971e-32, 1.390972e-32, 
    1.390971e-32, 1.390973e-32, 1.390972e-32, 1.390973e-32, 1.390974e-32, 
    1.390969e-32, 1.390971e-32, 1.390967e-32, 1.390968e-32, 1.390965e-32, 
    1.390967e-32, 1.390964e-32, 1.390965e-32, 1.390963e-32, 1.390963e-32, 
    1.390961e-32, 1.390963e-32, 1.39096e-32, 1.390962e-32, 1.390962e-32, 
    1.390963e-32, 1.390971e-32, 1.390969e-32, 1.390971e-32, 1.390971e-32, 
    1.390971e-32, 1.390972e-32, 1.390973e-32, 1.390974e-32, 1.390974e-32, 
    1.390973e-32, 1.390971e-32, 1.390971e-32, 1.39097e-32, 1.39097e-32, 
    1.390968e-32, 1.390968e-32, 1.390965e-32, 1.390966e-32, 1.390963e-32, 
    1.390964e-32, 1.390963e-32, 1.390964e-32, 1.390963e-32, 1.390965e-32, 
    1.390964e-32, 1.390965e-32, 1.390968e-32, 1.390967e-32, 1.39097e-32, 
    1.390972e-32, 1.390973e-32, 1.390974e-32, 1.390974e-32, 1.390974e-32, 
    1.390973e-32, 1.390972e-32, 1.390971e-32, 1.39097e-32, 1.39097e-32, 
    1.390968e-32, 1.390967e-32, 1.390965e-32, 1.390965e-32, 1.390965e-32, 
    1.390964e-32, 1.390963e-32, 1.390963e-32, 1.390963e-32, 1.390965e-32, 
    1.390964e-32, 1.390966e-32, 1.390965e-32, 1.39097e-32, 1.390971e-32, 
    1.390972e-32, 1.390972e-32, 1.390974e-32, 1.390973e-32, 1.390973e-32, 
    1.390972e-32, 1.390972e-32, 1.390972e-32, 1.39097e-32, 1.390971e-32, 
    1.390967e-32, 1.390969e-32, 1.390964e-32, 1.390965e-32, 1.390964e-32, 
    1.390965e-32, 1.390964e-32, 1.390965e-32, 1.390963e-32, 1.390962e-32, 
    1.390963e-32, 1.390962e-32, 1.390965e-32, 1.390963e-32, 1.390972e-32, 
    1.390972e-32, 1.390972e-32, 1.390973e-32, 1.390973e-32, 1.390974e-32, 
    1.390973e-32, 1.390973e-32, 1.390972e-32, 1.390971e-32, 1.390971e-32, 
    1.39097e-32, 1.390968e-32, 1.390967e-32, 1.390965e-32, 1.390964e-32, 
    1.390965e-32, 1.390965e-32, 1.390965e-32, 1.390965e-32, 1.390963e-32, 
    1.390964e-32, 1.390962e-32, 1.390962e-32, 1.390963e-32, 1.390962e-32, 
    1.390972e-32, 1.390972e-32, 1.390973e-32, 1.390973e-32, 1.390974e-32, 
    1.390973e-32, 1.390973e-32, 1.390971e-32, 1.390971e-32, 1.39097e-32, 
    1.390969e-32, 1.390968e-32, 1.390967e-32, 1.390966e-32, 1.390964e-32, 
    1.390964e-32, 1.390964e-32, 1.390964e-32, 1.390965e-32, 1.390964e-32, 
    1.390964e-32, 1.390964e-32, 1.390962e-32, 1.390963e-32, 1.390962e-32, 
    1.390962e-32, 1.390972e-32, 1.390972e-32, 1.390972e-32, 1.390971e-32, 
    1.390972e-32, 1.39097e-32, 1.39097e-32, 1.390968e-32, 1.390968e-32, 
    1.390967e-32, 1.390968e-32, 1.390968e-32, 1.390967e-32, 1.390968e-32, 
    1.390966e-32, 1.390967e-32, 1.390964e-32, 1.390966e-32, 1.390964e-32, 
    1.390964e-32, 1.390964e-32, 1.390963e-32, 1.390962e-32, 1.390961e-32, 
    1.390961e-32, 1.39096e-32, 1.390971e-32, 1.39097e-32, 1.39097e-32, 
    1.39097e-32, 1.390969e-32, 1.390968e-32, 1.390966e-32, 1.390967e-32, 
    1.390966e-32, 1.390966e-32, 1.390967e-32, 1.390966e-32, 1.39097e-32, 
    1.390969e-32, 1.39097e-32, 1.390971e-32, 1.390967e-32, 1.390969e-32, 
    1.390965e-32, 1.390966e-32, 1.390963e-32, 1.390965e-32, 1.390962e-32, 
    1.39096e-32, 1.390959e-32, 1.390958e-32, 1.39097e-32, 1.39097e-32, 
    1.39097e-32, 1.390969e-32, 1.390968e-32, 1.390966e-32, 1.390966e-32, 
    1.390966e-32, 1.390965e-32, 1.390965e-32, 1.390966e-32, 1.390965e-32, 
    1.390969e-32, 1.390967e-32, 1.390971e-32, 1.39097e-32, 1.390969e-32, 
    1.390969e-32, 1.390967e-32, 1.390967e-32, 1.390965e-32, 1.390966e-32, 
    1.390961e-32, 1.390963e-32, 1.390956e-32, 1.390958e-32, 1.390971e-32, 
    1.39097e-32, 1.390968e-32, 1.390969e-32, 1.390966e-32, 1.390966e-32, 
    1.390965e-32, 1.390964e-32, 1.390964e-32, 1.390964e-32, 1.390965e-32, 
    1.390964e-32, 1.390966e-32, 1.390965e-32, 1.390968e-32, 1.390967e-32, 
    1.390968e-32, 1.390968e-32, 1.390967e-32, 1.390966e-32, 1.390966e-32, 
    1.390965e-32, 1.390964e-32, 1.390966e-32, 1.39096e-32, 1.390964e-32, 
    1.390969e-32, 1.390968e-32, 1.390968e-32, 1.390968e-32, 1.390966e-32, 
    1.390967e-32, 1.390964e-32, 1.390965e-32, 1.390963e-32, 1.390964e-32, 
    1.390964e-32, 1.390965e-32, 1.390965e-32, 1.390967e-32, 1.390968e-32, 
    1.390968e-32, 1.390968e-32, 1.390967e-32, 1.390966e-32, 1.390964e-32, 
    1.390965e-32, 1.390963e-32, 1.390966e-32, 1.390965e-32, 1.390966e-32, 
    1.390964e-32, 1.390967e-32, 1.390965e-32, 1.390968e-32, 1.390967e-32, 
    1.390967e-32, 1.390965e-32, 1.390965e-32, 1.390964e-32, 1.390965e-32, 
    1.390966e-32, 1.390966e-32, 1.390967e-32, 1.390967e-32, 1.390968e-32, 
    1.390968e-32, 1.390968e-32, 1.390967e-32, 1.390966e-32, 1.390965e-32, 
    1.390963e-32, 1.390963e-32, 1.390961e-32, 1.390962e-32, 1.39096e-32, 
    1.390962e-32, 1.390959e-32, 1.390965e-32, 1.390962e-32, 1.390967e-32, 
    1.390966e-32, 1.390965e-32, 1.390963e-32, 1.390964e-32, 1.390963e-32, 
    1.390966e-32, 1.390967e-32, 1.390968e-32, 1.390968e-32, 1.390968e-32, 
    1.390968e-32, 1.390967e-32, 1.390967e-32, 1.390966e-32, 1.390967e-32, 
    1.390964e-32, 1.390963e-32, 1.390961e-32, 1.390959e-32, 1.390957e-32, 
    1.390957e-32, 1.390956e-32, 1.390956e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.55127e-15, 1.555453e-15, 1.55464e-15, 1.558011e-15, 1.556142e-15, 
    1.558348e-15, 1.552119e-15, 1.555618e-15, 1.553385e-15, 1.551647e-15, 
    1.564543e-15, 1.558162e-15, 1.571166e-15, 1.567103e-15, 1.577302e-15, 
    1.570534e-15, 1.578666e-15, 1.577108e-15, 1.581797e-15, 1.580455e-15, 
    1.586443e-15, 1.582417e-15, 1.589546e-15, 1.585483e-15, 1.586118e-15, 
    1.582284e-15, 1.559448e-15, 1.563749e-15, 1.559193e-15, 1.559806e-15, 
    1.559531e-15, 1.55618e-15, 1.55449e-15, 1.550951e-15, 1.551593e-15, 
    1.554193e-15, 1.560082e-15, 1.558085e-15, 1.563119e-15, 1.563006e-15, 
    1.568602e-15, 1.56608e-15, 1.575474e-15, 1.572807e-15, 1.580511e-15, 
    1.578574e-15, 1.58042e-15, 1.57986e-15, 1.580427e-15, 1.577587e-15, 
    1.578804e-15, 1.576304e-15, 1.566552e-15, 1.56942e-15, 1.560858e-15, 
    1.555699e-15, 1.552272e-15, 1.549837e-15, 1.550182e-15, 1.550837e-15, 
    1.554208e-15, 1.557376e-15, 1.559788e-15, 1.561401e-15, 1.562989e-15, 
    1.56779e-15, 1.570331e-15, 1.576012e-15, 1.574989e-15, 1.576723e-15, 
    1.578382e-15, 1.581163e-15, 1.580705e-15, 1.58193e-15, 1.576678e-15, 
    1.580169e-15, 1.574405e-15, 1.575982e-15, 1.563417e-15, 1.558624e-15, 
    1.556582e-15, 1.554796e-15, 1.550446e-15, 1.553451e-15, 1.552266e-15, 
    1.555084e-15, 1.556873e-15, 1.555988e-15, 1.561445e-15, 1.559324e-15, 
    1.570482e-15, 1.56568e-15, 1.578188e-15, 1.575199e-15, 1.578905e-15, 
    1.577014e-15, 1.580253e-15, 1.577338e-15, 1.582386e-15, 1.583483e-15, 
    1.582733e-15, 1.585616e-15, 1.577177e-15, 1.580419e-15, 1.555963e-15, 
    1.556108e-15, 1.55678e-15, 1.553823e-15, 1.553643e-15, 1.550933e-15, 
    1.553345e-15, 1.554371e-15, 1.556977e-15, 1.558516e-15, 1.55998e-15, 
    1.563196e-15, 1.566783e-15, 1.571796e-15, 1.575393e-15, 1.577802e-15, 
    1.576325e-15, 1.577629e-15, 1.576171e-15, 1.575488e-15, 1.583072e-15, 
    1.578815e-15, 1.585201e-15, 1.584848e-15, 1.581959e-15, 1.584888e-15, 
    1.556209e-15, 1.555379e-15, 1.552494e-15, 1.554752e-15, 1.550637e-15, 
    1.55294e-15, 1.554264e-15, 1.559368e-15, 1.560489e-15, 1.561528e-15, 
    1.563579e-15, 1.566209e-15, 1.570818e-15, 1.574824e-15, 1.578478e-15, 
    1.578211e-15, 1.578305e-15, 1.57912e-15, 1.577099e-15, 1.579452e-15, 
    1.579846e-15, 1.578815e-15, 1.584801e-15, 1.583092e-15, 1.584841e-15, 
    1.583728e-15, 1.555649e-15, 1.557046e-15, 1.556291e-15, 1.55771e-15, 
    1.55671e-15, 1.561153e-15, 1.562485e-15, 1.568709e-15, 1.566157e-15, 
    1.570219e-15, 1.56657e-15, 1.567216e-15, 1.57035e-15, 1.566767e-15, 
    1.574602e-15, 1.569291e-15, 1.579152e-15, 1.573853e-15, 1.579484e-15, 
    1.578463e-15, 1.580154e-15, 1.581668e-15, 1.583572e-15, 1.587082e-15, 
    1.58627e-15, 1.589204e-15, 1.559127e-15, 1.560937e-15, 1.560779e-15, 
    1.562672e-15, 1.564072e-15, 1.567105e-15, 1.571964e-15, 1.570138e-15, 
    1.573491e-15, 1.574162e-15, 1.56907e-15, 1.572197e-15, 1.562149e-15, 
    1.563773e-15, 1.562806e-15, 1.55927e-15, 1.570558e-15, 1.564768e-15, 
    1.575452e-15, 1.572322e-15, 1.581452e-15, 1.576913e-15, 1.585822e-15, 
    1.589623e-15, 1.5932e-15, 1.597371e-15, 1.561925e-15, 1.560696e-15, 
    1.562898e-15, 1.56594e-15, 1.568764e-15, 1.572513e-15, 1.572896e-15, 
    1.573598e-15, 1.575415e-15, 1.576942e-15, 1.573819e-15, 1.577325e-15, 
    1.564148e-15, 1.57106e-15, 1.56023e-15, 1.563494e-15, 1.565761e-15, 
    1.564768e-15, 1.569929e-15, 1.571144e-15, 1.576078e-15, 1.573529e-15, 
    1.588684e-15, 1.581986e-15, 1.600546e-15, 1.595368e-15, 1.560266e-15, 
    1.561922e-15, 1.567676e-15, 1.564939e-15, 1.572763e-15, 1.574685e-15, 
    1.576249e-15, 1.578245e-15, 1.578461e-15, 1.579643e-15, 1.577705e-15, 
    1.579567e-15, 1.57252e-15, 1.575671e-15, 1.56702e-15, 1.569127e-15, 
    1.568158e-15, 1.567094e-15, 1.570376e-15, 1.573867e-15, 1.573943e-15, 
    1.575062e-15, 1.57821e-15, 1.572795e-15, 1.589545e-15, 1.579206e-15, 
    1.563726e-15, 1.566909e-15, 1.567365e-15, 1.566132e-15, 1.574492e-15, 
    1.571466e-15, 1.579614e-15, 1.577414e-15, 1.581019e-15, 1.579228e-15, 
    1.578964e-15, 1.576662e-15, 1.575229e-15, 1.571604e-15, 1.568653e-15, 
    1.566311e-15, 1.566856e-15, 1.569427e-15, 1.574081e-15, 1.57848e-15, 
    1.577516e-15, 1.580745e-15, 1.572196e-15, 1.575782e-15, 1.574396e-15, 
    1.57801e-15, 1.570089e-15, 1.576831e-15, 1.568363e-15, 1.569107e-15, 
    1.571405e-15, 1.576024e-15, 1.577048e-15, 1.578138e-15, 1.577465e-15, 
    1.574199e-15, 1.573665e-15, 1.57135e-15, 1.57071e-15, 1.568945e-15, 
    1.567482e-15, 1.568818e-15, 1.57022e-15, 1.574201e-15, 1.577785e-15, 
    1.581689e-15, 1.582644e-15, 1.587196e-15, 1.583489e-15, 1.589603e-15, 
    1.584403e-15, 1.593401e-15, 1.577223e-15, 1.584253e-15, 1.57151e-15, 
    1.572886e-15, 1.57537e-15, 1.581065e-15, 1.577993e-15, 1.581586e-15, 
    1.573644e-15, 1.569516e-15, 1.568448e-15, 1.566453e-15, 1.568494e-15, 
    1.568328e-15, 1.570279e-15, 1.569652e-15, 1.574333e-15, 1.57182e-15, 
    1.578957e-15, 1.581558e-15, 1.588896e-15, 1.593386e-15, 1.597954e-15, 
    1.599968e-15, 1.600581e-15, 1.600837e-15 ;

 LITR3N_vr =
  7.964089e-06, 7.96408e-06, 7.964082e-06, 7.964075e-06, 7.964079e-06, 
    7.964075e-06, 7.964087e-06, 7.96408e-06, 7.964084e-06, 7.964088e-06, 
    7.964062e-06, 7.964075e-06, 7.964049e-06, 7.964057e-06, 7.964037e-06, 
    7.96405e-06, 7.964034e-06, 7.964037e-06, 7.964028e-06, 7.96403e-06, 
    7.964019e-06, 7.964027e-06, 7.964012e-06, 7.96402e-06, 7.964019e-06, 
    7.964027e-06, 7.964072e-06, 7.964064e-06, 7.964073e-06, 7.964071e-06, 
    7.964072e-06, 7.964079e-06, 7.964082e-06, 7.964089e-06, 7.964088e-06, 
    7.964083e-06, 7.964071e-06, 7.964075e-06, 7.964065e-06, 7.964065e-06, 
    7.964054e-06, 7.964059e-06, 7.96404e-06, 7.964046e-06, 7.96403e-06, 
    7.964034e-06, 7.96403e-06, 7.964031e-06, 7.96403e-06, 7.964036e-06, 
    7.964034e-06, 7.964039e-06, 7.964059e-06, 7.964052e-06, 7.964069e-06, 
    7.964079e-06, 7.964087e-06, 7.964091e-06, 7.964091e-06, 7.964089e-06, 
    7.964083e-06, 7.964077e-06, 7.964071e-06, 7.964069e-06, 7.964065e-06, 
    7.964056e-06, 7.96405e-06, 7.964039e-06, 7.964041e-06, 7.964038e-06, 
    7.964035e-06, 7.964029e-06, 7.96403e-06, 7.964028e-06, 7.964038e-06, 
    7.964031e-06, 7.964042e-06, 7.964039e-06, 7.964064e-06, 7.964074e-06, 
    7.964078e-06, 7.964081e-06, 7.96409e-06, 7.964084e-06, 7.964087e-06, 
    7.964081e-06, 7.964078e-06, 7.964079e-06, 7.964069e-06, 7.964072e-06, 
    7.96405e-06, 7.96406e-06, 7.964035e-06, 7.964041e-06, 7.964034e-06, 
    7.964038e-06, 7.964031e-06, 7.964037e-06, 7.964027e-06, 7.964024e-06, 
    7.964026e-06, 7.96402e-06, 7.964037e-06, 7.96403e-06, 7.964079e-06, 
    7.964079e-06, 7.964078e-06, 7.964084e-06, 7.964084e-06, 7.964089e-06, 
    7.964085e-06, 7.964082e-06, 7.964078e-06, 7.964074e-06, 7.964071e-06, 
    7.964065e-06, 7.964058e-06, 7.964048e-06, 7.96404e-06, 7.964036e-06, 
    7.964039e-06, 7.964036e-06, 7.964039e-06, 7.96404e-06, 7.964025e-06, 
    7.964034e-06, 7.964021e-06, 7.964021e-06, 7.964028e-06, 7.964021e-06, 
    7.964079e-06, 7.96408e-06, 7.964086e-06, 7.964081e-06, 7.96409e-06, 
    7.964085e-06, 7.964083e-06, 7.964072e-06, 7.96407e-06, 7.964069e-06, 
    7.964064e-06, 7.964059e-06, 7.964049e-06, 7.964041e-06, 7.964034e-06, 
    7.964035e-06, 7.964035e-06, 7.964033e-06, 7.964037e-06, 7.964032e-06, 
    7.964031e-06, 7.964034e-06, 7.964022e-06, 7.964025e-06, 7.964022e-06, 
    7.964024e-06, 7.96408e-06, 7.964077e-06, 7.964079e-06, 7.964076e-06, 
    7.964078e-06, 7.964069e-06, 7.964067e-06, 7.964054e-06, 7.964059e-06, 
    7.964051e-06, 7.964059e-06, 7.964057e-06, 7.96405e-06, 7.964058e-06, 
    7.964042e-06, 7.964053e-06, 7.964033e-06, 7.964044e-06, 7.964032e-06, 
    7.964034e-06, 7.964031e-06, 7.964028e-06, 7.964024e-06, 7.964018e-06, 
    7.964019e-06, 7.964013e-06, 7.964073e-06, 7.964069e-06, 7.964069e-06, 
    7.964066e-06, 7.964063e-06, 7.964057e-06, 7.964048e-06, 7.964051e-06, 
    7.964044e-06, 7.964043e-06, 7.964053e-06, 7.964047e-06, 7.964067e-06, 
    7.964064e-06, 7.964066e-06, 7.964073e-06, 7.96405e-06, 7.964062e-06, 
    7.96404e-06, 7.964047e-06, 7.964029e-06, 7.964038e-06, 7.964019e-06, 
    7.964012e-06, 7.964005e-06, 7.963997e-06, 7.964068e-06, 7.964069e-06, 
    7.964066e-06, 7.964059e-06, 7.964054e-06, 7.964047e-06, 7.964046e-06, 
    7.964044e-06, 7.96404e-06, 7.964038e-06, 7.964044e-06, 7.964037e-06, 
    7.964063e-06, 7.964049e-06, 7.96407e-06, 7.964064e-06, 7.964059e-06, 
    7.964062e-06, 7.964051e-06, 7.964049e-06, 7.964039e-06, 7.964044e-06, 
    7.964014e-06, 7.964028e-06, 7.96399e-06, 7.964e-06, 7.96407e-06, 
    7.964068e-06, 7.964056e-06, 7.964061e-06, 7.964046e-06, 7.964042e-06, 
    7.964039e-06, 7.964035e-06, 7.964034e-06, 7.964032e-06, 7.964036e-06, 
    7.964032e-06, 7.964047e-06, 7.96404e-06, 7.964058e-06, 7.964053e-06, 
    7.964055e-06, 7.964057e-06, 7.96405e-06, 7.964044e-06, 7.964043e-06, 
    7.964041e-06, 7.964035e-06, 7.964046e-06, 7.964012e-06, 7.964033e-06, 
    7.964064e-06, 7.964058e-06, 7.964057e-06, 7.964059e-06, 7.964042e-06, 
    7.964049e-06, 7.964032e-06, 7.964037e-06, 7.964029e-06, 7.964033e-06, 
    7.964033e-06, 7.964038e-06, 7.964041e-06, 7.964049e-06, 7.964054e-06, 
    7.964059e-06, 7.964058e-06, 7.964052e-06, 7.964043e-06, 7.964034e-06, 
    7.964037e-06, 7.964029e-06, 7.964047e-06, 7.964039e-06, 7.964042e-06, 
    7.964035e-06, 7.964051e-06, 7.964038e-06, 7.964055e-06, 7.964053e-06, 
    7.964049e-06, 7.964039e-06, 7.964038e-06, 7.964035e-06, 7.964037e-06, 
    7.964043e-06, 7.964044e-06, 7.964049e-06, 7.964049e-06, 7.964053e-06, 
    7.964057e-06, 7.964054e-06, 7.964051e-06, 7.964043e-06, 7.964036e-06, 
    7.964028e-06, 7.964026e-06, 7.964017e-06, 7.964024e-06, 7.964012e-06, 
    7.964022e-06, 7.964005e-06, 7.964037e-06, 7.964023e-06, 7.964049e-06, 
    7.964046e-06, 7.96404e-06, 7.964029e-06, 7.964036e-06, 7.964029e-06, 
    7.964044e-06, 7.964052e-06, 7.964054e-06, 7.964059e-06, 7.964054e-06, 
    7.964055e-06, 7.96405e-06, 7.964052e-06, 7.964043e-06, 7.964048e-06, 
    7.964033e-06, 7.964029e-06, 7.964014e-06, 7.964005e-06, 7.963996e-06, 
    7.963991e-06, 7.96399e-06, 7.963989e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.604594e-14, 5.619708e-14, 5.616772e-14, 5.628951e-14, 5.622197e-14, 
    5.630169e-14, 5.607661e-14, 5.620306e-14, 5.612236e-14, 5.605958e-14, 
    5.65255e-14, 5.629494e-14, 5.676479e-14, 5.6618e-14, 5.698647e-14, 
    5.674193e-14, 5.703574e-14, 5.697947e-14, 5.714888e-14, 5.710037e-14, 
    5.731673e-14, 5.717126e-14, 5.742883e-14, 5.728203e-14, 5.730499e-14, 
    5.716645e-14, 5.634141e-14, 5.649681e-14, 5.633219e-14, 5.635437e-14, 
    5.634442e-14, 5.622336e-14, 5.616228e-14, 5.603441e-14, 5.605764e-14, 
    5.615157e-14, 5.636433e-14, 5.629217e-14, 5.647405e-14, 5.646995e-14, 
    5.667214e-14, 5.658101e-14, 5.692041e-14, 5.682406e-14, 5.710239e-14, 
    5.703244e-14, 5.70991e-14, 5.707889e-14, 5.709937e-14, 5.699675e-14, 
    5.704072e-14, 5.69504e-14, 5.659807e-14, 5.670171e-14, 5.639237e-14, 
    5.620598e-14, 5.608215e-14, 5.599419e-14, 5.600663e-14, 5.603033e-14, 
    5.615211e-14, 5.626657e-14, 5.635372e-14, 5.641197e-14, 5.646936e-14, 
    5.66428e-14, 5.673461e-14, 5.693987e-14, 5.690288e-14, 5.696556e-14, 
    5.702548e-14, 5.712595e-14, 5.710942e-14, 5.715366e-14, 5.696393e-14, 
    5.709004e-14, 5.68818e-14, 5.693878e-14, 5.648481e-14, 5.631165e-14, 
    5.623786e-14, 5.617335e-14, 5.601619e-14, 5.612474e-14, 5.608195e-14, 
    5.618375e-14, 5.624837e-14, 5.621642e-14, 5.641357e-14, 5.633695e-14, 
    5.674005e-14, 5.656656e-14, 5.701849e-14, 5.691048e-14, 5.704437e-14, 
    5.697607e-14, 5.709306e-14, 5.698777e-14, 5.717014e-14, 5.720979e-14, 
    5.718269e-14, 5.728683e-14, 5.698193e-14, 5.709909e-14, 5.621552e-14, 
    5.622073e-14, 5.624502e-14, 5.613821e-14, 5.613168e-14, 5.603377e-14, 
    5.612091e-14, 5.615799e-14, 5.625213e-14, 5.630776e-14, 5.636063e-14, 
    5.647682e-14, 5.660643e-14, 5.678752e-14, 5.691748e-14, 5.700454e-14, 
    5.695117e-14, 5.699828e-14, 5.694561e-14, 5.692092e-14, 5.719492e-14, 
    5.704112e-14, 5.727185e-14, 5.72591e-14, 5.715471e-14, 5.726054e-14, 
    5.622439e-14, 5.61944e-14, 5.609017e-14, 5.617174e-14, 5.60231e-14, 
    5.61063e-14, 5.615411e-14, 5.633852e-14, 5.637904e-14, 5.641655e-14, 
    5.649065e-14, 5.658567e-14, 5.67522e-14, 5.689693e-14, 5.702897e-14, 
    5.70193e-14, 5.70227e-14, 5.705216e-14, 5.697915e-14, 5.706415e-14, 
    5.70784e-14, 5.704112e-14, 5.725739e-14, 5.719564e-14, 5.725883e-14, 
    5.721863e-14, 5.620415e-14, 5.625462e-14, 5.622735e-14, 5.627862e-14, 
    5.624249e-14, 5.640303e-14, 5.645112e-14, 5.667601e-14, 5.65838e-14, 
    5.673057e-14, 5.659872e-14, 5.662209e-14, 5.673528e-14, 5.660586e-14, 
    5.688892e-14, 5.669703e-14, 5.705331e-14, 5.686185e-14, 5.70653e-14, 
    5.70284e-14, 5.708951e-14, 5.71442e-14, 5.7213e-14, 5.733981e-14, 
    5.731047e-14, 5.741647e-14, 5.632984e-14, 5.639522e-14, 5.638949e-14, 
    5.645791e-14, 5.650848e-14, 5.661806e-14, 5.679361e-14, 5.672763e-14, 
    5.684876e-14, 5.687302e-14, 5.668904e-14, 5.680202e-14, 5.643898e-14, 
    5.649767e-14, 5.646276e-14, 5.633498e-14, 5.674279e-14, 5.653363e-14, 
    5.691962e-14, 5.680653e-14, 5.71364e-14, 5.69724e-14, 5.72943e-14, 
    5.74316e-14, 5.756084e-14, 5.771153e-14, 5.643092e-14, 5.638651e-14, 
    5.646605e-14, 5.657598e-14, 5.667798e-14, 5.681343e-14, 5.682729e-14, 
    5.685264e-14, 5.691828e-14, 5.697346e-14, 5.686062e-14, 5.69873e-14, 
    5.651122e-14, 5.676095e-14, 5.636968e-14, 5.648758e-14, 5.656952e-14, 
    5.653361e-14, 5.672009e-14, 5.6764e-14, 5.694224e-14, 5.685016e-14, 
    5.73977e-14, 5.71557e-14, 5.782627e-14, 5.763919e-14, 5.637098e-14, 
    5.643079e-14, 5.663869e-14, 5.653981e-14, 5.682248e-14, 5.689192e-14, 
    5.69484e-14, 5.702052e-14, 5.702833e-14, 5.707104e-14, 5.700104e-14, 
    5.706829e-14, 5.681371e-14, 5.692753e-14, 5.661498e-14, 5.66911e-14, 
    5.66561e-14, 5.661767e-14, 5.673624e-14, 5.686237e-14, 5.686511e-14, 
    5.690553e-14, 5.701928e-14, 5.682362e-14, 5.742881e-14, 5.705527e-14, 
    5.649597e-14, 5.661098e-14, 5.662745e-14, 5.658291e-14, 5.688496e-14, 
    5.67756e-14, 5.707001e-14, 5.69905e-14, 5.712076e-14, 5.705604e-14, 
    5.704652e-14, 5.696337e-14, 5.691155e-14, 5.678061e-14, 5.667397e-14, 
    5.658937e-14, 5.660905e-14, 5.670197e-14, 5.687009e-14, 5.702901e-14, 
    5.699421e-14, 5.711086e-14, 5.6802e-14, 5.693155e-14, 5.688147e-14, 
    5.701203e-14, 5.672586e-14, 5.696944e-14, 5.666351e-14, 5.669037e-14, 
    5.677343e-14, 5.694031e-14, 5.697728e-14, 5.701665e-14, 5.699237e-14, 
    5.687437e-14, 5.685507e-14, 5.677142e-14, 5.67483e-14, 5.668453e-14, 
    5.663169e-14, 5.667996e-14, 5.673061e-14, 5.687443e-14, 5.700391e-14, 
    5.714497e-14, 5.717948e-14, 5.734394e-14, 5.721001e-14, 5.743088e-14, 
    5.724302e-14, 5.756809e-14, 5.698362e-14, 5.723759e-14, 5.677722e-14, 
    5.682691e-14, 5.691665e-14, 5.712242e-14, 5.701142e-14, 5.714126e-14, 
    5.685432e-14, 5.670515e-14, 5.666659e-14, 5.659451e-14, 5.666823e-14, 
    5.666224e-14, 5.673275e-14, 5.67101e-14, 5.687921e-14, 5.678841e-14, 
    5.704627e-14, 5.714024e-14, 5.740535e-14, 5.756758e-14, 5.77326e-14, 
    5.780536e-14, 5.78275e-14, 5.783675e-14 ;

 LITTERC =
  6.210302e-05, 6.210287e-05, 6.21029e-05, 6.210276e-05, 6.210284e-05, 
    6.210276e-05, 6.210299e-05, 6.210286e-05, 6.210294e-05, 6.2103e-05, 
    6.210252e-05, 6.210276e-05, 6.210227e-05, 6.210242e-05, 6.210204e-05, 
    6.21023e-05, 6.210199e-05, 6.210204e-05, 6.210187e-05, 6.210192e-05, 
    6.21017e-05, 6.210185e-05, 6.210158e-05, 6.210173e-05, 6.210171e-05, 
    6.210186e-05, 6.210271e-05, 6.210255e-05, 6.210272e-05, 6.21027e-05, 
    6.210271e-05, 6.210284e-05, 6.21029e-05, 6.210303e-05, 6.210301e-05, 
    6.210291e-05, 6.210269e-05, 6.210276e-05, 6.210258e-05, 6.210258e-05, 
    6.210237e-05, 6.210247e-05, 6.210211e-05, 6.210221e-05, 6.210192e-05, 
    6.210199e-05, 6.210192e-05, 6.210194e-05, 6.210192e-05, 6.210203e-05, 
    6.210199e-05, 6.210208e-05, 6.210244e-05, 6.210234e-05, 6.210266e-05, 
    6.210285e-05, 6.210298e-05, 6.210308e-05, 6.210306e-05, 6.210304e-05, 
    6.210291e-05, 6.210279e-05, 6.21027e-05, 6.210264e-05, 6.210258e-05, 
    6.21024e-05, 6.210231e-05, 6.210209e-05, 6.210212e-05, 6.210206e-05, 
    6.2102e-05, 6.21019e-05, 6.210191e-05, 6.210187e-05, 6.210207e-05, 
    6.210194e-05, 6.210215e-05, 6.210209e-05, 6.210256e-05, 6.210274e-05, 
    6.210282e-05, 6.210289e-05, 6.210306e-05, 6.210294e-05, 6.210298e-05, 
    6.210288e-05, 6.210281e-05, 6.210284e-05, 6.210264e-05, 6.210272e-05, 
    6.21023e-05, 6.210248e-05, 6.210201e-05, 6.210212e-05, 6.210198e-05, 
    6.210205e-05, 6.210193e-05, 6.210204e-05, 6.210185e-05, 6.21018e-05, 
    6.210183e-05, 6.210172e-05, 6.210204e-05, 6.210192e-05, 6.210284e-05, 
    6.210284e-05, 6.210282e-05, 6.210292e-05, 6.210293e-05, 6.210303e-05, 
    6.210295e-05, 6.21029e-05, 6.210281e-05, 6.210275e-05, 6.210269e-05, 
    6.210258e-05, 6.210244e-05, 6.210225e-05, 6.210211e-05, 6.210202e-05, 
    6.210208e-05, 6.210203e-05, 6.210208e-05, 6.210211e-05, 6.210183e-05, 
    6.210199e-05, 6.210175e-05, 6.210175e-05, 6.210186e-05, 6.210175e-05, 
    6.210284e-05, 6.210287e-05, 6.210298e-05, 6.210289e-05, 6.210305e-05, 
    6.210296e-05, 6.210291e-05, 6.210271e-05, 6.210268e-05, 6.210263e-05, 
    6.210256e-05, 6.210246e-05, 6.210228e-05, 6.210213e-05, 6.210199e-05, 
    6.210201e-05, 6.2102e-05, 6.210197e-05, 6.210205e-05, 6.210196e-05, 
    6.210194e-05, 6.210199e-05, 6.210176e-05, 6.210183e-05, 6.210175e-05, 
    6.21018e-05, 6.210286e-05, 6.21028e-05, 6.210283e-05, 6.210278e-05, 
    6.210282e-05, 6.210265e-05, 6.21026e-05, 6.210236e-05, 6.210246e-05, 
    6.210231e-05, 6.210244e-05, 6.210242e-05, 6.21023e-05, 6.210244e-05, 
    6.210214e-05, 6.210234e-05, 6.210197e-05, 6.210217e-05, 6.210196e-05, 
    6.210199e-05, 6.210194e-05, 6.210188e-05, 6.21018e-05, 6.210167e-05, 
    6.21017e-05, 6.210159e-05, 6.210273e-05, 6.210266e-05, 6.210266e-05, 
    6.210259e-05, 6.210254e-05, 6.210242e-05, 6.210224e-05, 6.210231e-05, 
    6.210218e-05, 6.210216e-05, 6.210235e-05, 6.210223e-05, 6.210261e-05, 
    6.210255e-05, 6.210259e-05, 6.210272e-05, 6.210229e-05, 6.210251e-05, 
    6.210211e-05, 6.210223e-05, 6.210188e-05, 6.210206e-05, 6.210172e-05, 
    6.210158e-05, 6.210144e-05, 6.210129e-05, 6.210262e-05, 6.210266e-05, 
    6.210258e-05, 6.210247e-05, 6.210236e-05, 6.210222e-05, 6.21022e-05, 
    6.210218e-05, 6.210211e-05, 6.210205e-05, 6.210218e-05, 6.210204e-05, 
    6.210254e-05, 6.210228e-05, 6.210268e-05, 6.210256e-05, 6.210247e-05, 
    6.210251e-05, 6.210232e-05, 6.210227e-05, 6.210209e-05, 6.210218e-05, 
    6.210162e-05, 6.210186e-05, 6.210116e-05, 6.210136e-05, 6.210268e-05, 
    6.210262e-05, 6.21024e-05, 6.210251e-05, 6.210221e-05, 6.210214e-05, 
    6.210208e-05, 6.210201e-05, 6.210199e-05, 6.210195e-05, 6.210202e-05, 
    6.210196e-05, 6.210222e-05, 6.21021e-05, 6.210243e-05, 6.210235e-05, 
    6.210239e-05, 6.210242e-05, 6.21023e-05, 6.210217e-05, 6.210217e-05, 
    6.210212e-05, 6.210201e-05, 6.210221e-05, 6.210158e-05, 6.210197e-05, 
    6.210255e-05, 6.210243e-05, 6.210242e-05, 6.210246e-05, 6.210215e-05, 
    6.210226e-05, 6.210196e-05, 6.210204e-05, 6.21019e-05, 6.210197e-05, 
    6.210198e-05, 6.210207e-05, 6.210212e-05, 6.210226e-05, 6.210236e-05, 
    6.210245e-05, 6.210244e-05, 6.210234e-05, 6.210216e-05, 6.210199e-05, 
    6.210203e-05, 6.210191e-05, 6.210223e-05, 6.21021e-05, 6.210215e-05, 
    6.210202e-05, 6.210231e-05, 6.210206e-05, 6.210238e-05, 6.210235e-05, 
    6.210226e-05, 6.210209e-05, 6.210205e-05, 6.210201e-05, 6.210204e-05, 
    6.210216e-05, 6.210218e-05, 6.210226e-05, 6.210229e-05, 6.210236e-05, 
    6.210241e-05, 6.210236e-05, 6.210231e-05, 6.210216e-05, 6.210202e-05, 
    6.210188e-05, 6.210184e-05, 6.210167e-05, 6.21018e-05, 6.210158e-05, 
    6.210178e-05, 6.210143e-05, 6.210204e-05, 6.210178e-05, 6.210226e-05, 
    6.21022e-05, 6.210211e-05, 6.21019e-05, 6.210202e-05, 6.210188e-05, 
    6.210218e-05, 6.210234e-05, 6.210237e-05, 6.210245e-05, 6.210237e-05, 
    6.210238e-05, 6.210231e-05, 6.210233e-05, 6.210215e-05, 6.210225e-05, 
    6.210198e-05, 6.210188e-05, 6.21016e-05, 6.210143e-05, 6.210127e-05, 
    6.210119e-05, 6.210116e-05, 6.210116e-05 ;

 LITTERC_HR =
  9.042218e-13, 9.066582e-13, 9.06185e-13, 9.081482e-13, 9.070596e-13, 
    9.083447e-13, 9.047163e-13, 9.067546e-13, 9.054538e-13, 9.044417e-13, 
    9.119526e-13, 9.082358e-13, 9.158099e-13, 9.134437e-13, 9.193833e-13, 
    9.154413e-13, 9.201776e-13, 9.192704e-13, 9.220014e-13, 9.212194e-13, 
    9.247071e-13, 9.223622e-13, 9.265142e-13, 9.241478e-13, 9.245178e-13, 
    9.222847e-13, 9.08985e-13, 9.1149e-13, 9.088363e-13, 9.091937e-13, 
    9.090335e-13, 9.070819e-13, 9.060972e-13, 9.04036e-13, 9.044105e-13, 
    9.059246e-13, 9.093545e-13, 9.081912e-13, 9.111232e-13, 9.11057e-13, 
    9.143163e-13, 9.128474e-13, 9.183185e-13, 9.167654e-13, 9.212521e-13, 
    9.201243e-13, 9.21199e-13, 9.208733e-13, 9.212032e-13, 9.195491e-13, 
    9.202579e-13, 9.18802e-13, 9.131223e-13, 9.14793e-13, 9.098064e-13, 
    9.068017e-13, 9.048056e-13, 9.033876e-13, 9.035881e-13, 9.039702e-13, 
    9.059335e-13, 9.077785e-13, 9.091833e-13, 9.101225e-13, 9.110475e-13, 
    9.138434e-13, 9.153234e-13, 9.186321e-13, 9.180359e-13, 9.190463e-13, 
    9.200121e-13, 9.216318e-13, 9.213653e-13, 9.220785e-13, 9.190202e-13, 
    9.210529e-13, 9.17696e-13, 9.186147e-13, 9.112964e-13, 9.085052e-13, 
    9.073157e-13, 9.062758e-13, 9.037423e-13, 9.05492e-13, 9.048023e-13, 
    9.064434e-13, 9.074851e-13, 9.0697e-13, 9.101482e-13, 9.08913e-13, 
    9.154111e-13, 9.126145e-13, 9.198995e-13, 9.181583e-13, 9.203168e-13, 
    9.192158e-13, 9.211016e-13, 9.194044e-13, 9.22344e-13, 9.229834e-13, 
    9.225464e-13, 9.242251e-13, 9.193102e-13, 9.211988e-13, 9.069555e-13, 
    9.070395e-13, 9.074311e-13, 9.057092e-13, 9.05604e-13, 9.040256e-13, 
    9.054304e-13, 9.060281e-13, 9.075457e-13, 9.084425e-13, 9.092948e-13, 
    9.111677e-13, 9.132571e-13, 9.161764e-13, 9.182712e-13, 9.196746e-13, 
    9.188143e-13, 9.195738e-13, 9.187247e-13, 9.183267e-13, 9.227437e-13, 
    9.202643e-13, 9.239838e-13, 9.237782e-13, 9.220953e-13, 9.238014e-13, 
    9.070985e-13, 9.06615e-13, 9.049348e-13, 9.062498e-13, 9.038537e-13, 
    9.051949e-13, 9.059656e-13, 9.089383e-13, 9.095915e-13, 9.101963e-13, 
    9.113908e-13, 9.129225e-13, 9.156069e-13, 9.1794e-13, 9.200684e-13, 
    9.199126e-13, 9.199674e-13, 9.204423e-13, 9.192653e-13, 9.206355e-13, 
    9.208652e-13, 9.202643e-13, 9.237507e-13, 9.227553e-13, 9.237739e-13, 
    9.231258e-13, 9.067723e-13, 9.075858e-13, 9.071462e-13, 9.079726e-13, 
    9.073903e-13, 9.099781e-13, 9.107536e-13, 9.143787e-13, 9.128923e-13, 
    9.152582e-13, 9.131329e-13, 9.135095e-13, 9.153342e-13, 9.13248e-13, 
    9.178109e-13, 9.147175e-13, 9.204609e-13, 9.173745e-13, 9.206541e-13, 
    9.200592e-13, 9.210443e-13, 9.219259e-13, 9.23035e-13, 9.250792e-13, 
    9.246061e-13, 9.26315e-13, 9.087983e-13, 9.098524e-13, 9.0976e-13, 
    9.10863e-13, 9.116782e-13, 9.134447e-13, 9.162744e-13, 9.152108e-13, 
    9.171635e-13, 9.175547e-13, 9.145887e-13, 9.164101e-13, 9.105579e-13, 
    9.115039e-13, 9.10941e-13, 9.088812e-13, 9.154553e-13, 9.120836e-13, 
    9.183058e-13, 9.164827e-13, 9.218002e-13, 9.191566e-13, 9.243456e-13, 
    9.265587e-13, 9.28642e-13, 9.310713e-13, 9.10428e-13, 9.097119e-13, 
    9.109943e-13, 9.127663e-13, 9.144105e-13, 9.165938e-13, 9.168174e-13, 
    9.17226e-13, 9.182842e-13, 9.191737e-13, 9.173547e-13, 9.193967e-13, 
    9.117223e-13, 9.157479e-13, 9.094407e-13, 9.113412e-13, 9.12662e-13, 
    9.120832e-13, 9.150894e-13, 9.157972e-13, 9.186703e-13, 9.17186e-13, 
    9.260123e-13, 9.221113e-13, 9.329207e-13, 9.299051e-13, 9.094616e-13, 
    9.104257e-13, 9.137772e-13, 9.121832e-13, 9.167398e-13, 9.178593e-13, 
    9.187697e-13, 9.199323e-13, 9.200581e-13, 9.207467e-13, 9.196182e-13, 
    9.207023e-13, 9.165985e-13, 9.184332e-13, 9.133949e-13, 9.14622e-13, 
    9.140578e-13, 9.134383e-13, 9.153496e-13, 9.173828e-13, 9.174271e-13, 
    9.180785e-13, 9.199124e-13, 9.167583e-13, 9.265139e-13, 9.204924e-13, 
    9.114765e-13, 9.133304e-13, 9.13596e-13, 9.12878e-13, 9.17747e-13, 
    9.159842e-13, 9.2073e-13, 9.194484e-13, 9.215481e-13, 9.205049e-13, 
    9.203514e-13, 9.190109e-13, 9.181757e-13, 9.16065e-13, 9.143459e-13, 
    9.129821e-13, 9.132994e-13, 9.147972e-13, 9.175073e-13, 9.200693e-13, 
    9.195082e-13, 9.213886e-13, 9.164097e-13, 9.184981e-13, 9.176907e-13, 
    9.197955e-13, 9.151824e-13, 9.19109e-13, 9.141773e-13, 9.146103e-13, 
    9.159492e-13, 9.186392e-13, 9.192352e-13, 9.1987e-13, 9.194785e-13, 
    9.175762e-13, 9.172653e-13, 9.159169e-13, 9.15544e-13, 9.145161e-13, 
    9.136643e-13, 9.144423e-13, 9.15259e-13, 9.175773e-13, 9.196646e-13, 
    9.219383e-13, 9.224947e-13, 9.251457e-13, 9.229868e-13, 9.265471e-13, 
    9.23519e-13, 9.287591e-13, 9.193374e-13, 9.234315e-13, 9.160103e-13, 
    9.168112e-13, 9.182579e-13, 9.21575e-13, 9.197856e-13, 9.218786e-13, 
    9.172531e-13, 9.148484e-13, 9.142268e-13, 9.13065e-13, 9.142534e-13, 
    9.141568e-13, 9.152933e-13, 9.149282e-13, 9.176543e-13, 9.161906e-13, 
    9.203472e-13, 9.218622e-13, 9.261357e-13, 9.287508e-13, 9.314109e-13, 
    9.325837e-13, 9.329406e-13, 9.330898e-13 ;

 LITTERC_LOSS =
  1.67461e-12, 1.679122e-12, 1.678246e-12, 1.681882e-12, 1.679866e-12, 
    1.682246e-12, 1.675526e-12, 1.679301e-12, 1.676892e-12, 1.675017e-12, 
    1.688928e-12, 1.682044e-12, 1.696071e-12, 1.691689e-12, 1.70269e-12, 
    1.695389e-12, 1.70416e-12, 1.70248e-12, 1.707538e-12, 1.70609e-12, 
    1.712549e-12, 1.708206e-12, 1.715896e-12, 1.711514e-12, 1.712199e-12, 
    1.708063e-12, 1.683432e-12, 1.688071e-12, 1.683156e-12, 1.683818e-12, 
    1.683522e-12, 1.679907e-12, 1.678084e-12, 1.674266e-12, 1.67496e-12, 
    1.677764e-12, 1.684116e-12, 1.681962e-12, 1.687392e-12, 1.687269e-12, 
    1.693305e-12, 1.690585e-12, 1.700717e-12, 1.697841e-12, 1.706151e-12, 
    1.704062e-12, 1.706052e-12, 1.705449e-12, 1.70606e-12, 1.702996e-12, 
    1.704309e-12, 1.701613e-12, 1.691094e-12, 1.694188e-12, 1.684953e-12, 
    1.679388e-12, 1.675691e-12, 1.673065e-12, 1.673437e-12, 1.674144e-12, 
    1.67778e-12, 1.681197e-12, 1.683799e-12, 1.685538e-12, 1.687251e-12, 
    1.69243e-12, 1.695171e-12, 1.701298e-12, 1.700194e-12, 1.702065e-12, 
    1.703854e-12, 1.706854e-12, 1.70636e-12, 1.707681e-12, 1.702017e-12, 
    1.705782e-12, 1.699565e-12, 1.701266e-12, 1.687713e-12, 1.682543e-12, 
    1.68034e-12, 1.678414e-12, 1.673722e-12, 1.676963e-12, 1.675685e-12, 
    1.678725e-12, 1.680654e-12, 1.6797e-12, 1.685586e-12, 1.683298e-12, 
    1.695333e-12, 1.690154e-12, 1.703646e-12, 1.700421e-12, 1.704418e-12, 
    1.702379e-12, 1.705872e-12, 1.702729e-12, 1.708173e-12, 1.709357e-12, 
    1.708548e-12, 1.711657e-12, 1.702554e-12, 1.706052e-12, 1.679673e-12, 
    1.679829e-12, 1.680554e-12, 1.677365e-12, 1.67717e-12, 1.674247e-12, 
    1.676848e-12, 1.677955e-12, 1.680766e-12, 1.682427e-12, 1.684005e-12, 
    1.687474e-12, 1.691344e-12, 1.69675e-12, 1.70063e-12, 1.703229e-12, 
    1.701636e-12, 1.703042e-12, 1.70147e-12, 1.700733e-12, 1.708913e-12, 
    1.704321e-12, 1.71121e-12, 1.710829e-12, 1.707712e-12, 1.710872e-12, 
    1.679938e-12, 1.679042e-12, 1.675931e-12, 1.678366e-12, 1.673928e-12, 
    1.676412e-12, 1.67784e-12, 1.683345e-12, 1.684555e-12, 1.685675e-12, 
    1.687887e-12, 1.690724e-12, 1.695696e-12, 1.700016e-12, 1.703958e-12, 
    1.70367e-12, 1.703771e-12, 1.704651e-12, 1.702471e-12, 1.705009e-12, 
    1.705434e-12, 1.704321e-12, 1.710778e-12, 1.708934e-12, 1.710821e-12, 
    1.709621e-12, 1.679334e-12, 1.68084e-12, 1.680026e-12, 1.681557e-12, 
    1.680478e-12, 1.685271e-12, 1.686707e-12, 1.693421e-12, 1.690668e-12, 
    1.69505e-12, 1.691114e-12, 1.691811e-12, 1.695191e-12, 1.691327e-12, 
    1.699777e-12, 1.694048e-12, 1.704685e-12, 1.698969e-12, 1.705043e-12, 
    1.703941e-12, 1.705766e-12, 1.707398e-12, 1.709453e-12, 1.713238e-12, 
    1.712362e-12, 1.715527e-12, 1.683086e-12, 1.685038e-12, 1.684867e-12, 
    1.68691e-12, 1.688419e-12, 1.691691e-12, 1.696932e-12, 1.694962e-12, 
    1.698578e-12, 1.699303e-12, 1.69381e-12, 1.697183e-12, 1.686345e-12, 
    1.688097e-12, 1.687054e-12, 1.683239e-12, 1.695415e-12, 1.68917e-12, 
    1.700694e-12, 1.697318e-12, 1.707166e-12, 1.70227e-12, 1.71188e-12, 
    1.715979e-12, 1.719837e-12, 1.724336e-12, 1.686104e-12, 1.684778e-12, 
    1.687153e-12, 1.690435e-12, 1.69348e-12, 1.697524e-12, 1.697937e-12, 
    1.698694e-12, 1.700654e-12, 1.702301e-12, 1.698933e-12, 1.702714e-12, 
    1.688501e-12, 1.695957e-12, 1.684276e-12, 1.687796e-12, 1.690242e-12, 
    1.68917e-12, 1.694737e-12, 1.696048e-12, 1.701369e-12, 1.69862e-12, 
    1.714967e-12, 1.707742e-12, 1.727761e-12, 1.722176e-12, 1.684314e-12, 
    1.6861e-12, 1.692307e-12, 1.689355e-12, 1.697794e-12, 1.699867e-12, 
    1.701553e-12, 1.703706e-12, 1.703939e-12, 1.705215e-12, 1.703125e-12, 
    1.705132e-12, 1.697532e-12, 1.70093e-12, 1.691599e-12, 1.693872e-12, 
    1.692827e-12, 1.691679e-12, 1.695219e-12, 1.698985e-12, 1.699066e-12, 
    1.700273e-12, 1.703669e-12, 1.697828e-12, 1.715895e-12, 1.704744e-12, 
    1.688046e-12, 1.691479e-12, 1.691971e-12, 1.690641e-12, 1.699659e-12, 
    1.696394e-12, 1.705184e-12, 1.70281e-12, 1.706699e-12, 1.704767e-12, 
    1.704482e-12, 1.702e-12, 1.700453e-12, 1.696544e-12, 1.69336e-12, 
    1.690835e-12, 1.691422e-12, 1.694196e-12, 1.699215e-12, 1.70396e-12, 
    1.702921e-12, 1.706403e-12, 1.697182e-12, 1.70105e-12, 1.699555e-12, 
    1.703453e-12, 1.694909e-12, 1.702181e-12, 1.693048e-12, 1.69385e-12, 
    1.696329e-12, 1.701312e-12, 1.702415e-12, 1.703591e-12, 1.702866e-12, 
    1.699343e-12, 1.698767e-12, 1.69627e-12, 1.695579e-12, 1.693675e-12, 
    1.692098e-12, 1.693539e-12, 1.695051e-12, 1.699345e-12, 1.70321e-12, 
    1.707422e-12, 1.708452e-12, 1.713362e-12, 1.709363e-12, 1.715957e-12, 
    1.710349e-12, 1.720054e-12, 1.702605e-12, 1.710187e-12, 1.696443e-12, 
    1.697926e-12, 1.700605e-12, 1.706749e-12, 1.703435e-12, 1.707311e-12, 
    1.698744e-12, 1.694291e-12, 1.69314e-12, 1.690988e-12, 1.693189e-12, 
    1.69301e-12, 1.695115e-12, 1.694439e-12, 1.699487e-12, 1.696777e-12, 
    1.704475e-12, 1.70728e-12, 1.715195e-12, 1.720038e-12, 1.724965e-12, 
    1.727137e-12, 1.727798e-12, 1.728074e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  4.221994e-18, 4.220502e-18, 4.220785e-18, 4.219598e-18, 4.220246e-18, 
    4.219477e-18, 4.221678e-18, 4.220454e-18, 4.221228e-18, 4.221842e-18, 
    4.217337e-18, 4.219542e-18, 4.214933e-18, 4.216355e-18, 4.212751e-18, 
    4.21517e-18, 4.212259e-18, 4.212792e-18, 4.211119e-18, 4.211596e-18, 
    4.209518e-18, 4.210898e-18, 4.208397e-18, 4.209832e-18, 4.209618e-18, 
    4.210948e-18, 4.219071e-18, 4.21762e-18, 4.219163e-18, 4.218954e-18, 
    4.219042e-18, 4.220242e-18, 4.220866e-18, 4.222088e-18, 4.221861e-18, 
    4.220953e-18, 4.21886e-18, 4.219551e-18, 4.217756e-18, 4.217795e-18, 
    4.215819e-18, 4.21671e-18, 4.213374e-18, 4.214314e-18, 4.211576e-18, 
    4.212268e-18, 4.211613e-18, 4.211808e-18, 4.21161e-18, 4.212624e-18, 
    4.212191e-18, 4.213075e-18, 4.216549e-18, 4.215536e-18, 4.218576e-18, 
    4.220451e-18, 4.22163e-18, 4.222488e-18, 4.222367e-18, 4.222141e-18, 
    4.220948e-18, 4.219804e-18, 4.218941e-18, 4.218369e-18, 4.217801e-18, 
    4.216159e-18, 4.215229e-18, 4.213197e-18, 4.21354e-18, 4.212941e-18, 
    4.212335e-18, 4.211352e-18, 4.21151e-18, 4.211083e-18, 4.21294e-18, 
    4.211714e-18, 4.213741e-18, 4.213189e-18, 4.217743e-18, 4.21936e-18, 
    4.220131e-18, 4.220734e-18, 4.222275e-18, 4.221216e-18, 4.221635e-18, 
    4.220617e-18, 4.219984e-18, 4.220293e-18, 4.218353e-18, 4.21911e-18, 
    4.215175e-18, 4.216867e-18, 4.212406e-18, 4.213467e-18, 4.212148e-18, 
    4.212816e-18, 4.21168e-18, 4.212702e-18, 4.210916e-18, 4.210538e-18, 
    4.210798e-18, 4.209768e-18, 4.212762e-18, 4.211622e-18, 4.220307e-18, 
    4.220256e-18, 4.220014e-18, 4.221085e-18, 4.221145e-18, 4.222099e-18, 
    4.221242e-18, 4.220884e-18, 4.21994e-18, 4.2194e-18, 4.21888e-18, 
    4.217738e-18, 4.216479e-18, 4.214695e-18, 4.2134e-18, 4.212537e-18, 
    4.21306e-18, 4.212599e-18, 4.213118e-18, 4.213357e-18, 4.210686e-18, 
    4.212193e-18, 4.209916e-18, 4.210038e-18, 4.211076e-18, 4.210025e-18, 
    4.22022e-18, 4.22051e-18, 4.221547e-18, 4.220735e-18, 4.222202e-18, 
    4.221393e-18, 4.220934e-18, 4.219116e-18, 4.218694e-18, 4.218332e-18, 
    4.217597e-18, 4.216665e-18, 4.215039e-18, 4.213612e-18, 4.212297e-18, 
    4.212391e-18, 4.212359e-18, 4.212075e-18, 4.212791e-18, 4.211957e-18, 
    4.211825e-18, 4.212182e-18, 4.210056e-18, 4.210661e-18, 4.210041e-18, 
    4.210433e-18, 4.220413e-18, 4.219921e-18, 4.220189e-18, 4.219691e-18, 
    4.220049e-18, 4.218486e-18, 4.218018e-18, 4.215805e-18, 4.216689e-18, 
    4.215256e-18, 4.216536e-18, 4.216315e-18, 4.21525e-18, 4.21646e-18, 
    4.213708e-18, 4.215609e-18, 4.212064e-18, 4.213996e-18, 4.211945e-18, 
    4.212302e-18, 4.211701e-18, 4.211174e-18, 4.210492e-18, 4.209265e-18, 
    4.209545e-18, 4.208504e-18, 4.219179e-18, 4.218551e-18, 4.218589e-18, 
    4.217919e-18, 4.217428e-18, 4.216342e-18, 4.214624e-18, 4.215264e-18, 
    4.21407e-18, 4.213836e-18, 4.21564e-18, 4.214549e-18, 4.218117e-18, 
    4.217559e-18, 4.217878e-18, 4.21914e-18, 4.215141e-18, 4.217202e-18, 
    4.213382e-18, 4.214493e-18, 4.211251e-18, 4.21288e-18, 4.209703e-18, 
    4.208395e-18, 4.207082e-18, 4.205647e-18, 4.218189e-18, 4.218617e-18, 
    4.217834e-18, 4.216784e-18, 4.21576e-18, 4.214428e-18, 4.214282e-18, 
    4.214038e-18, 4.213384e-18, 4.212844e-18, 4.213978e-18, 4.212707e-18, 
    4.217465e-18, 4.214954e-18, 4.218796e-18, 4.217662e-18, 4.216838e-18, 
    4.217181e-18, 4.215333e-18, 4.214904e-18, 4.213169e-18, 4.214055e-18, 
    4.208733e-18, 4.211087e-18, 4.204497e-18, 4.206345e-18, 4.218772e-18, 
    4.218182e-18, 4.216158e-18, 4.217117e-18, 4.21433e-18, 4.213653e-18, 
    4.213087e-18, 4.212394e-18, 4.212306e-18, 4.211893e-18, 4.212572e-18, 
    4.211913e-18, 4.214425e-18, 4.213299e-18, 4.216367e-18, 4.21563e-18, 
    4.215963e-18, 4.216342e-18, 4.215176e-18, 4.213965e-18, 4.21391e-18, 
    4.213527e-18, 4.212499e-18, 4.214318e-18, 4.208482e-18, 4.212131e-18, 
    4.217541e-18, 4.216446e-18, 4.216255e-18, 4.216685e-18, 4.213721e-18, 
    4.214798e-18, 4.211899e-18, 4.212675e-18, 4.211396e-18, 4.212034e-18, 
    4.212129e-18, 4.212943e-18, 4.213457e-18, 4.214754e-18, 4.215802e-18, 
    4.216619e-18, 4.216426e-18, 4.215529e-18, 4.213883e-18, 4.212311e-18, 
    4.212659e-18, 4.211493e-18, 4.214532e-18, 4.213271e-18, 4.213768e-18, 
    4.212469e-18, 4.215287e-18, 4.212974e-18, 4.21589e-18, 4.215628e-18, 
    4.214819e-18, 4.213206e-18, 4.212806e-18, 4.212432e-18, 4.212657e-18, 
    4.213837e-18, 4.214018e-18, 4.214832e-18, 4.215071e-18, 4.215683e-18, 
    4.216203e-18, 4.215735e-18, 4.215249e-18, 4.213825e-18, 4.212558e-18, 
    4.21117e-18, 4.21082e-18, 4.209272e-18, 4.210571e-18, 4.208467e-18, 
    4.210314e-18, 4.20709e-18, 4.212797e-18, 4.210312e-18, 4.214773e-18, 
    4.214284e-18, 4.213431e-18, 4.211418e-18, 4.212474e-18, 4.211225e-18, 
    4.214023e-18, 4.215512e-18, 4.215862e-18, 4.216574e-18, 4.215846e-18, 
    4.215903e-18, 4.215209e-18, 4.21543e-18, 4.213777e-18, 4.214663e-18, 
    4.212139e-18, 4.211228e-18, 4.208623e-18, 4.207048e-18, 4.205401e-18, 
    4.20469e-18, 4.204471e-18, 4.204381e-18 ;

 MEG_acetic_acid =
  6.33299e-19, 6.330752e-19, 6.331177e-19, 6.329397e-19, 6.330368e-19, 
    6.329215e-19, 6.332517e-19, 6.330681e-19, 6.331842e-19, 6.332763e-19, 
    6.326004e-19, 6.329313e-19, 6.322399e-19, 6.324532e-19, 6.319126e-19, 
    6.322755e-19, 6.318388e-19, 6.319188e-19, 6.316678e-19, 6.317394e-19, 
    6.314276e-19, 6.316347e-19, 6.312595e-19, 6.314747e-19, 6.314427e-19, 
    6.316422e-19, 6.328606e-19, 6.326429e-19, 6.328745e-19, 6.328432e-19, 
    6.328563e-19, 6.330363e-19, 6.331299e-19, 6.333132e-19, 6.332791e-19, 
    6.331429e-19, 6.32829e-19, 6.329327e-19, 6.326634e-19, 6.326693e-19, 
    6.323729e-19, 6.325065e-19, 6.320061e-19, 6.321471e-19, 6.317363e-19, 
    6.318402e-19, 6.317419e-19, 6.317711e-19, 6.317416e-19, 6.318936e-19, 
    6.318287e-19, 6.319612e-19, 6.324823e-19, 6.323303e-19, 6.327864e-19, 
    6.330677e-19, 6.332444e-19, 6.333732e-19, 6.33355e-19, 6.333212e-19, 
    6.331422e-19, 6.329706e-19, 6.328412e-19, 6.327553e-19, 6.326702e-19, 
    6.324239e-19, 6.322844e-19, 6.319796e-19, 6.32031e-19, 6.319412e-19, 
    6.318503e-19, 6.317028e-19, 6.317265e-19, 6.316624e-19, 6.319409e-19, 
    6.31757e-19, 6.320611e-19, 6.319783e-19, 6.326614e-19, 6.32904e-19, 
    6.330197e-19, 6.331101e-19, 6.333413e-19, 6.331824e-19, 6.332453e-19, 
    6.330926e-19, 6.329976e-19, 6.33044e-19, 6.327529e-19, 6.328666e-19, 
    6.322762e-19, 6.3253e-19, 6.318609e-19, 6.320201e-19, 6.318223e-19, 
    6.319225e-19, 6.317519e-19, 6.319053e-19, 6.316374e-19, 6.315807e-19, 
    6.316197e-19, 6.314651e-19, 6.319142e-19, 6.317433e-19, 6.330459e-19, 
    6.330385e-19, 6.33002e-19, 6.331627e-19, 6.331718e-19, 6.333149e-19, 
    6.331862e-19, 6.331326e-19, 6.32991e-19, 6.3291e-19, 6.32832e-19, 
    6.326607e-19, 6.324719e-19, 6.322043e-19, 6.320099e-19, 6.318806e-19, 
    6.31959e-19, 6.318899e-19, 6.319676e-19, 6.320035e-19, 6.316029e-19, 
    6.318289e-19, 6.314874e-19, 6.315058e-19, 6.316614e-19, 6.315036e-19, 
    6.33033e-19, 6.330764e-19, 6.332321e-19, 6.331102e-19, 6.333303e-19, 
    6.332089e-19, 6.331402e-19, 6.328674e-19, 6.32804e-19, 6.327498e-19, 
    6.326395e-19, 6.324998e-19, 6.322559e-19, 6.320417e-19, 6.318444e-19, 
    6.318586e-19, 6.318537e-19, 6.318112e-19, 6.319186e-19, 6.317935e-19, 
    6.317738e-19, 6.318272e-19, 6.315083e-19, 6.315992e-19, 6.315062e-19, 
    6.31565e-19, 6.33062e-19, 6.329882e-19, 6.330282e-19, 6.329537e-19, 
    6.330073e-19, 6.327729e-19, 6.327027e-19, 6.323707e-19, 6.325033e-19, 
    6.322884e-19, 6.324803e-19, 6.324471e-19, 6.322874e-19, 6.32469e-19, 
    6.320562e-19, 6.323413e-19, 6.318095e-19, 6.320994e-19, 6.317917e-19, 
    6.318453e-19, 6.317552e-19, 6.31676e-19, 6.315738e-19, 6.313897e-19, 
    6.314317e-19, 6.312756e-19, 6.328769e-19, 6.327827e-19, 6.327883e-19, 
    6.326878e-19, 6.326142e-19, 6.324513e-19, 6.321936e-19, 6.322896e-19, 
    6.321105e-19, 6.320754e-19, 6.32346e-19, 6.321824e-19, 6.327175e-19, 
    6.326338e-19, 6.326817e-19, 6.32871e-19, 6.322712e-19, 6.325803e-19, 
    6.320072e-19, 6.321739e-19, 6.316876e-19, 6.319319e-19, 6.314555e-19, 
    6.312592e-19, 6.310623e-19, 6.30847e-19, 6.327283e-19, 6.327926e-19, 
    6.326751e-19, 6.325176e-19, 6.32364e-19, 6.321642e-19, 6.321423e-19, 
    6.321057e-19, 6.320076e-19, 6.319265e-19, 6.320967e-19, 6.31906e-19, 
    6.326197e-19, 6.322431e-19, 6.328194e-19, 6.326493e-19, 6.325257e-19, 
    6.325772e-19, 6.322999e-19, 6.322355e-19, 6.319753e-19, 6.321083e-19, 
    6.3131e-19, 6.31663e-19, 6.306744e-19, 6.309518e-19, 6.328158e-19, 
    6.327273e-19, 6.324236e-19, 6.325676e-19, 6.321495e-19, 6.320478e-19, 
    6.31963e-19, 6.31859e-19, 6.318458e-19, 6.317839e-19, 6.318857e-19, 
    6.317869e-19, 6.321638e-19, 6.319948e-19, 6.324551e-19, 6.323445e-19, 
    6.323945e-19, 6.324512e-19, 6.322764e-19, 6.320947e-19, 6.320864e-19, 
    6.32029e-19, 6.318748e-19, 6.321476e-19, 6.312723e-19, 6.318196e-19, 
    6.326311e-19, 6.324669e-19, 6.324382e-19, 6.325027e-19, 6.320582e-19, 
    6.322197e-19, 6.317848e-19, 6.319013e-19, 6.317094e-19, 6.318051e-19, 
    6.318194e-19, 6.319414e-19, 6.320186e-19, 6.322131e-19, 6.323702e-19, 
    6.324927e-19, 6.32464e-19, 6.323293e-19, 6.320825e-19, 6.318466e-19, 
    6.318988e-19, 6.317239e-19, 6.321799e-19, 6.319907e-19, 6.320651e-19, 
    6.318703e-19, 6.32293e-19, 6.31946e-19, 6.323835e-19, 6.323441e-19, 
    6.322228e-19, 6.319808e-19, 6.319209e-19, 6.318648e-19, 6.318985e-19, 
    6.320755e-19, 6.321027e-19, 6.322247e-19, 6.322606e-19, 6.323524e-19, 
    6.324304e-19, 6.323602e-19, 6.322873e-19, 6.320737e-19, 6.318837e-19, 
    6.316755e-19, 6.316229e-19, 6.313907e-19, 6.315855e-19, 6.312701e-19, 
    6.315471e-19, 6.310635e-19, 6.319195e-19, 6.315467e-19, 6.322158e-19, 
    6.321426e-19, 6.320147e-19, 6.317127e-19, 6.318711e-19, 6.316838e-19, 
    6.321034e-19, 6.323267e-19, 6.323793e-19, 6.324861e-19, 6.323768e-19, 
    6.323855e-19, 6.322813e-19, 6.323145e-19, 6.320665e-19, 6.321995e-19, 
    6.318209e-19, 6.316842e-19, 6.312934e-19, 6.310571e-19, 6.308101e-19, 
    6.307035e-19, 6.306706e-19, 6.306571e-19 ;

 MEG_acetone =
  1.325731e-16, 1.325484e-16, 1.325531e-16, 1.325334e-16, 1.325442e-16, 
    1.325314e-16, 1.325679e-16, 1.325476e-16, 1.325604e-16, 1.325706e-16, 
    1.32496e-16, 1.325325e-16, 1.324562e-16, 1.324798e-16, 1.324201e-16, 
    1.324602e-16, 1.32412e-16, 1.324208e-16, 1.323932e-16, 1.32401e-16, 
    1.323667e-16, 1.323895e-16, 1.323482e-16, 1.323719e-16, 1.323684e-16, 
    1.323903e-16, 1.325247e-16, 1.325007e-16, 1.325262e-16, 1.325228e-16, 
    1.325242e-16, 1.325441e-16, 1.325544e-16, 1.325747e-16, 1.325709e-16, 
    1.325559e-16, 1.325212e-16, 1.325327e-16, 1.32503e-16, 1.325036e-16, 
    1.324709e-16, 1.324857e-16, 1.324304e-16, 1.32446e-16, 1.324007e-16, 
    1.324121e-16, 1.324013e-16, 1.324045e-16, 1.324013e-16, 1.32418e-16, 
    1.324109e-16, 1.324255e-16, 1.32483e-16, 1.324662e-16, 1.325165e-16, 
    1.325476e-16, 1.325671e-16, 1.325813e-16, 1.325793e-16, 1.325755e-16, 
    1.325558e-16, 1.325368e-16, 1.325226e-16, 1.325131e-16, 1.325037e-16, 
    1.324765e-16, 1.324611e-16, 1.324275e-16, 1.324332e-16, 1.324233e-16, 
    1.324133e-16, 1.32397e-16, 1.323996e-16, 1.323926e-16, 1.324233e-16, 
    1.32403e-16, 1.324365e-16, 1.324274e-16, 1.325027e-16, 1.325295e-16, 
    1.325423e-16, 1.325522e-16, 1.325778e-16, 1.325602e-16, 1.325672e-16, 
    1.325503e-16, 1.325398e-16, 1.325449e-16, 1.325128e-16, 1.325254e-16, 
    1.324602e-16, 1.324882e-16, 1.324144e-16, 1.32432e-16, 1.324102e-16, 
    1.324212e-16, 1.324024e-16, 1.324193e-16, 1.323898e-16, 1.323836e-16, 
    1.323879e-16, 1.323708e-16, 1.324203e-16, 1.324015e-16, 1.325452e-16, 
    1.325443e-16, 1.325403e-16, 1.32558e-16, 1.325591e-16, 1.325749e-16, 
    1.325607e-16, 1.325547e-16, 1.325391e-16, 1.325302e-16, 1.325216e-16, 
    1.325027e-16, 1.324818e-16, 1.324523e-16, 1.324309e-16, 1.324166e-16, 
    1.324252e-16, 1.324176e-16, 1.324262e-16, 1.324301e-16, 1.32386e-16, 
    1.324109e-16, 1.323733e-16, 1.323753e-16, 1.323924e-16, 1.323751e-16, 
    1.325437e-16, 1.325485e-16, 1.325657e-16, 1.325523e-16, 1.325766e-16, 
    1.325632e-16, 1.325556e-16, 1.325255e-16, 1.325185e-16, 1.325125e-16, 
    1.325003e-16, 1.324849e-16, 1.32458e-16, 1.324344e-16, 1.324126e-16, 
    1.324142e-16, 1.324136e-16, 1.324089e-16, 1.324208e-16, 1.32407e-16, 
    1.324048e-16, 1.324107e-16, 1.323756e-16, 1.323856e-16, 1.323754e-16, 
    1.323818e-16, 1.325469e-16, 1.325388e-16, 1.325432e-16, 1.32535e-16, 
    1.325409e-16, 1.32515e-16, 1.325073e-16, 1.324707e-16, 1.324853e-16, 
    1.324616e-16, 1.324828e-16, 1.324791e-16, 1.324615e-16, 1.324815e-16, 
    1.32436e-16, 1.324674e-16, 1.324088e-16, 1.324407e-16, 1.324068e-16, 
    1.324127e-16, 1.324028e-16, 1.323941e-16, 1.323828e-16, 1.323625e-16, 
    1.323671e-16, 1.3235e-16, 1.325265e-16, 1.325161e-16, 1.325167e-16, 
    1.325057e-16, 1.324975e-16, 1.324796e-16, 1.324511e-16, 1.324617e-16, 
    1.32442e-16, 1.324381e-16, 1.324679e-16, 1.324499e-16, 1.325089e-16, 
    1.324997e-16, 1.32505e-16, 1.325259e-16, 1.324597e-16, 1.324938e-16, 
    1.324306e-16, 1.32449e-16, 1.323953e-16, 1.324223e-16, 1.323698e-16, 
    1.323482e-16, 1.323265e-16, 1.323028e-16, 1.325101e-16, 1.325172e-16, 
    1.325042e-16, 1.324869e-16, 1.324699e-16, 1.324479e-16, 1.324455e-16, 
    1.324414e-16, 1.324306e-16, 1.324217e-16, 1.324404e-16, 1.324194e-16, 
    1.324981e-16, 1.324566e-16, 1.325202e-16, 1.325014e-16, 1.324878e-16, 
    1.324934e-16, 1.324629e-16, 1.324558e-16, 1.32427e-16, 1.324417e-16, 
    1.323537e-16, 1.323926e-16, 1.322838e-16, 1.323143e-16, 1.325198e-16, 
    1.3251e-16, 1.324765e-16, 1.324924e-16, 1.324463e-16, 1.32435e-16, 
    1.324257e-16, 1.324142e-16, 1.324128e-16, 1.324059e-16, 1.324172e-16, 
    1.324063e-16, 1.324478e-16, 1.324292e-16, 1.3248e-16, 1.324678e-16, 
    1.324733e-16, 1.324796e-16, 1.324603e-16, 1.324402e-16, 1.324393e-16, 
    1.32433e-16, 1.32416e-16, 1.324461e-16, 1.323496e-16, 1.324099e-16, 
    1.324994e-16, 1.324813e-16, 1.324781e-16, 1.324852e-16, 1.324362e-16, 
    1.32454e-16, 1.32406e-16, 1.324189e-16, 1.323977e-16, 1.324083e-16, 
    1.324099e-16, 1.324233e-16, 1.324318e-16, 1.324533e-16, 1.324706e-16, 
    1.324841e-16, 1.32481e-16, 1.324661e-16, 1.324389e-16, 1.324128e-16, 
    1.324186e-16, 1.323993e-16, 1.324496e-16, 1.324287e-16, 1.324369e-16, 
    1.324155e-16, 1.324621e-16, 1.324238e-16, 1.324721e-16, 1.324677e-16, 
    1.324544e-16, 1.324276e-16, 1.32421e-16, 1.324148e-16, 1.324186e-16, 
    1.324381e-16, 1.324411e-16, 1.324546e-16, 1.324585e-16, 1.324686e-16, 
    1.324772e-16, 1.324695e-16, 1.324615e-16, 1.324379e-16, 1.324169e-16, 
    1.32394e-16, 1.323882e-16, 1.323626e-16, 1.323841e-16, 1.323493e-16, 
    1.323798e-16, 1.323266e-16, 1.324209e-16, 1.323798e-16, 1.324536e-16, 
    1.324455e-16, 1.324314e-16, 1.323981e-16, 1.324156e-16, 1.323949e-16, 
    1.324412e-16, 1.324658e-16, 1.324716e-16, 1.324834e-16, 1.324713e-16, 
    1.324723e-16, 1.324608e-16, 1.324645e-16, 1.324371e-16, 1.324518e-16, 
    1.3241e-16, 1.32395e-16, 1.323519e-16, 1.323259e-16, 1.322988e-16, 
    1.32287e-16, 1.322834e-16, 1.322819e-16 ;

 MEG_carene_3 =
  5.257811e-17, 5.256785e-17, 5.25698e-17, 5.256164e-17, 5.256609e-17, 
    5.25608e-17, 5.257595e-17, 5.256752e-17, 5.257285e-17, 5.257707e-17, 
    5.254608e-17, 5.256125e-17, 5.252955e-17, 5.253933e-17, 5.251455e-17, 
    5.253118e-17, 5.251117e-17, 5.251483e-17, 5.250334e-17, 5.250662e-17, 
    5.249234e-17, 5.250182e-17, 5.248465e-17, 5.24945e-17, 5.249303e-17, 
    5.250217e-17, 5.255801e-17, 5.254802e-17, 5.255865e-17, 5.255721e-17, 
    5.255781e-17, 5.256606e-17, 5.257036e-17, 5.257877e-17, 5.25772e-17, 
    5.257095e-17, 5.255656e-17, 5.256131e-17, 5.254896e-17, 5.254924e-17, 
    5.253565e-17, 5.254177e-17, 5.251883e-17, 5.25253e-17, 5.250648e-17, 
    5.251123e-17, 5.250673e-17, 5.250807e-17, 5.250672e-17, 5.251368e-17, 
    5.251071e-17, 5.251677e-17, 5.254067e-17, 5.25337e-17, 5.255461e-17, 
    5.25675e-17, 5.257561e-17, 5.258152e-17, 5.258069e-17, 5.257913e-17, 
    5.257092e-17, 5.256305e-17, 5.255712e-17, 5.255318e-17, 5.254928e-17, 
    5.253798e-17, 5.253159e-17, 5.251762e-17, 5.251997e-17, 5.251586e-17, 
    5.25117e-17, 5.250494e-17, 5.250603e-17, 5.250309e-17, 5.251584e-17, 
    5.250742e-17, 5.252135e-17, 5.251756e-17, 5.254887e-17, 5.256e-17, 
    5.25653e-17, 5.256945e-17, 5.258005e-17, 5.257276e-17, 5.257565e-17, 
    5.256865e-17, 5.256429e-17, 5.256642e-17, 5.255307e-17, 5.255828e-17, 
    5.253122e-17, 5.254285e-17, 5.251218e-17, 5.251947e-17, 5.251041e-17, 
    5.2515e-17, 5.250719e-17, 5.251422e-17, 5.250195e-17, 5.249935e-17, 
    5.250114e-17, 5.249406e-17, 5.251462e-17, 5.250679e-17, 5.256651e-17, 
    5.256617e-17, 5.25645e-17, 5.257186e-17, 5.257228e-17, 5.257885e-17, 
    5.257294e-17, 5.257048e-17, 5.256399e-17, 5.256027e-17, 5.25567e-17, 
    5.254884e-17, 5.254019e-17, 5.252792e-17, 5.251901e-17, 5.251308e-17, 
    5.251667e-17, 5.251351e-17, 5.251707e-17, 5.251871e-17, 5.250037e-17, 
    5.251071e-17, 5.249508e-17, 5.249592e-17, 5.250304e-17, 5.249583e-17, 
    5.256592e-17, 5.256791e-17, 5.257504e-17, 5.256946e-17, 5.257955e-17, 
    5.257398e-17, 5.257083e-17, 5.255832e-17, 5.255541e-17, 5.255293e-17, 
    5.254787e-17, 5.254147e-17, 5.253028e-17, 5.252046e-17, 5.251143e-17, 
    5.251208e-17, 5.251185e-17, 5.250991e-17, 5.251482e-17, 5.250909e-17, 
    5.250819e-17, 5.251064e-17, 5.249604e-17, 5.25002e-17, 5.249594e-17, 
    5.249863e-17, 5.256724e-17, 5.256386e-17, 5.25657e-17, 5.256228e-17, 
    5.256474e-17, 5.255399e-17, 5.255077e-17, 5.253555e-17, 5.254163e-17, 
    5.253178e-17, 5.254058e-17, 5.253905e-17, 5.253173e-17, 5.254006e-17, 
    5.252113e-17, 5.25342e-17, 5.250983e-17, 5.252311e-17, 5.250901e-17, 
    5.251147e-17, 5.250734e-17, 5.250371e-17, 5.249904e-17, 5.249061e-17, 
    5.249253e-17, 5.248539e-17, 5.255876e-17, 5.255443e-17, 5.25547e-17, 
    5.255009e-17, 5.254671e-17, 5.253924e-17, 5.252743e-17, 5.253183e-17, 
    5.252362e-17, 5.252201e-17, 5.253442e-17, 5.252692e-17, 5.255145e-17, 
    5.254761e-17, 5.25498e-17, 5.255848e-17, 5.253098e-17, 5.254516e-17, 
    5.251888e-17, 5.252652e-17, 5.250425e-17, 5.251543e-17, 5.249362e-17, 
    5.248464e-17, 5.247564e-17, 5.246579e-17, 5.255195e-17, 5.255489e-17, 
    5.25495e-17, 5.254228e-17, 5.253524e-17, 5.252608e-17, 5.252508e-17, 
    5.25234e-17, 5.25189e-17, 5.251519e-17, 5.252299e-17, 5.251425e-17, 
    5.254696e-17, 5.25297e-17, 5.255612e-17, 5.254832e-17, 5.254265e-17, 
    5.254502e-17, 5.25323e-17, 5.252935e-17, 5.251742e-17, 5.252352e-17, 
    5.248696e-17, 5.250312e-17, 5.245791e-17, 5.247058e-17, 5.255595e-17, 
    5.25519e-17, 5.253798e-17, 5.254458e-17, 5.252541e-17, 5.252074e-17, 
    5.251686e-17, 5.25121e-17, 5.251149e-17, 5.250865e-17, 5.251332e-17, 
    5.250879e-17, 5.252606e-17, 5.251832e-17, 5.253942e-17, 5.253435e-17, 
    5.253664e-17, 5.253924e-17, 5.253123e-17, 5.252289e-17, 5.252251e-17, 
    5.251988e-17, 5.251282e-17, 5.252532e-17, 5.248524e-17, 5.251029e-17, 
    5.254749e-17, 5.253996e-17, 5.253864e-17, 5.25416e-17, 5.252122e-17, 
    5.252863e-17, 5.25087e-17, 5.251403e-17, 5.250524e-17, 5.250962e-17, 
    5.251028e-17, 5.251587e-17, 5.25194e-17, 5.252832e-17, 5.253553e-17, 
    5.254115e-17, 5.253982e-17, 5.253365e-17, 5.252233e-17, 5.251153e-17, 
    5.251392e-17, 5.250591e-17, 5.25268e-17, 5.251813e-17, 5.252154e-17, 
    5.251261e-17, 5.253199e-17, 5.251608e-17, 5.253613e-17, 5.253433e-17, 
    5.252877e-17, 5.251767e-17, 5.251493e-17, 5.251236e-17, 5.251391e-17, 
    5.252201e-17, 5.252326e-17, 5.252886e-17, 5.25305e-17, 5.253471e-17, 
    5.253829e-17, 5.253507e-17, 5.253173e-17, 5.252193e-17, 5.251323e-17, 
    5.250369e-17, 5.250128e-17, 5.249065e-17, 5.249957e-17, 5.248513e-17, 
    5.249781e-17, 5.247569e-17, 5.251486e-17, 5.24978e-17, 5.252845e-17, 
    5.252509e-17, 5.251922e-17, 5.25054e-17, 5.251265e-17, 5.250407e-17, 
    5.25233e-17, 5.253353e-17, 5.253594e-17, 5.254084e-17, 5.253583e-17, 
    5.253623e-17, 5.253145e-17, 5.253297e-17, 5.25216e-17, 5.25277e-17, 
    5.251035e-17, 5.250409e-17, 5.24862e-17, 5.24754e-17, 5.246411e-17, 
    5.245923e-17, 5.245773e-17, 5.245712e-17 ;

 MEG_ethanol =
  4.221994e-18, 4.220502e-18, 4.220785e-18, 4.219598e-18, 4.220246e-18, 
    4.219477e-18, 4.221678e-18, 4.220454e-18, 4.221228e-18, 4.221842e-18, 
    4.217337e-18, 4.219542e-18, 4.214933e-18, 4.216355e-18, 4.212751e-18, 
    4.21517e-18, 4.212259e-18, 4.212792e-18, 4.211119e-18, 4.211596e-18, 
    4.209518e-18, 4.210898e-18, 4.208397e-18, 4.209832e-18, 4.209618e-18, 
    4.210948e-18, 4.219071e-18, 4.21762e-18, 4.219163e-18, 4.218954e-18, 
    4.219042e-18, 4.220242e-18, 4.220866e-18, 4.222088e-18, 4.221861e-18, 
    4.220953e-18, 4.21886e-18, 4.219551e-18, 4.217756e-18, 4.217795e-18, 
    4.215819e-18, 4.21671e-18, 4.213374e-18, 4.214314e-18, 4.211576e-18, 
    4.212268e-18, 4.211613e-18, 4.211808e-18, 4.21161e-18, 4.212624e-18, 
    4.212191e-18, 4.213075e-18, 4.216549e-18, 4.215536e-18, 4.218576e-18, 
    4.220451e-18, 4.22163e-18, 4.222488e-18, 4.222367e-18, 4.222141e-18, 
    4.220948e-18, 4.219804e-18, 4.218941e-18, 4.218369e-18, 4.217801e-18, 
    4.216159e-18, 4.215229e-18, 4.213197e-18, 4.21354e-18, 4.212941e-18, 
    4.212335e-18, 4.211352e-18, 4.21151e-18, 4.211083e-18, 4.21294e-18, 
    4.211714e-18, 4.213741e-18, 4.213189e-18, 4.217743e-18, 4.21936e-18, 
    4.220131e-18, 4.220734e-18, 4.222275e-18, 4.221216e-18, 4.221635e-18, 
    4.220617e-18, 4.219984e-18, 4.220293e-18, 4.218353e-18, 4.21911e-18, 
    4.215175e-18, 4.216867e-18, 4.212406e-18, 4.213467e-18, 4.212148e-18, 
    4.212816e-18, 4.21168e-18, 4.212702e-18, 4.210916e-18, 4.210538e-18, 
    4.210798e-18, 4.209768e-18, 4.212762e-18, 4.211622e-18, 4.220307e-18, 
    4.220256e-18, 4.220014e-18, 4.221085e-18, 4.221145e-18, 4.222099e-18, 
    4.221242e-18, 4.220884e-18, 4.21994e-18, 4.2194e-18, 4.21888e-18, 
    4.217738e-18, 4.216479e-18, 4.214695e-18, 4.2134e-18, 4.212537e-18, 
    4.21306e-18, 4.212599e-18, 4.213118e-18, 4.213357e-18, 4.210686e-18, 
    4.212193e-18, 4.209916e-18, 4.210038e-18, 4.211076e-18, 4.210025e-18, 
    4.22022e-18, 4.22051e-18, 4.221547e-18, 4.220735e-18, 4.222202e-18, 
    4.221393e-18, 4.220934e-18, 4.219116e-18, 4.218694e-18, 4.218332e-18, 
    4.217597e-18, 4.216665e-18, 4.215039e-18, 4.213612e-18, 4.212297e-18, 
    4.212391e-18, 4.212359e-18, 4.212075e-18, 4.212791e-18, 4.211957e-18, 
    4.211825e-18, 4.212182e-18, 4.210056e-18, 4.210661e-18, 4.210041e-18, 
    4.210433e-18, 4.220413e-18, 4.219921e-18, 4.220189e-18, 4.219691e-18, 
    4.220049e-18, 4.218486e-18, 4.218018e-18, 4.215805e-18, 4.216689e-18, 
    4.215256e-18, 4.216536e-18, 4.216315e-18, 4.21525e-18, 4.21646e-18, 
    4.213708e-18, 4.215609e-18, 4.212064e-18, 4.213996e-18, 4.211945e-18, 
    4.212302e-18, 4.211701e-18, 4.211174e-18, 4.210492e-18, 4.209265e-18, 
    4.209545e-18, 4.208504e-18, 4.219179e-18, 4.218551e-18, 4.218589e-18, 
    4.217919e-18, 4.217428e-18, 4.216342e-18, 4.214624e-18, 4.215264e-18, 
    4.21407e-18, 4.213836e-18, 4.21564e-18, 4.214549e-18, 4.218117e-18, 
    4.217559e-18, 4.217878e-18, 4.21914e-18, 4.215141e-18, 4.217202e-18, 
    4.213382e-18, 4.214493e-18, 4.211251e-18, 4.21288e-18, 4.209703e-18, 
    4.208395e-18, 4.207082e-18, 4.205647e-18, 4.218189e-18, 4.218617e-18, 
    4.217834e-18, 4.216784e-18, 4.21576e-18, 4.214428e-18, 4.214282e-18, 
    4.214038e-18, 4.213384e-18, 4.212844e-18, 4.213978e-18, 4.212707e-18, 
    4.217465e-18, 4.214954e-18, 4.218796e-18, 4.217662e-18, 4.216838e-18, 
    4.217181e-18, 4.215333e-18, 4.214904e-18, 4.213169e-18, 4.214055e-18, 
    4.208733e-18, 4.211087e-18, 4.204497e-18, 4.206345e-18, 4.218772e-18, 
    4.218182e-18, 4.216158e-18, 4.217117e-18, 4.21433e-18, 4.213653e-18, 
    4.213087e-18, 4.212394e-18, 4.212306e-18, 4.211893e-18, 4.212572e-18, 
    4.211913e-18, 4.214425e-18, 4.213299e-18, 4.216367e-18, 4.21563e-18, 
    4.215963e-18, 4.216342e-18, 4.215176e-18, 4.213965e-18, 4.21391e-18, 
    4.213527e-18, 4.212499e-18, 4.214318e-18, 4.208482e-18, 4.212131e-18, 
    4.217541e-18, 4.216446e-18, 4.216255e-18, 4.216685e-18, 4.213721e-18, 
    4.214798e-18, 4.211899e-18, 4.212675e-18, 4.211396e-18, 4.212034e-18, 
    4.212129e-18, 4.212943e-18, 4.213457e-18, 4.214754e-18, 4.215802e-18, 
    4.216619e-18, 4.216426e-18, 4.215529e-18, 4.213883e-18, 4.212311e-18, 
    4.212659e-18, 4.211493e-18, 4.214532e-18, 4.213271e-18, 4.213768e-18, 
    4.212469e-18, 4.215287e-18, 4.212974e-18, 4.21589e-18, 4.215628e-18, 
    4.214819e-18, 4.213206e-18, 4.212806e-18, 4.212432e-18, 4.212657e-18, 
    4.213837e-18, 4.214018e-18, 4.214832e-18, 4.215071e-18, 4.215683e-18, 
    4.216203e-18, 4.215735e-18, 4.215249e-18, 4.213825e-18, 4.212558e-18, 
    4.21117e-18, 4.21082e-18, 4.209272e-18, 4.210571e-18, 4.208467e-18, 
    4.210314e-18, 4.20709e-18, 4.212797e-18, 4.210312e-18, 4.214773e-18, 
    4.214284e-18, 4.213431e-18, 4.211418e-18, 4.212474e-18, 4.211225e-18, 
    4.214023e-18, 4.215512e-18, 4.215862e-18, 4.216574e-18, 4.215846e-18, 
    4.215903e-18, 4.215209e-18, 4.21543e-18, 4.213777e-18, 4.214663e-18, 
    4.212139e-18, 4.211228e-18, 4.208623e-18, 4.207048e-18, 4.205401e-18, 
    4.20469e-18, 4.204471e-18, 4.204381e-18 ;

 MEG_formaldehyde =
  8.443987e-19, 8.441003e-19, 8.441569e-19, 8.439196e-19, 8.440491e-19, 
    8.438954e-19, 8.443356e-19, 8.440907e-19, 8.442456e-19, 8.443684e-19, 
    8.434673e-19, 8.439083e-19, 8.429866e-19, 8.432709e-19, 8.425502e-19, 
    8.43034e-19, 8.424517e-19, 8.425584e-19, 8.422237e-19, 8.423192e-19, 
    8.419035e-19, 8.421796e-19, 8.416793e-19, 8.419663e-19, 8.419236e-19, 
    8.421896e-19, 8.438141e-19, 8.435239e-19, 8.438326e-19, 8.437909e-19, 
    8.438084e-19, 8.440484e-19, 8.441732e-19, 8.444177e-19, 8.443722e-19, 
    8.441906e-19, 8.43772e-19, 8.439102e-19, 8.435511e-19, 8.43559e-19, 
    8.431638e-19, 8.43342e-19, 8.426747e-19, 8.428629e-19, 8.423151e-19, 
    8.424535e-19, 8.423226e-19, 8.423615e-19, 8.423221e-19, 8.425248e-19, 
    8.424382e-19, 8.426149e-19, 8.433097e-19, 8.431071e-19, 8.437152e-19, 
    8.440903e-19, 8.443259e-19, 8.444976e-19, 8.444733e-19, 8.444282e-19, 
    8.441896e-19, 8.439608e-19, 8.437882e-19, 8.436738e-19, 8.435602e-19, 
    8.432318e-19, 8.430458e-19, 8.426395e-19, 8.427079e-19, 8.425882e-19, 
    8.424671e-19, 8.422704e-19, 8.42302e-19, 8.422165e-19, 8.425878e-19, 
    8.423427e-19, 8.427481e-19, 8.426378e-19, 8.435486e-19, 8.43872e-19, 
    8.440262e-19, 8.441468e-19, 8.44455e-19, 8.442432e-19, 8.443271e-19, 
    8.441234e-19, 8.439968e-19, 8.440586e-19, 8.436706e-19, 8.438221e-19, 
    8.430349e-19, 8.433734e-19, 8.424812e-19, 8.426935e-19, 8.424297e-19, 
    8.425633e-19, 8.423359e-19, 8.425405e-19, 8.421832e-19, 8.421076e-19, 
    8.421596e-19, 8.419535e-19, 8.425523e-19, 8.423244e-19, 8.440612e-19, 
    8.440513e-19, 8.440027e-19, 8.442169e-19, 8.44229e-19, 8.444198e-19, 
    8.442482e-19, 8.441768e-19, 8.43988e-19, 8.438799e-19, 8.43776e-19, 
    8.435476e-19, 8.432958e-19, 8.42939e-19, 8.426799e-19, 8.425074e-19, 
    8.426119e-19, 8.425198e-19, 8.426235e-19, 8.426713e-19, 8.421372e-19, 
    8.424385e-19, 8.419832e-19, 8.420077e-19, 8.422152e-19, 8.420049e-19, 
    8.44044e-19, 8.441019e-19, 8.443095e-19, 8.44147e-19, 8.444404e-19, 
    8.442785e-19, 8.441869e-19, 8.438231e-19, 8.437386e-19, 8.436664e-19, 
    8.435193e-19, 8.43333e-19, 8.430078e-19, 8.427223e-19, 8.424593e-19, 
    8.424782e-19, 8.424717e-19, 8.424149e-19, 8.425581e-19, 8.423913e-19, 
    8.423651e-19, 8.424364e-19, 8.420111e-19, 8.421322e-19, 8.420082e-19, 
    8.420866e-19, 8.440826e-19, 8.439842e-19, 8.440377e-19, 8.439383e-19, 
    8.440098e-19, 8.436972e-19, 8.436036e-19, 8.43161e-19, 8.433377e-19, 
    8.430512e-19, 8.433071e-19, 8.432628e-19, 8.430499e-19, 8.43292e-19, 
    8.427416e-19, 8.431217e-19, 8.424127e-19, 8.427992e-19, 8.423889e-19, 
    8.424604e-19, 8.423402e-19, 8.422346e-19, 8.420985e-19, 8.418529e-19, 
    8.419089e-19, 8.417007e-19, 8.438359e-19, 8.437102e-19, 8.437177e-19, 
    8.435838e-19, 8.434856e-19, 8.432684e-19, 8.429248e-19, 8.430528e-19, 
    8.42814e-19, 8.427672e-19, 8.43128e-19, 8.429099e-19, 8.436234e-19, 
    8.435117e-19, 8.435755e-19, 8.43828e-19, 8.430282e-19, 8.434404e-19, 
    8.426763e-19, 8.428984e-19, 8.422502e-19, 8.425759e-19, 8.419406e-19, 
    8.416789e-19, 8.414164e-19, 8.411293e-19, 8.436378e-19, 8.437235e-19, 
    8.435668e-19, 8.433568e-19, 8.431519e-19, 8.428856e-19, 8.428564e-19, 
    8.428076e-19, 8.426768e-19, 8.425687e-19, 8.427956e-19, 8.425413e-19, 
    8.434929e-19, 8.429908e-19, 8.437592e-19, 8.435324e-19, 8.433676e-19, 
    8.434362e-19, 8.430665e-19, 8.429807e-19, 8.426338e-19, 8.42811e-19, 
    8.417466e-19, 8.422173e-19, 8.408993e-19, 8.41269e-19, 8.437544e-19, 
    8.436363e-19, 8.432315e-19, 8.434234e-19, 8.428659e-19, 8.427305e-19, 
    8.426174e-19, 8.424787e-19, 8.424611e-19, 8.423786e-19, 8.425143e-19, 
    8.423826e-19, 8.428851e-19, 8.426597e-19, 8.432735e-19, 8.431261e-19, 
    8.431926e-19, 8.432683e-19, 8.430352e-19, 8.427929e-19, 8.42782e-19, 
    8.427054e-19, 8.424998e-19, 8.428635e-19, 8.416964e-19, 8.424262e-19, 
    8.435081e-19, 8.432892e-19, 8.432509e-19, 8.433369e-19, 8.427442e-19, 
    8.429595e-19, 8.423798e-19, 8.42535e-19, 8.422792e-19, 8.424068e-19, 
    8.424259e-19, 8.425885e-19, 8.426915e-19, 8.429508e-19, 8.431603e-19, 
    8.433237e-19, 8.432853e-19, 8.431057e-19, 8.427767e-19, 8.424622e-19, 
    8.425317e-19, 8.422986e-19, 8.429065e-19, 8.426543e-19, 8.427535e-19, 
    8.424937e-19, 8.430574e-19, 8.425947e-19, 8.431779e-19, 8.431255e-19, 
    8.429637e-19, 8.426411e-19, 8.425612e-19, 8.424863e-19, 8.425314e-19, 
    8.427673e-19, 8.428036e-19, 8.429663e-19, 8.430141e-19, 8.431365e-19, 
    8.432406e-19, 8.431469e-19, 8.430498e-19, 8.427649e-19, 8.425117e-19, 
    8.422341e-19, 8.421639e-19, 8.418543e-19, 8.421141e-19, 8.416935e-19, 
    8.420628e-19, 8.414179e-19, 8.425593e-19, 8.420623e-19, 8.429545e-19, 
    8.428568e-19, 8.426862e-19, 8.422836e-19, 8.424948e-19, 8.422451e-19, 
    8.428045e-19, 8.431023e-19, 8.431723e-19, 8.433148e-19, 8.431691e-19, 
    8.431807e-19, 8.430417e-19, 8.43086e-19, 8.427553e-19, 8.429327e-19, 
    8.424278e-19, 8.422455e-19, 8.417246e-19, 8.414095e-19, 8.410801e-19, 
    8.409379e-19, 8.408942e-19, 8.408762e-19 ;

 MEG_isoprene =
  6.667447e-19, 6.664678e-19, 6.665204e-19, 6.663001e-19, 6.664203e-19, 
    6.662776e-19, 6.666862e-19, 6.66459e-19, 6.666027e-19, 6.667167e-19, 
    6.658802e-19, 6.662896e-19, 6.65434e-19, 6.656979e-19, 6.650289e-19, 
    6.65478e-19, 6.649375e-19, 6.650365e-19, 6.647258e-19, 6.648144e-19, 
    6.644284e-19, 6.646848e-19, 6.642202e-19, 6.644867e-19, 6.64447e-19, 
    6.646941e-19, 6.662022e-19, 6.659328e-19, 6.662194e-19, 6.661806e-19, 
    6.661969e-19, 6.664197e-19, 6.665355e-19, 6.667624e-19, 6.667202e-19, 
    6.665516e-19, 6.661631e-19, 6.662914e-19, 6.65958e-19, 6.659654e-19, 
    6.655985e-19, 6.657639e-19, 6.651445e-19, 6.653192e-19, 6.648106e-19, 
    6.649391e-19, 6.648175e-19, 6.648537e-19, 6.648171e-19, 6.650053e-19, 
    6.649249e-19, 6.650889e-19, 6.657339e-19, 6.655459e-19, 6.661103e-19, 
    6.664585e-19, 6.666772e-19, 6.668366e-19, 6.668141e-19, 6.667722e-19, 
    6.665507e-19, 6.663383e-19, 6.661781e-19, 6.660719e-19, 6.659665e-19, 
    6.656617e-19, 6.65489e-19, 6.651117e-19, 6.651753e-19, 6.650642e-19, 
    6.649517e-19, 6.647691e-19, 6.647984e-19, 6.647191e-19, 6.650639e-19, 
    6.648362e-19, 6.652126e-19, 6.651102e-19, 6.659557e-19, 6.662559e-19, 
    6.663991e-19, 6.665109e-19, 6.667971e-19, 6.666005e-19, 6.666783e-19, 
    6.664893e-19, 6.663718e-19, 6.664291e-19, 6.66069e-19, 6.662096e-19, 
    6.654788e-19, 6.65793e-19, 6.649648e-19, 6.651619e-19, 6.64917e-19, 
    6.65041e-19, 6.648299e-19, 6.650198e-19, 6.646881e-19, 6.64618e-19, 
    6.646662e-19, 6.644749e-19, 6.650308e-19, 6.648192e-19, 6.664316e-19, 
    6.664224e-19, 6.663772e-19, 6.665761e-19, 6.665873e-19, 6.667644e-19, 
    6.666052e-19, 6.665388e-19, 6.663636e-19, 6.662633e-19, 6.661668e-19, 
    6.659547e-19, 6.657211e-19, 6.653898e-19, 6.651493e-19, 6.649892e-19, 
    6.650862e-19, 6.650007e-19, 6.650969e-19, 6.651413e-19, 6.646454e-19, 
    6.649252e-19, 6.645024e-19, 6.645251e-19, 6.647178e-19, 6.645226e-19, 
    6.664156e-19, 6.664693e-19, 6.666619e-19, 6.665112e-19, 6.667835e-19, 
    6.666333e-19, 6.665482e-19, 6.662105e-19, 6.661321e-19, 6.660651e-19, 
    6.659285e-19, 6.657556e-19, 6.654537e-19, 6.651886e-19, 6.649444e-19, 
    6.64962e-19, 6.64956e-19, 6.649033e-19, 6.650362e-19, 6.648813e-19, 
    6.64857e-19, 6.649231e-19, 6.645283e-19, 6.646408e-19, 6.645256e-19, 
    6.645984e-19, 6.664514e-19, 6.663601e-19, 6.664097e-19, 6.663174e-19, 
    6.663838e-19, 6.660937e-19, 6.660067e-19, 6.655959e-19, 6.657599e-19, 
    6.65494e-19, 6.657315e-19, 6.656904e-19, 6.654928e-19, 6.657175e-19, 
    6.652066e-19, 6.655594e-19, 6.649012e-19, 6.652601e-19, 6.648791e-19, 
    6.649455e-19, 6.648339e-19, 6.647359e-19, 6.646094e-19, 6.643814e-19, 
    6.644334e-19, 6.642401e-19, 6.662224e-19, 6.661057e-19, 6.661127e-19, 
    6.659883e-19, 6.658972e-19, 6.656956e-19, 6.653766e-19, 6.654954e-19, 
    6.652737e-19, 6.652303e-19, 6.655653e-19, 6.653627e-19, 6.660251e-19, 
    6.659214e-19, 6.659807e-19, 6.662151e-19, 6.654726e-19, 6.658553e-19, 
    6.65146e-19, 6.653522e-19, 6.647503e-19, 6.650527e-19, 6.644629e-19, 
    6.642199e-19, 6.639761e-19, 6.637094e-19, 6.660385e-19, 6.661181e-19, 
    6.659726e-19, 6.657777e-19, 6.655875e-19, 6.653402e-19, 6.653131e-19, 
    6.652679e-19, 6.651464e-19, 6.650461e-19, 6.652567e-19, 6.650206e-19, 
    6.65904e-19, 6.65438e-19, 6.661512e-19, 6.659407e-19, 6.657876e-19, 
    6.658514e-19, 6.655082e-19, 6.654285e-19, 6.651065e-19, 6.65271e-19, 
    6.642827e-19, 6.647198e-19, 6.634957e-19, 6.638392e-19, 6.661467e-19, 
    6.660371e-19, 6.656613e-19, 6.658396e-19, 6.65322e-19, 6.651962e-19, 
    6.650912e-19, 6.649625e-19, 6.649461e-19, 6.648695e-19, 6.649955e-19, 
    6.648732e-19, 6.653397e-19, 6.651306e-19, 6.657003e-19, 6.655634e-19, 
    6.656253e-19, 6.656955e-19, 6.654791e-19, 6.652542e-19, 6.65244e-19, 
    6.651729e-19, 6.649821e-19, 6.653197e-19, 6.642362e-19, 6.649138e-19, 
    6.659181e-19, 6.657149e-19, 6.656793e-19, 6.657592e-19, 6.65209e-19, 
    6.654089e-19, 6.648707e-19, 6.650148e-19, 6.647773e-19, 6.648957e-19, 
    6.649134e-19, 6.650644e-19, 6.6516e-19, 6.654007e-19, 6.655953e-19, 
    6.657469e-19, 6.657112e-19, 6.655446e-19, 6.652392e-19, 6.649471e-19, 
    6.650118e-19, 6.647952e-19, 6.653596e-19, 6.651255e-19, 6.652176e-19, 
    6.649764e-19, 6.654997e-19, 6.650702e-19, 6.656116e-19, 6.65563e-19, 
    6.654128e-19, 6.651132e-19, 6.65039e-19, 6.649696e-19, 6.650114e-19, 
    6.652304e-19, 6.652641e-19, 6.654152e-19, 6.654596e-19, 6.655731e-19, 
    6.656698e-19, 6.655828e-19, 6.654927e-19, 6.652282e-19, 6.649931e-19, 
    6.647353e-19, 6.646702e-19, 6.643827e-19, 6.64624e-19, 6.642334e-19, 
    6.645763e-19, 6.639775e-19, 6.650373e-19, 6.645759e-19, 6.654041e-19, 
    6.653135e-19, 6.651552e-19, 6.647814e-19, 6.649775e-19, 6.647456e-19, 
    6.65265e-19, 6.655415e-19, 6.656064e-19, 6.657387e-19, 6.656034e-19, 
    6.656141e-19, 6.654852e-19, 6.655263e-19, 6.652193e-19, 6.653839e-19, 
    6.649153e-19, 6.64746e-19, 6.642623e-19, 6.639697e-19, 6.636638e-19, 
    6.635317e-19, 6.63491e-19, 6.634743e-19 ;

 MEG_methanol =
  9.493388e-17, 9.491827e-17, 9.492123e-17, 9.490882e-17, 9.491559e-17, 
    9.490755e-17, 9.493059e-17, 9.491776e-17, 9.492587e-17, 9.49323e-17, 
    9.488515e-17, 9.490822e-17, 9.486e-17, 9.487488e-17, 9.483717e-17, 
    9.486248e-17, 9.483202e-17, 9.48376e-17, 9.482012e-17, 9.482511e-17, 
    9.480338e-17, 9.481781e-17, 9.479169e-17, 9.480667e-17, 9.480443e-17, 
    9.481833e-17, 9.490329e-17, 9.48881e-17, 9.490426e-17, 9.490208e-17, 
    9.4903e-17, 9.491555e-17, 9.492209e-17, 9.493488e-17, 9.49325e-17, 
    9.492299e-17, 9.490109e-17, 9.490833e-17, 9.488954e-17, 9.488996e-17, 
    9.486927e-17, 9.48786e-17, 9.484368e-17, 9.485354e-17, 9.482489e-17, 
    9.483212e-17, 9.482528e-17, 9.482732e-17, 9.482525e-17, 9.483585e-17, 
    9.483132e-17, 9.484056e-17, 9.487691e-17, 9.486631e-17, 9.489812e-17, 
    9.491774e-17, 9.493008e-17, 9.493907e-17, 9.49378e-17, 9.493543e-17, 
    9.492294e-17, 9.491097e-17, 9.490194e-17, 9.489596e-17, 9.489002e-17, 
    9.487283e-17, 9.48631e-17, 9.484184e-17, 9.484542e-17, 9.483916e-17, 
    9.483283e-17, 9.482255e-17, 9.482421e-17, 9.481974e-17, 9.483914e-17, 
    9.482633e-17, 9.484752e-17, 9.484175e-17, 9.48894e-17, 9.490633e-17, 
    9.491439e-17, 9.49207e-17, 9.493684e-17, 9.492574e-17, 9.493014e-17, 
    9.491948e-17, 9.491285e-17, 9.491609e-17, 9.489579e-17, 9.490372e-17, 
    9.486253e-17, 9.488024e-17, 9.483357e-17, 9.484467e-17, 9.483088e-17, 
    9.483786e-17, 9.482597e-17, 9.483667e-17, 9.4818e-17, 9.481405e-17, 
    9.481677e-17, 9.4806e-17, 9.483728e-17, 9.482537e-17, 9.491623e-17, 
    9.491571e-17, 9.491317e-17, 9.492438e-17, 9.4925e-17, 9.4935e-17, 
    9.492602e-17, 9.492228e-17, 9.491239e-17, 9.490674e-17, 9.49013e-17, 
    9.488936e-17, 9.487618e-17, 9.485751e-17, 9.484396e-17, 9.483494e-17, 
    9.48404e-17, 9.483559e-17, 9.484101e-17, 9.484351e-17, 9.481559e-17, 
    9.483133e-17, 9.480755e-17, 9.480883e-17, 9.481967e-17, 9.480869e-17, 
    9.491532e-17, 9.491836e-17, 9.492922e-17, 9.492072e-17, 9.493607e-17, 
    9.49276e-17, 9.49228e-17, 9.490377e-17, 9.489935e-17, 9.489557e-17, 
    9.488788e-17, 9.487813e-17, 9.486111e-17, 9.484617e-17, 9.483242e-17, 
    9.483341e-17, 9.483307e-17, 9.48301e-17, 9.483759e-17, 9.482887e-17, 
    9.48275e-17, 9.483122e-17, 9.480901e-17, 9.481533e-17, 9.480886e-17, 
    9.481295e-17, 9.491735e-17, 9.49122e-17, 9.491499e-17, 9.490979e-17, 
    9.491353e-17, 9.489718e-17, 9.489228e-17, 9.486913e-17, 9.487838e-17, 
    9.486338e-17, 9.487678e-17, 9.487445e-17, 9.486331e-17, 9.487599e-17, 
    9.484718e-17, 9.486707e-17, 9.482999e-17, 9.485019e-17, 9.482875e-17, 
    9.483249e-17, 9.48262e-17, 9.482069e-17, 9.481357e-17, 9.480075e-17, 
    9.480367e-17, 9.479281e-17, 9.490444e-17, 9.489786e-17, 9.489826e-17, 
    9.489125e-17, 9.488611e-17, 9.487475e-17, 9.485677e-17, 9.486347e-17, 
    9.485097e-17, 9.484852e-17, 9.486741e-17, 9.485599e-17, 9.489332e-17, 
    9.488748e-17, 9.489082e-17, 9.490402e-17, 9.486218e-17, 9.488374e-17, 
    9.484377e-17, 9.485539e-17, 9.48215e-17, 9.483851e-17, 9.480533e-17, 
    9.479166e-17, 9.477798e-17, 9.4763e-17, 9.489407e-17, 9.489855e-17, 
    9.489036e-17, 9.487937e-17, 9.486866e-17, 9.485473e-17, 9.48532e-17, 
    9.485064e-17, 9.484379e-17, 9.483814e-17, 9.485001e-17, 9.483671e-17, 
    9.488648e-17, 9.486023e-17, 9.490042e-17, 9.488856e-17, 9.487994e-17, 
    9.488353e-17, 9.486418e-17, 9.48597e-17, 9.484154e-17, 9.485082e-17, 
    9.47952e-17, 9.481977e-17, 9.475101e-17, 9.477028e-17, 9.490017e-17, 
    9.4894e-17, 9.487282e-17, 9.488286e-17, 9.485369e-17, 9.48466e-17, 
    9.484068e-17, 9.483344e-17, 9.483252e-17, 9.48282e-17, 9.48353e-17, 
    9.482842e-17, 9.485469e-17, 9.48429e-17, 9.487502e-17, 9.48673e-17, 
    9.487079e-17, 9.487474e-17, 9.486255e-17, 9.484986e-17, 9.484929e-17, 
    9.484528e-17, 9.483453e-17, 9.485357e-17, 9.479257e-17, 9.483068e-17, 
    9.48873e-17, 9.487583e-17, 9.487383e-17, 9.487834e-17, 9.484732e-17, 
    9.485859e-17, 9.482827e-17, 9.483638e-17, 9.482302e-17, 9.482968e-17, 
    9.483068e-17, 9.483918e-17, 9.484456e-17, 9.485813e-17, 9.486909e-17, 
    9.487764e-17, 9.487563e-17, 9.486623e-17, 9.484902e-17, 9.483257e-17, 
    9.483621e-17, 9.482403e-17, 9.485581e-17, 9.484262e-17, 9.48478e-17, 
    9.483423e-17, 9.486371e-17, 9.483949e-17, 9.487001e-17, 9.486727e-17, 
    9.485881e-17, 9.484192e-17, 9.483775e-17, 9.483384e-17, 9.483619e-17, 
    9.484852e-17, 9.485043e-17, 9.485894e-17, 9.486144e-17, 9.486785e-17, 
    9.48733e-17, 9.486839e-17, 9.486331e-17, 9.48484e-17, 9.483516e-17, 
    9.482065e-17, 9.481699e-17, 9.480081e-17, 9.481438e-17, 9.479242e-17, 
    9.481169e-17, 9.477804e-17, 9.483765e-17, 9.481167e-17, 9.485833e-17, 
    9.485322e-17, 9.484428e-17, 9.482324e-17, 9.483428e-17, 9.482123e-17, 
    9.485048e-17, 9.486606e-17, 9.486972e-17, 9.487718e-17, 9.486956e-17, 
    9.487016e-17, 9.486289e-17, 9.486521e-17, 9.48479e-17, 9.485718e-17, 
    9.483078e-17, 9.482126e-17, 9.479405e-17, 9.477761e-17, 9.476044e-17, 
    9.475303e-17, 9.475075e-17, 9.474981e-17 ;

 MEG_pinene_a =
  8.100023e-17, 8.098319e-17, 8.098641e-17, 8.097287e-17, 8.098026e-17, 
    8.097148e-17, 8.099663e-17, 8.098264e-17, 8.099148e-17, 8.09985e-17, 
    8.094703e-17, 8.097222e-17, 8.091959e-17, 8.093582e-17, 8.089468e-17, 
    8.09223e-17, 8.088906e-17, 8.089515e-17, 8.087606e-17, 8.08815e-17, 
    8.085779e-17, 8.087354e-17, 8.084502e-17, 8.086138e-17, 8.085894e-17, 
    8.087411e-17, 8.096684e-17, 8.095027e-17, 8.09679e-17, 8.096552e-17, 
    8.096652e-17, 8.098022e-17, 8.098735e-17, 8.100132e-17, 8.099872e-17, 
    8.098834e-17, 8.096444e-17, 8.097233e-17, 8.095183e-17, 8.095228e-17, 
    8.092971e-17, 8.093989e-17, 8.090178e-17, 8.091253e-17, 8.088127e-17, 
    8.088916e-17, 8.088169e-17, 8.088392e-17, 8.088167e-17, 8.089323e-17, 
    8.088829e-17, 8.089837e-17, 8.093804e-17, 8.092647e-17, 8.09612e-17, 
    8.098261e-17, 8.099607e-17, 8.100588e-17, 8.100449e-17, 8.100192e-17, 
    8.098829e-17, 8.097522e-17, 8.096536e-17, 8.095883e-17, 8.095235e-17, 
    8.093359e-17, 8.092297e-17, 8.089977e-17, 8.090368e-17, 8.089685e-17, 
    8.088994e-17, 8.087872e-17, 8.088052e-17, 8.087565e-17, 8.089683e-17, 
    8.088284e-17, 8.090597e-17, 8.089968e-17, 8.095167e-17, 8.097015e-17, 
    8.097895e-17, 8.098584e-17, 8.100345e-17, 8.099134e-17, 8.099614e-17, 
    8.098451e-17, 8.097728e-17, 8.09808e-17, 8.095865e-17, 8.09673e-17, 
    8.092235e-17, 8.094167e-17, 8.089075e-17, 8.090286e-17, 8.08878e-17, 
    8.089543e-17, 8.088245e-17, 8.089412e-17, 8.087375e-17, 8.086943e-17, 
    8.08724e-17, 8.086065e-17, 8.08948e-17, 8.08818e-17, 8.098096e-17, 
    8.098039e-17, 8.097761e-17, 8.098985e-17, 8.099054e-17, 8.100144e-17, 
    8.099164e-17, 8.098755e-17, 8.097677e-17, 8.09706e-17, 8.096466e-17, 
    8.095162e-17, 8.093725e-17, 8.091688e-17, 8.090208e-17, 8.089224e-17, 
    8.08982e-17, 8.089295e-17, 8.089887e-17, 8.090159e-17, 8.087112e-17, 
    8.08883e-17, 8.086234e-17, 8.086373e-17, 8.087557e-17, 8.086358e-17, 
    8.097997e-17, 8.098328e-17, 8.099513e-17, 8.098585e-17, 8.100261e-17, 
    8.099336e-17, 8.098813e-17, 8.096736e-17, 8.096253e-17, 8.095841e-17, 
    8.095001e-17, 8.093938e-17, 8.09208e-17, 8.09045e-17, 8.088949e-17, 
    8.089057e-17, 8.08902e-17, 8.088696e-17, 8.089513e-17, 8.088561e-17, 
    8.088412e-17, 8.088819e-17, 8.086393e-17, 8.087083e-17, 8.086377e-17, 
    8.086823e-17, 8.098217e-17, 8.097655e-17, 8.097961e-17, 8.097393e-17, 
    8.097802e-17, 8.096016e-17, 8.095482e-17, 8.092954e-17, 8.093964e-17, 
    8.092328e-17, 8.09379e-17, 8.093537e-17, 8.092321e-17, 8.093704e-17, 
    8.09056e-17, 8.092731e-17, 8.088684e-17, 8.090889e-17, 8.088548e-17, 
    8.088956e-17, 8.08827e-17, 8.087668e-17, 8.086891e-17, 8.085491e-17, 
    8.085811e-17, 8.084624e-17, 8.096808e-17, 8.096091e-17, 8.096134e-17, 
    8.095369e-17, 8.094809e-17, 8.093569e-17, 8.091606e-17, 8.092337e-17, 
    8.090974e-17, 8.090707e-17, 8.092767e-17, 8.091521e-17, 8.095595e-17, 
    8.094958e-17, 8.095322e-17, 8.096763e-17, 8.092197e-17, 8.094551e-17, 
    8.090188e-17, 8.091456e-17, 8.087756e-17, 8.089615e-17, 8.085992e-17, 
    8.084499e-17, 8.083004e-17, 8.081368e-17, 8.095678e-17, 8.096167e-17, 
    8.095272e-17, 8.094073e-17, 8.092904e-17, 8.091383e-17, 8.091216e-17, 
    8.090938e-17, 8.09019e-17, 8.089574e-17, 8.090869e-17, 8.089417e-17, 
    8.09485e-17, 8.091984e-17, 8.09637e-17, 8.095076e-17, 8.094134e-17, 
    8.094527e-17, 8.092416e-17, 8.091926e-17, 8.089945e-17, 8.090957e-17, 
    8.084885e-17, 8.087569e-17, 8.080058e-17, 8.082164e-17, 8.096343e-17, 
    8.09567e-17, 8.093357e-17, 8.094454e-17, 8.091271e-17, 8.090497e-17, 
    8.089852e-17, 8.08906e-17, 8.08896e-17, 8.088489e-17, 8.089263e-17, 
    8.088512e-17, 8.09138e-17, 8.090093e-17, 8.093598e-17, 8.092755e-17, 
    8.093136e-17, 8.093568e-17, 8.092236e-17, 8.090853e-17, 8.090791e-17, 
    8.090353e-17, 8.08918e-17, 8.091256e-17, 8.084599e-17, 8.08876e-17, 
    8.094938e-17, 8.093687e-17, 8.093469e-17, 8.09396e-17, 8.090575e-17, 
    8.091805e-17, 8.088496e-17, 8.089382e-17, 8.087922e-17, 8.08865e-17, 
    8.088758e-17, 8.089687e-17, 8.090274e-17, 8.091755e-17, 8.092951e-17, 
    8.093884e-17, 8.093665e-17, 8.092639e-17, 8.09076e-17, 8.088965e-17, 
    8.089363e-17, 8.088032e-17, 8.091502e-17, 8.090062e-17, 8.090628e-17, 
    8.089145e-17, 8.092364e-17, 8.089721e-17, 8.093052e-17, 8.092753e-17, 
    8.091829e-17, 8.089987e-17, 8.089531e-17, 8.089104e-17, 8.089361e-17, 
    8.090707e-17, 8.090914e-17, 8.091843e-17, 8.092117e-17, 8.092815e-17, 
    8.09341e-17, 8.092875e-17, 8.09232e-17, 8.090693e-17, 8.089248e-17, 
    8.087664e-17, 8.087264e-17, 8.085499e-17, 8.08698e-17, 8.084582e-17, 
    8.086686e-17, 8.083012e-17, 8.089519e-17, 8.086684e-17, 8.091776e-17, 
    8.091219e-17, 8.090244e-17, 8.087947e-17, 8.089152e-17, 8.087727e-17, 
    8.09092e-17, 8.09262e-17, 8.09302e-17, 8.093833e-17, 8.093001e-17, 
    8.093068e-17, 8.092274e-17, 8.092527e-17, 8.090638e-17, 8.091651e-17, 
    8.08877e-17, 8.08773e-17, 8.084759e-17, 8.082964e-17, 8.081089e-17, 
    8.080279e-17, 8.08003e-17, 8.079927e-17 ;

 MEG_thujene_a =
  1.951962e-18, 1.951581e-18, 1.951654e-18, 1.951351e-18, 1.951516e-18, 
    1.95132e-18, 1.951882e-18, 1.951569e-18, 1.951767e-18, 1.951924e-18, 
    1.950773e-18, 1.951336e-18, 1.95016e-18, 1.950523e-18, 1.949603e-18, 
    1.95022e-18, 1.949477e-18, 1.949613e-18, 1.949186e-18, 1.949308e-18, 
    1.948778e-18, 1.94913e-18, 1.948493e-18, 1.948858e-18, 1.948804e-18, 
    1.949143e-18, 1.951216e-18, 1.950846e-18, 1.95124e-18, 1.951186e-18, 
    1.951209e-18, 1.951515e-18, 1.951675e-18, 1.951987e-18, 1.951929e-18, 
    1.951697e-18, 1.951162e-18, 1.951339e-18, 1.95088e-18, 1.95089e-18, 
    1.950386e-18, 1.950613e-18, 1.949761e-18, 1.950002e-18, 1.949303e-18, 
    1.949479e-18, 1.949313e-18, 1.949362e-18, 1.949312e-18, 1.94957e-18, 
    1.94946e-18, 1.949685e-18, 1.950572e-18, 1.950313e-18, 1.95109e-18, 
    1.951568e-18, 1.95187e-18, 1.952089e-18, 1.952058e-18, 1.952e-18, 
    1.951695e-18, 1.951403e-18, 1.951183e-18, 1.951037e-18, 1.950892e-18, 
    1.950473e-18, 1.950235e-18, 1.949717e-18, 1.949804e-18, 1.949651e-18, 
    1.949497e-18, 1.949246e-18, 1.949286e-18, 1.949177e-18, 1.949651e-18, 
    1.949338e-18, 1.949855e-18, 1.949714e-18, 1.950877e-18, 1.95129e-18, 
    1.951487e-18, 1.951641e-18, 1.952035e-18, 1.951764e-18, 1.951871e-18, 
    1.951611e-18, 1.951449e-18, 1.951528e-18, 1.951033e-18, 1.951226e-18, 
    1.950221e-18, 1.950653e-18, 1.949515e-18, 1.949785e-18, 1.949449e-18, 
    1.949619e-18, 1.949329e-18, 1.94959e-18, 1.949135e-18, 1.949038e-18, 
    1.949105e-18, 1.948842e-18, 1.949605e-18, 1.949315e-18, 1.951532e-18, 
    1.951519e-18, 1.951457e-18, 1.95173e-18, 1.951746e-18, 1.951989e-18, 
    1.95177e-18, 1.951679e-18, 1.951438e-18, 1.9513e-18, 1.951167e-18, 
    1.950876e-18, 1.950554e-18, 1.950099e-18, 1.949768e-18, 1.949548e-18, 
    1.949681e-18, 1.949564e-18, 1.949696e-18, 1.949757e-18, 1.949076e-18, 
    1.94946e-18, 1.94888e-18, 1.948911e-18, 1.949175e-18, 1.948908e-18, 
    1.95151e-18, 1.951584e-18, 1.951848e-18, 1.951641e-18, 1.952016e-18, 
    1.951809e-18, 1.951692e-18, 1.951227e-18, 1.95112e-18, 1.951027e-18, 
    1.95084e-18, 1.950602e-18, 1.950187e-18, 1.949822e-18, 1.949487e-18, 
    1.949511e-18, 1.949503e-18, 1.94943e-18, 1.949613e-18, 1.9494e-18, 
    1.949367e-18, 1.949457e-18, 1.948915e-18, 1.94907e-18, 1.948912e-18, 
    1.949012e-18, 1.951559e-18, 1.951433e-18, 1.951501e-18, 1.951374e-18, 
    1.951466e-18, 1.951067e-18, 1.950947e-18, 1.950382e-18, 1.950608e-18, 
    1.950242e-18, 1.950569e-18, 1.950512e-18, 1.95024e-18, 1.95055e-18, 
    1.949847e-18, 1.950332e-18, 1.949428e-18, 1.949921e-18, 1.949397e-18, 
    1.949488e-18, 1.949335e-18, 1.9492e-18, 1.949027e-18, 1.948714e-18, 
    1.948785e-18, 1.94852e-18, 1.951244e-18, 1.951083e-18, 1.951093e-18, 
    1.950922e-18, 1.950797e-18, 1.950519e-18, 1.950081e-18, 1.950244e-18, 
    1.949939e-18, 1.94988e-18, 1.95034e-18, 1.950062e-18, 1.950972e-18, 
    1.95083e-18, 1.950911e-18, 1.951234e-18, 1.950213e-18, 1.950739e-18, 
    1.949764e-18, 1.950047e-18, 1.94922e-18, 1.949636e-18, 1.948826e-18, 
    1.948492e-18, 1.948158e-18, 1.947792e-18, 1.950991e-18, 1.9511e-18, 
    1.9509e-18, 1.950632e-18, 1.950371e-18, 1.950031e-18, 1.949994e-18, 
    1.949931e-18, 1.949764e-18, 1.949626e-18, 1.949916e-18, 1.949591e-18, 
    1.950806e-18, 1.950165e-18, 1.951146e-18, 1.950856e-18, 1.950646e-18, 
    1.950734e-18, 1.950262e-18, 1.950152e-18, 1.949709e-18, 1.949936e-18, 
    1.948578e-18, 1.949178e-18, 1.9475e-18, 1.94797e-18, 1.95114e-18, 
    1.950989e-18, 1.950472e-18, 1.950717e-18, 1.950006e-18, 1.949833e-18, 
    1.949688e-18, 1.949511e-18, 1.949489e-18, 1.949384e-18, 1.949557e-18, 
    1.949389e-18, 1.95003e-18, 1.949742e-18, 1.950526e-18, 1.950338e-18, 
    1.950423e-18, 1.950519e-18, 1.950222e-18, 1.949912e-18, 1.949898e-18, 
    1.949801e-18, 1.949538e-18, 1.950003e-18, 1.948514e-18, 1.949444e-18, 
    1.950825e-18, 1.950546e-18, 1.950497e-18, 1.950607e-18, 1.94985e-18, 
    1.950125e-18, 1.949385e-18, 1.949583e-18, 1.949257e-18, 1.94942e-18, 
    1.949444e-18, 1.949652e-18, 1.949783e-18, 1.950114e-18, 1.950381e-18, 
    1.95059e-18, 1.950541e-18, 1.950312e-18, 1.949892e-18, 1.94949e-18, 
    1.949579e-18, 1.949282e-18, 1.950057e-18, 1.949735e-18, 1.949862e-18, 
    1.949531e-18, 1.95025e-18, 1.949659e-18, 1.950404e-18, 1.950337e-18, 
    1.950131e-18, 1.949719e-18, 1.949617e-18, 1.949521e-18, 1.949579e-18, 
    1.94988e-18, 1.949926e-18, 1.950134e-18, 1.950195e-18, 1.950351e-18, 
    1.950484e-18, 1.950364e-18, 1.95024e-18, 1.949877e-18, 1.949553e-18, 
    1.9492e-18, 1.94911e-18, 1.948716e-18, 1.949047e-18, 1.948511e-18, 
    1.948981e-18, 1.94816e-18, 1.949614e-18, 1.948981e-18, 1.950119e-18, 
    1.949994e-18, 1.949776e-18, 1.949263e-18, 1.949532e-18, 1.949214e-18, 
    1.949927e-18, 1.950307e-18, 1.950397e-18, 1.950579e-18, 1.950393e-18, 
    1.950408e-18, 1.95023e-18, 1.950287e-18, 1.949864e-18, 1.950091e-18, 
    1.949447e-18, 1.949214e-18, 1.94855e-18, 1.948149e-18, 1.94773e-18, 
    1.947549e-18, 1.947493e-18, 1.94747e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  2.08774e-25, 2.747033e-26, 3.626074e-25, 1.373513e-25, 3.735955e-25, 
    1.263632e-25, -1.593273e-25, -2.142678e-25, 3.681014e-25, 1.318573e-25, 
    -3.021726e-25, 2.08774e-25, -8.790471e-26, -1.15375e-25, -8.790471e-26, 
    -2.582202e-25, -2.032797e-25, 2.14268e-25, 2.252561e-25, -2.417381e-25, 
    1.648223e-26, -3.845834e-25, -4.944636e-26, -1.318571e-25, -1.483393e-25, 
    -4.120536e-25, -8.241066e-26, 6.592868e-26, 1.153751e-25, -2.747024e-25, 
    4.724883e-25, 2.637145e-25, -1.043869e-25, 2.582204e-25, 3.845843e-26, 
    -1.977857e-25, -2.142678e-25, 5.494135e-27, 3.626074e-25, -1.15375e-25, 
    -1.20869e-25, -6.592851e-26, -1.098801e-26, 5.494135e-27, 1.04387e-25, 
    -4.065596e-25, 9.339893e-26, -8.790471e-26, 1.098819e-26, 1.758097e-25, 
    -3.790893e-25, -8.790471e-26, 3.845835e-25, 2.692085e-25, -3.241488e-25, 
    1.867978e-25, -8.790471e-26, -2.197611e-26, 6.373098e-25, 6.263217e-25, 
    8.590255e-32, 8.241083e-26, 1.153751e-25, -1.813035e-25, -1.483393e-25, 
    -1.758095e-25, -3.076667e-25, -1.20869e-25, 4.175479e-25, 3.18655e-25, 
    -2.527262e-25, -1.373511e-25, -5.384167e-25, 4.999586e-25, -1.922916e-25, 
    2.801966e-25, -2.142678e-25, 2.417383e-25, -2.142678e-25, 2.801966e-25, 
    -5.494041e-26, -7.691661e-26, 4.395241e-25, -4.615001e-25, -4.395231e-26, 
    -1.263631e-25, 6.043463e-26, 3.461252e-25, 1.538335e-25, 5.494135e-27, 
    -1.428452e-25, 2.637145e-25, -4.175477e-25, -4.834763e-25, -3.955715e-25, 
    8.241083e-26, 3.790895e-25, -1.098801e-26, 8.790488e-26, -3.021726e-25, 
    1.428454e-25, 2.417383e-25, -2.747016e-26, 8.790488e-26, -3.681012e-25, 
    2.801966e-25, -1.373511e-25, -1.318571e-25, 2.747033e-26, -1.703155e-25, 
    -1.813035e-25, 1.977859e-25, 3.406311e-25, 2.14268e-25, 3.351371e-25, 
    3.021728e-25, -5.384167e-25, 1.428454e-25, -4.120536e-25, 8.241083e-26, 
    -1.593273e-25, -9.88928e-26, 2.527264e-25, 8.590077e-32, 1.703156e-25, 
    2.747033e-26, 2.032799e-25, 1.648216e-25, -3.186548e-25, 4.615002e-25, 
    2.747033e-26, -2.966786e-25, -2.856905e-25, -1.098801e-26, -9.88928e-26, 
    -2.637143e-25, -9.339876e-26, 1.648216e-25, -2.637143e-25, 1.098811e-25, 
    1.263632e-25, -6.592851e-26, 1.758097e-25, -1.538333e-25, -2.637143e-25, 
    -1.648206e-26, -1.648214e-25, -9.88928e-26, -4.944636e-26, -1.098801e-26, 
    -2.197619e-25, 4.3403e-25, 2.637145e-25, -1.648206e-26, 1.867978e-25, 
    -1.043869e-25, -3.296421e-26, -3.241488e-25, -5.054525e-25, 1.648223e-26, 
    1.04387e-25, -1.318571e-25, -4.010655e-25, -3.296429e-25, -9.88928e-26, 
    6.043463e-26, -5.65887e-25, -5.494041e-26, -3.845826e-26, -2.197619e-25, 
    -5.933573e-25, -6.592851e-26, 2.14268e-25, -5.933573e-25, 1.758097e-25, 
    5.329229e-25, 3.955717e-25, 2.197621e-25, -5.164406e-25, -1.813035e-25, 
    2.197628e-26, -2.417381e-25, -3.241488e-25, 2.08774e-25, -3.351369e-25, 
    -1.648214e-25, -6.592851e-26, -4.50512e-25, 1.04387e-25, -5.60393e-25, 
    -1.648206e-26, -3.021726e-25, -1.813035e-25, -1.648206e-26, 
    -4.779822e-25, 1.428454e-25, 2.417383e-25, 1.483394e-25, 2.362442e-25, 
    7.691678e-26, -3.845826e-26, -5.493964e-27, -1.922916e-25, -1.043869e-25, 
    -6.482978e-25, 9.339893e-26, -2.417381e-25, -3.296421e-26, -5.054525e-25, 
    -3.296421e-26, 9.889298e-26, -2.197611e-26, -1.263631e-25, 2.197628e-26, 
    -3.131607e-25, -1.15375e-25, -2.087738e-25, -2.032797e-25, -1.648214e-25, 
    2.801966e-25, -9.339876e-26, 6.208277e-25, 1.318573e-25, -1.098809e-25, 
    -2.3075e-25, -3.296421e-26, 3.131609e-25, -5.493964e-27, 2.747033e-26, 
    -1.813035e-25, -3.626072e-25, 4.999586e-25, 6.043463e-26, 1.263632e-25, 
    -3.021726e-25, -8.241066e-26, 2.197628e-26, 5.494135e-27, 2.966788e-25, 
    2.252561e-25, 6.043463e-26, 1.593275e-25, -2.747016e-26, 4.779824e-25, 
    -1.098809e-25, 1.373513e-25, 8.590102e-32, 4.065598e-25, 3.24149e-25, 
    1.538335e-25, -5.164406e-25, -7.691661e-26, 1.648223e-26, -5.878632e-25, 
    -4.395231e-26, 1.867978e-25, -8.790471e-26, -4.944644e-25, -9.88928e-26, 
    -9.88928e-26, -1.483393e-25, 3.461252e-25, -1.098801e-26, -2.692083e-25, 
    4.395248e-26, -9.339876e-26, 8.790488e-26, -6.263215e-25, -4.50512e-25, 
    6.592868e-26, -2.032797e-25, 3.681014e-25, -1.263631e-25, -1.098801e-26, 
    -8.790471e-26, -1.867976e-25, 2.692085e-25, -2.142678e-25, 8.241083e-26, 
    1.758097e-25, 8.790488e-26, 8.590033e-32, 1.153751e-25, -5.494041e-26, 
    -1.373511e-25, 1.593275e-25, 4.395248e-26, -4.395231e-26, -3.790893e-25, 
    -1.098809e-25, -5.164406e-25, -3.186548e-25, -8.241066e-26, 
    -2.747016e-26, -2.142678e-25, -8.241074e-25, -1.20869e-25, 8.790488e-26, 
    -2.36244e-25, -7.691661e-26, -1.648206e-26, 2.911847e-25, 3.790895e-25, 
    -3.900774e-25, 2.637145e-25, -2.36244e-25, -2.417381e-25, -4.944636e-26, 
    -4.395231e-26, -1.318571e-25, 4.615002e-25, -3.241488e-25, 2.032799e-25, 
    -2.966786e-25, 7.142273e-26, -3.571131e-25, -1.703155e-25, 1.648223e-26, 
    -7.142256e-26, -8.241066e-26, -1.20869e-25, -3.900774e-25, -3.845826e-26, 
    3.626074e-25, 1.977859e-25, 2.472323e-25, -2.747024e-25, -2.36244e-25, 
    8.241083e-26, 5.988515e-25, -5.823692e-25, 1.318573e-25, 1.648216e-25, 
    -2.087738e-25, -3.626072e-25, 5.109467e-25, 1.098819e-26, -9.88928e-26 ;

 M_LITR2C_TO_LEACHING =
  2.692085e-25, 1.538334e-25, -3.296424e-26, -1.428452e-25, -1.098809e-25, 
    5.494055e-26, -6.592854e-26, -1.703155e-25, 2.801966e-25, -2.747024e-25, 
    -1.15375e-25, 5.494105e-27, -1.867976e-25, 2.307501e-25, -4.944639e-26, 
    -1.648214e-25, 1.208691e-25, 3.351371e-25, 1.098811e-25, -1.758095e-25, 
    -1.373512e-25, -2.197619e-25, -2.087738e-25, 5.562049e-32, -1.318571e-25, 
    -3.296424e-26, -2.637143e-25, 1.922918e-25, 5.562085e-32, 7.691675e-26, 
    2.197625e-26, -2.747019e-26, -3.790894e-25, -2.911846e-25, -1.15375e-25, 
    1.263632e-25, -5.493994e-27, -4.230417e-25, -2.582203e-25, -1.043869e-25, 
    -3.845829e-26, -2.582203e-25, 3.296435e-26, -5.493994e-27, 3.296435e-26, 
    -5.494044e-26, -1.813036e-25, -5.494044e-26, 1.703156e-25, 5.56206e-32, 
    -3.296424e-26, 1.428453e-25, 1.64822e-26, -2.197614e-26, 9.33989e-26, 
    -3.955715e-25, -1.043869e-25, 1.04387e-25, -2.197619e-25, 5.494105e-27, 
    -1.648214e-25, 9.889295e-26, 6.592865e-26, 2.087739e-25, 2.472323e-25, 
    5.494055e-26, 3.296435e-26, -9.889284e-26, -1.538333e-25, -8.790474e-26, 
    -2.637143e-25, -1.043869e-25, -7.691664e-26, 1.208691e-25, 2.74703e-26, 
    6.592865e-26, 1.483394e-25, -8.241069e-26, 2.087739e-25, -2.747024e-25, 
    5.494055e-26, 2.74703e-26, 6.04346e-26, 1.208691e-25, -4.120537e-25, 
    9.889295e-26, 6.04346e-26, -1.922917e-25, 1.04387e-25, -2.911846e-25, 
    -9.339879e-26, 1.867977e-25, 2.14268e-25, -3.296424e-26, -2.197619e-25, 
    -1.648214e-25, -9.889284e-26, -2.472322e-25, -1.758095e-25, 1.318572e-25, 
    -4.395234e-26, 2.197625e-26, 1.098815e-26, -1.043869e-25, -7.691664e-26, 
    -1.867976e-25, -1.648209e-26, 4.010657e-25, -2.637143e-25, -1.648214e-25, 
    -9.339879e-26, 2.307501e-25, 3.84584e-26, 1.208691e-25, 6.592865e-26, 
    2.307501e-25, -3.626072e-25, 3.29643e-25, 2.307501e-25, 1.593275e-25, 
    1.098815e-26, 1.373513e-25, 2.527263e-25, 2.032799e-25, 6.592865e-26, 
    1.593275e-25, -6.373097e-25, -1.318571e-25, 1.04387e-25, -3.296424e-26, 
    2.307501e-25, 1.648215e-25, 1.977858e-25, -1.098804e-26, -9.339879e-26, 
    1.098815e-26, -1.703155e-25, -2.527262e-25, -1.373512e-25, 1.098815e-26, 
    -3.845829e-26, 8.24108e-26, 2.856906e-25, 5.494055e-26, -1.098809e-25, 
    1.483394e-25, 7.14227e-26, 2.197625e-26, -1.098809e-25, 4.395245e-26, 
    -3.845829e-26, -2.637143e-25, -1.538333e-25, 1.867977e-25, -2.25256e-25, 
    -2.25256e-25, 1.318572e-25, -3.845829e-26, -4.340298e-25, -1.703155e-25, 
    3.461252e-25, -2.142679e-25, -3.845829e-26, 2.74703e-26, -9.339879e-26, 
    6.04346e-26, 1.593275e-25, -1.263631e-25, -6.043449e-26, -1.428452e-25, 
    1.813037e-25, 6.592865e-26, 9.889295e-26, -1.15375e-25, -1.428452e-25, 
    -1.593274e-25, 2.74703e-26, -2.3075e-25, -4.395234e-26, -2.801965e-25, 
    1.703156e-25, -2.362441e-25, 3.296435e-26, 1.483394e-25, -5.494044e-26, 
    -9.339879e-26, -3.076667e-25, 7.691675e-26, 7.14227e-26, 1.373513e-25, 
    -3.516191e-25, -2.197619e-25, 6.04346e-26, -1.263631e-25, -2.582203e-25, 
    9.33989e-26, 1.428453e-25, -5.493994e-27, 2.14268e-25, -1.15375e-25, 
    -7.142259e-26, -6.043449e-26, 2.74703e-26, 1.813037e-25, 2.307501e-25, 
    2.087739e-25, -2.142679e-25, -2.747024e-25, -4.450179e-25, -5.493994e-27, 
    -8.241069e-26, -1.428452e-25, -8.790474e-26, 8.24108e-26, -1.977857e-25, 
    2.801966e-25, -4.395234e-26, -3.845829e-26, -1.648209e-26, 2.252561e-25, 
    1.263632e-25, 2.74703e-26, 2.692085e-25, -2.142679e-25, -2.747019e-26, 
    -2.747019e-26, 1.098811e-25, -1.20869e-25, -6.592854e-26, -3.461251e-25, 
    2.362442e-25, 1.263632e-25, 1.208691e-25, -2.637143e-25, 7.691675e-26, 
    1.098811e-25, -2.3075e-25, -5.384168e-25, 2.582204e-25, -9.339879e-26, 
    -1.428452e-25, 1.64822e-26, -3.735953e-25, -1.263631e-25, 5.494105e-27, 
    3.84584e-26, -2.197619e-25, -1.098804e-26, 1.64822e-26, -1.098804e-26, 
    3.84584e-26, -3.845829e-26, -5.494044e-26, -1.15375e-25, 1.64822e-26, 
    1.098811e-25, -2.966786e-25, 3.735954e-25, 1.703156e-25, 5.494055e-26, 
    -7.691664e-26, -9.889284e-26, -3.021727e-25, -7.691664e-26, 1.648215e-25, 
    -5.493994e-27, -2.747019e-26, 1.703156e-25, -4.065596e-25, -1.20869e-25, 
    -1.648209e-26, -2.032798e-25, -1.593274e-25, -5.493994e-27, 
    -7.691664e-26, 3.296435e-26, -1.538333e-25, -1.428452e-25, 9.889295e-26, 
    -3.516191e-25, -1.043869e-25, 8.24108e-26, 9.889295e-26, 6.04346e-26, 
    -1.098809e-25, -6.592854e-26, 1.318572e-25, 7.691675e-26, 4.94465e-26, 
    7.691675e-26, -2.747019e-26, -1.593274e-25, 1.593275e-25, -1.098804e-26, 
    -1.428452e-25, -1.922917e-25, 8.790485e-26, 2.087739e-25, -7.142259e-26, 
    -8.241069e-26, 5.494105e-27, -1.813036e-25, 1.977858e-25, -2.197614e-26, 
    2.307501e-25, 1.373513e-25, -2.856905e-25, -1.318571e-25, 1.64822e-26, 
    -8.790474e-26, 5.56205e-32, -1.15375e-25, -3.296424e-26, -1.593274e-25, 
    6.592865e-26, -3.735953e-25, 3.84584e-26, -7.142259e-26, -2.197619e-25, 
    1.098815e-26, -2.197614e-26, -7.691664e-26, -1.043869e-25, -2.582203e-25, 
    1.538334e-25, -3.296424e-26, 1.098815e-26, -3.296424e-26, 3.84584e-26, 
    -1.098809e-25, -2.472322e-25, 1.373513e-25, -3.021727e-25, -7.142259e-26, 
    3.296435e-26, 2.472323e-25, 5.494055e-26, 2.527263e-25 ;

 M_LITR3C_TO_LEACHING =
  2.747028e-26, -1.263631e-25, 3.845837e-26, 6.31816e-26, -1.09881e-25, 
    6.867565e-26, -3.296427e-26, -1.15375e-25, -1.071339e-25, -6.318154e-26, 
    -2.19762e-25, -1.400982e-25, -6.592857e-26, 2.747052e-27, 4.12054e-26, 
    4.395242e-26, -8.790477e-26, -2.746997e-27, 3.02173e-26, -1.483393e-25, 
    -2.747022e-26, -4.395237e-26, -7.691667e-26, -1.098807e-26, 
    -8.241047e-27, -4.395237e-26, 3.845837e-26, -9.614584e-26, 1.04387e-25, 
    -5.494022e-27, -1.428453e-25, 2.781044e-32, -6.043452e-26, -2.170149e-25, 
    1.730626e-25, -3.296427e-26, 2.472325e-26, -7.416964e-26, -1.098807e-26, 
    -4.395237e-26, -1.648212e-26, -8.241047e-27, 1.92292e-26, -2.747022e-26, 
    1.813037e-25, 8.241077e-26, 1.538334e-25, -8.515774e-26, 8.241077e-26, 
    2.747052e-27, -1.208691e-25, -1.620744e-25, -2.47232e-26, 4.12054e-26, 
    1.153751e-25, 1.373515e-26, 4.12054e-26, 1.153751e-25, -5.494022e-27, 
    6.31816e-26, -5.494022e-27, -7.691667e-26, 1.92292e-26, 5.21935e-26, 
    6.043457e-26, -3.021725e-26, 3.571135e-26, -9.339881e-26, 1.07134e-25, 
    -1.895447e-25, 5.21935e-26, 1.648218e-26, 1.483394e-25, 8.241102e-27, 
    2.472325e-26, -8.790477e-26, -5.219344e-26, -1.09881e-25, 3.571135e-26, 
    -9.339881e-26, 2.781044e-32, -1.37351e-26, -6.043452e-26, -3.845832e-26, 
    4.395242e-26, -3.296427e-26, 1.620745e-25, -3.845832e-26, 1.016399e-25, 
    -4.395237e-26, 2.747052e-27, 8.515779e-26, 4.12054e-26, -8.241071e-26, 
    -4.395237e-26, -6.318154e-26, 1.92292e-26, -3.021725e-26, -1.071339e-25, 
    1.04387e-25, -1.18122e-25, -3.845832e-26, 3.845837e-26, -3.845832e-26, 
    9.065185e-26, 7.966375e-26, -3.57113e-26, -1.922915e-26, 9.065185e-26, 
    -4.395237e-26, -1.071339e-25, 2.747052e-27, -1.236161e-25, -1.18122e-25, 
    -4.120535e-26, -9.065179e-26, -4.944642e-26, 2.747028e-26, 2.781031e-32, 
    -1.373512e-25, 1.236161e-25, 2.197623e-26, -2.746997e-27, -7.142262e-26, 
    1.236161e-25, -1.098807e-26, -1.318572e-25, -4.669939e-26, -2.47232e-26, 
    -1.37351e-26, -1.565804e-25, 6.867565e-26, 1.648218e-26, -5.768749e-26, 
    -8.515774e-26, -1.346042e-25, 3.571135e-26, -8.241071e-26, 2.747052e-27, 
    1.758096e-25, 4.669945e-26, 2.781037e-32, -2.115209e-25, -4.120535e-26, 
    8.515779e-26, 1.04387e-25, -2.747022e-26, -6.043452e-26, -6.318154e-26, 
    -7.966369e-26, -6.592857e-26, -9.614584e-26, 1.098813e-26, 8.790482e-26, 
    2.747028e-26, -6.043452e-26, -6.592857e-26, -2.47232e-26, 7.691672e-26, 
    1.291102e-25, 1.098813e-26, 1.098813e-26, -9.065179e-26, 4.12054e-26, 
    -1.977858e-25, 6.592862e-26, -9.339881e-26, -9.614584e-26, -2.747022e-26, 
    -1.675685e-25, 7.416969e-26, -4.395237e-26, -1.648215e-25, 1.92292e-26, 
    -2.197617e-26, 1.09881e-25, 3.02173e-26, -8.241047e-27, -9.339881e-26, 
    -9.889287e-26, 4.395242e-26, -1.648212e-26, -1.263631e-25, -3.57113e-26, 
    -1.648212e-26, -5.494022e-27, -1.098807e-26, 5.21935e-26, 1.318572e-25, 
    -1.291101e-25, -2.005328e-25, -1.455923e-25, -8.241047e-27, 
    -2.747022e-26, -1.016399e-25, -8.241047e-27, -6.592857e-26, 
    -1.291101e-25, -2.197617e-26, 3.571135e-26, 6.043457e-26, -3.57113e-26, 
    -7.416964e-26, 2.197623e-26, 8.515779e-26, -1.37351e-26, -1.15375e-25, 
    -1.263631e-25, 4.944647e-26, 5.494053e-26, 8.241102e-27, 1.620745e-25, 
    4.669945e-26, -5.494047e-26, 1.12628e-25, -3.845832e-26, -1.428453e-25, 
    7.416969e-26, -6.592857e-26, 2.747052e-27, 1.373515e-26, -7.142262e-26, 
    -1.263631e-25, -1.09881e-25, 1.07134e-25, -4.120535e-26, -1.043869e-25, 
    -8.515774e-26, 8.790482e-26, -1.648212e-26, 1.318572e-25, 1.181221e-25, 
    -2.747022e-26, 4.944647e-26, -1.016399e-25, 3.845837e-26, -8.515774e-26, 
    2.197623e-26, 4.944647e-26, -1.043869e-25, -2.170149e-25, -6.043452e-26, 
    6.592862e-26, -6.043452e-26, 9.339887e-26, -4.120535e-26, 4.944647e-26, 
    -6.592857e-26, 6.592862e-26, 6.043457e-26, -8.241047e-27, 5.494077e-27, 
    -1.922915e-26, -7.691667e-26, 9.614589e-26, -1.15375e-25, -3.296427e-26, 
    -2.47232e-26, -1.37351e-26, -5.494022e-27, -3.021725e-26, -1.346042e-25, 
    -4.669939e-26, 1.648218e-26, -5.768749e-26, -8.241047e-27, 4.944647e-26, 
    -1.538334e-25, -8.241047e-27, 4.669945e-26, 4.395242e-26, -7.142262e-26, 
    -2.032798e-25, 7.966375e-26, -3.296427e-26, 1.208691e-25, -9.065179e-26, 
    8.790482e-26, 8.515779e-26, 2.781028e-32, -6.592857e-26, 5.494053e-26, 
    -4.120535e-26, -4.944642e-26, -1.37351e-26, 1.648218e-26, 6.31816e-26, 
    -6.318154e-26, -8.241071e-26, -1.043869e-25, -3.845832e-26, 
    -7.966369e-26, 4.12054e-26, -5.768749e-26, 3.571135e-26, 1.263632e-25, 
    -1.318572e-25, -1.09881e-25, 7.966375e-26, 1.510864e-25, -9.614584e-26, 
    -6.318154e-26, -1.922915e-26, -3.845832e-26, -1.15375e-25, -9.065179e-26, 
    -6.592857e-26, 1.373515e-26, -9.614584e-26, -6.592857e-26, 3.02173e-26, 
    -1.400982e-25, 2.472325e-26, 1.373513e-25, -1.922915e-26, 1.291102e-25, 
    -7.691667e-26, -3.57113e-26, 8.241077e-26, 1.785566e-25, -8.241047e-27, 
    4.395242e-26, -8.241047e-27, 2.197623e-26, -1.236161e-25, 1.648218e-26, 
    4.12054e-26, 2.747052e-27, 5.768755e-26, -1.813036e-25, -3.845832e-26, 
    4.669945e-26, -5.768749e-26, -2.47232e-26, -1.12628e-25, 1.098813e-26, 
    -1.236161e-25, 3.845837e-26 ;

 M_SOIL1C_TO_LEACHING =
  -2.299818e-20, 1.964273e-20, -1.736818e-21, 3.479114e-20, -4.149414e-20, 
    7.574352e-21, 1.166661e-20, 1.640348e-20, 8.18336e-21, 1.325442e-20, 
    -1.442944e-20, -4.522789e-20, -3.696816e-20, 1.113988e-20, -1.372939e-20, 
    1.877064e-21, 8.317385e-21, -4.730668e-21, -1.283609e-21, -2.969226e-21, 
    -2.391365e-20, 3.795937e-21, -5.380928e-21, 4.032192e-20, 7.337154e-21, 
    -7.616728e-22, 4.475261e-20, 8.869545e-21, -1.492169e-20, 1.051815e-20, 
    1.676857e-21, 5.7776e-21, -1.072737e-20, 4.055433e-20, -3.782401e-20, 
    4.019809e-20, 3.039469e-20, -1.75279e-20, 5.344452e-21, -1.072963e-20, 
    -2.395266e-20, 3.423444e-20, 3.903387e-21, -2.782631e-21, -6.36523e-20, 
    -5.816349e-21, -4.286193e-21, 2.084602e-20, -1.083197e-20, -1.273618e-20, 
    2.958411e-20, -4.133098e-20, 3.702897e-20, 6.928016e-21, 5.105261e-21, 
    7.064201e-20, 2.684275e-20, 2.25761e-21, 5.351807e-21, 2.071908e-20, 
    -3.569645e-20, -5.105833e-21, -2.915407e-20, -2.73675e-20, 7.491557e-23, 
    -1.517672e-20, 3.726702e-20, 2.627125e-21, 7.082126e-21, -1.136041e-20, 
    -7.761519e-21, -8.675023e-21, -9.963441e-21, -1.10231e-20, -6.764901e-21, 
    5.651226e-21, -1.452418e-20, 1.91471e-20, 9.99821e-21, -3.678036e-21, 
    1.742244e-20, 1.029845e-20, -2.884729e-20, -2.359332e-20, 3.325485e-21, 
    -7.602061e-21, -6.33515e-21, 6.989396e-21, 2.432559e-20, -1.060157e-20, 
    -5.366226e-21, 3.383494e-20, 2.13917e-20, 3.048149e-20, -1.213056e-20, 
    -4.939732e-20, 1.057753e-20, 7.44769e-21, 1.91143e-20, 7.039908e-22, 
    -1.478453e-20, 6.397909e-21, 1.440373e-20, -3.375466e-20, 3.432861e-20, 
    1.046615e-20, -8.233137e-22, 4.419421e-20, 2.980124e-20, 1.856749e-20, 
    -1.488271e-21, -3.033129e-21, 8.186756e-21, -1.356571e-20, 6.537583e-21, 
    -6.916448e-21, 6.770838e-21, -1.584396e-20, 1.509953e-20, 1.279723e-20, 
    -5.336034e-20, 1.326846e-21, -3.399245e-20, -1.664662e-20, -1.42516e-20, 
    -2.715628e-20, 1.208945e-21, -2.679183e-20, -2.791964e-21, -2.252884e-20, 
    8.529412e-21, -6.342783e-20, 1.192502e-20, -1.40274e-20, -7.011741e-21, 
    3.223277e-22, 7.308588e-21, -8.037187e-21, -1.63193e-21, -3.009301e-20, 
    -1.619115e-20, -1.489144e-20, -2.580655e-20, -4.734243e-20, 
    -5.731209e-20, 1.632996e-20, -2.745541e-20, 1.50616e-20, 1.416679e-20, 
    -5.018466e-21, -5.054937e-21, 4.709457e-21, -3.303796e-20, 4.274325e-21, 
    -1.548998e-20, -1.450635e-20, -1.557535e-20, 8.236075e-22, 7.015399e-21, 
    3.00489e-20, -1.730908e-20, -3.417708e-20, 1.769042e-21, 3.956565e-20, 
    -9.381292e-21, -3.507466e-23, -1.180117e-21, -1.899358e-20, 
    -1.529092e-20, -1.692436e-21, 1.246844e-21, -3.894306e-20, 5.481584e-20, 
    -5.640776e-21, -2.459586e-20, -1.240254e-20, 2.463011e-20, -3.171223e-20, 
    -3.563683e-20, -1.533618e-20, -3.485307e-20, 2.064726e-20, 8.548362e-21, 
    8.205967e-21, -1.504353e-20, -5.971127e-22, 1.633048e-21, 5.49818e-20, 
    8.252055e-21, -1.676822e-20, 1.131432e-20, 2.556565e-20, -2.569119e-20, 
    -1.282607e-20, 1.463413e-20, 1.453746e-20, 7.752581e-22, -1.55756e-21, 
    -8.548378e-21, 2.298827e-20, -2.504174e-20, 6.279436e-21, -9.099404e-21, 
    -1.789064e-20, 1.314586e-20, -1.880785e-20, -9.238506e-21, 4.088847e-21, 
    -5.846294e-21, -5.253411e-21, 1.094183e-22, -1.728388e-20, 3.671372e-20, 
    -8.131249e-22, 3.346287e-20, 4.526208e-20, 4.038808e-21, 1.466524e-20, 
    9.569316e-21, 9.449726e-21, -4.295246e-20, 6.515237e-21, -1.892317e-20, 
    2.693913e-20, 6.170884e-21, 1.977532e-20, -4.848569e-21, -3.861545e-21, 
    1.921919e-20, -8.340538e-21, -2.950719e-20, 2.026218e-20, 9.091215e-21, 
    1.944651e-20, 2.462218e-20, -3.296918e-21, -1.889207e-20, -3.516179e-20, 
    3.072975e-20, 9.980112e-21, -2.088195e-20, -1.120661e-20, 2.22348e-20, 
    6.077036e-21, -1.165897e-20, 9.779653e-21, 3.530123e-20, 2.092464e-20, 
    1.690219e-20, -3.37052e-20, -1.639878e-22, 4.207855e-20, 1.919755e-21, 
    -5.388833e-21, 7.69622e-21, -9.760703e-21, -3.343862e-21, -1.538365e-20, 
    -2.235694e-20, -1.412635e-20, -1.893251e-20, 1.961312e-21, 1.929043e-20, 
    1.479361e-20, 1.436583e-20, -3.296165e-22, -2.828728e-21, -1.285832e-20, 
    3.225789e-20, 7.862176e-21, -2.066483e-21, 5.462091e-21, 1.032082e-20, 
    -1.228467e-21, -1.169516e-20, 2.506945e-20, -4.332793e-20, 1.364911e-20, 
    -2.536363e-21, 3.435858e-20, -4.389963e-21, 1.763678e-21, -1.353857e-20, 
    -7.263363e-22, 2.415949e-21, 2.302192e-20, -1.986779e-20, -1.968598e-20, 
    -2.473723e-20, -7.468608e-21, -1.541364e-20, -6.176791e-20, 
    -3.644961e-21, -2.567903e-20, -1.175027e-20, -1.130216e-20, 
    -8.026164e-21, -1.591208e-20, -2.563974e-20, -3.439448e-20, 
    -2.452266e-20, 1.336017e-20, -3.045123e-20, 2.677433e-21, -5.829623e-21, 
    1.016756e-20, 3.438299e-21, -2.15568e-20, -2.447291e-20, 3.824528e-20, 
    3.779969e-20, 2.468494e-20, 6.885064e-21, -8.145461e-21, -8.423407e-21, 
    -8.673333e-21, 7.733825e-21, 2.42928e-20, -2.353961e-20, 1.727911e-20, 
    1.747672e-20, -8.955793e-21, 2.825298e-20, 7.200026e-21, 1.884118e-21, 
    -8.932875e-21, 2.543419e-20, -4.139462e-20, 6.453641e-20, -5.585634e-21, 
    -2.687979e-20, -4.436582e-20, -1.923617e-20, 2.541495e-20, -1.057582e-20, 
    -5.999369e-22, 4.063694e-21, -3.313327e-21 ;

 M_SOIL2C_TO_LEACHING =
  -4.493445e-21, 9.829709e-21, 1.426996e-20, -5.448506e-21, 2.907576e-20, 
    -5.083507e-22, 4.600039e-21, 4.304688e-20, -4.773627e-21, -1.910684e-21, 
    4.384861e-21, -3.636651e-20, 4.642297e-20, -2.873961e-20, 1.082856e-21, 
    -1.070531e-20, -6.8616e-21, 1.945102e-20, -2.609598e-21, 2.896152e-20, 
    -3.985356e-21, 1.251847e-20, 6.944704e-21, -9.71238e-21, 3.028698e-20, 
    -4.10268e-20, -9.006673e-21, 4.3467e-21, -5.048891e-20, 2.453424e-20, 
    1.937159e-20, 3.154314e-20, 2.766532e-21, -3.02321e-20, -1.691889e-20, 
    9.466968e-21, 2.034843e-20, 1.208986e-20, 3.153747e-20, -1.002618e-20, 
    -3.108964e-20, 5.055224e-20, -8.737781e-21, -1.90931e-20, -1.332341e-20, 
    -1.986779e-20, 2.828043e-20, 1.779231e-21, -1.928931e-20, -8.829132e-21, 
    -6.563586e-21, 2.761856e-20, -1.588552e-20, 1.327081e-20, 2.627361e-20, 
    4.108106e-20, 2.43219e-20, 1.557764e-20, -5.809552e-20, -2.544238e-20, 
    -1.717731e-20, 3.507642e-20, -1.414587e-20, 1.417811e-20, -6.514345e-20, 
    -4.253091e-20, -2.189777e-20, 9.084707e-21, -3.538093e-20, -2.037863e-20, 
    2.231311e-20, -9.54528e-21, -1.824744e-20, 2.525605e-20, -6.948394e-21, 
    6.070789e-21, 2.677037e-20, 3.69433e-20, 1.334461e-20, -3.772505e-20, 
    -3.976905e-21, 3.504446e-20, -6.388576e-21, -1.666808e-20, 1.443595e-20, 
    1.201492e-20, 2.223028e-20, 1.217496e-20, 1.696075e-20, 1.815868e-20, 
    -1.050205e-20, -1.821464e-20, -2.278951e-20, -2.492669e-20, 
    -1.648376e-20, -2.936555e-20, -9.575797e-21, 1.761752e-20, -2.299366e-20, 
    1.295531e-20, -7.568987e-21, 1.265193e-20, -4.099314e-21, -9.886531e-21, 
    -2.696912e-20, 6.465492e-21, -4.547159e-21, 2.106515e-20, -1.009601e-20, 
    6.904292e-21, -1.401788e-21, -8.744872e-22, 1.553436e-20, -3.036644e-20, 
    -2.864883e-20, 3.290083e-20, -9.939127e-21, 1.32024e-20, -1.839305e-20, 
    -1.055573e-20, -2.182397e-20, -1.715753e-20, 9.640834e-21, -2.480481e-20, 
    -3.526219e-20, -4.588143e-21, 2.594451e-20, -1.429513e-20, -2.222009e-20, 
    -7.798845e-21, 2.84037e-20, -2.141399e-21, 1.696355e-20, 2.434327e-21, 
    1.16304e-20, 1.538196e-20, 8.660604e-21, -5.92304e-20, -4.990783e-21, 
    2.836951e-20, -3.829078e-20, -1.978947e-20, -6.731543e-21, -2.197129e-20, 
    -1.862628e-20, -7.092416e-20, 7.541555e-21, -1.939757e-20, 9.802822e-21, 
    -1.563671e-20, 2.964632e-20, 1.184981e-20, -1.925878e-20, -1.518888e-20, 
    -4.51126e-21, -1.090632e-20, 1.905689e-20, 6.480734e-21, 1.45236e-20, 
    -2.910826e-20, -1.057611e-20, -4.153797e-20, -2.74424e-20, 2.114149e-20, 
    -2.541778e-20, -2.525775e-20, -2.287094e-20, 2.354808e-20, 2.046772e-20, 
    -2.897792e-20, -1.615918e-20, -8.366559e-21, -6.364834e-21, 9.317962e-21, 
    -2.056726e-20, -1.198609e-20, 3.217556e-22, 1.27698e-20, -1.920815e-20, 
    -2.594901e-21, 3.785486e-21, -1.426348e-20, 9.082454e-21, -1.269828e-20, 
    -1.625644e-20, -4.520554e-20, -2.450881e-20, -1.976995e-20, 5.741102e-20, 
    -2.805084e-20, 1.751348e-20, -6.153014e-20, -7.883404e-21, 1.236835e-20, 
    -1.62918e-20, -2.994913e-20, 5.846321e-21, -1.781628e-20, 6.246655e-21, 
    1.303501e-20, 1.379925e-20, -1.523664e-20, 1.40568e-20, 4.171144e-21, 
    1.4337e-20, 3.798857e-20, 7.020485e-21, 1.519876e-20, -3.010801e-20, 
    5.562643e-20, 5.634966e-20, 1.529566e-21, 1.265729e-20, 3.504532e-20, 
    3.174106e-20, 2.981988e-20, -1.178817e-20, -8.205705e-21, 1.151273e-21, 
    -1.917198e-20, -3.221773e-20, -1.879481e-20, -2.892618e-20, 
    -1.382015e-20, -3.49557e-20, -5.397386e-20, -2.520487e-20, 3.916661e-21, 
    7.001552e-21, 4.340031e-20, -6.149446e-22, 2.197046e-20, -8.472302e-21, 
    8.978963e-21, -8.380143e-21, 2.178726e-21, 1.790562e-20, -4.455384e-20, 
    -3.179612e-21, -3.080635e-20, -1.868652e-20, 3.585593e-20, -2.051438e-20, 
    1.827884e-20, -2.676837e-20, 2.156613e-20, -3.350049e-20, 2.16207e-20, 
    9.510232e-21, -2.402053e-20, 1.754767e-20, -1.299543e-20, -2.360151e-20, 
    -2.636465e-20, -3.411092e-20, -3.186321e-20, 2.194839e-20, 5.389144e-21, 
    1.479926e-20, 1.584025e-20, 3.573435e-20, -3.986784e-21, -1.372799e-20, 
    9.337762e-21, 1.729407e-20, 8.618484e-21, 5.761882e-20, -1.086196e-20, 
    -2.198741e-20, 7.069527e-23, 6.383783e-21, 8.07386e-20, -3.266162e-20, 
    1.718522e-20, -1.029422e-20, -7.738339e-21, -1.484364e-20, 1.106269e-20, 
    -1.696378e-21, 3.250668e-20, 4.264147e-20, 2.874835e-20, 1.684454e-20, 
    -3.859247e-20, 4.589572e-21, -1.983499e-20, 2.226251e-20, -3.235543e-20, 
    -1.160344e-21, -9.860815e-21, 2.39818e-20, 1.615382e-20, 1.388519e-20, 
    9.644509e-21, -7.432709e-21, -4.196886e-21, -1.976713e-20, -3.637641e-20, 
    2.359925e-20, 1.911456e-20, 1.053541e-20, 9.805674e-21, 1.116843e-20, 
    -2.277171e-20, 5.408724e-20, -3.531025e-20, 5.053525e-21, 5.12053e-21, 
    -5.464631e-21, 6.264749e-21, -4.504467e-21, 2.875571e-20, -1.443905e-20, 
    3.763513e-20, 1.898527e-21, -2.188789e-20, 1.288689e-20, -1.261713e-20, 
    4.704017e-20, 1.78553e-20, 2.104054e-20, -3.649376e-20, 1.119754e-20, 
    -1.603989e-20, 2.205921e-20, 7.875216e-21, -1.675207e-20, 2.884122e-21, 
    -7.251478e-21, 1.72446e-20, 1.718242e-20, -1.672436e-20, 2.497756e-20, 
    -3.584799e-20, -1.040139e-20, 1.326233e-20, 2.446298e-20, 3.995356e-20 ;

 M_SOIL3C_TO_LEACHING =
  1.681969e-21, -2.398377e-20, 9.102228e-21, 1.592481e-20, -1.622082e-20, 
    7.910821e-21, 2.353309e-20, -8.085175e-23, -8.055564e-21, 2.962172e-21, 
    1.112093e-20, -1.133327e-20, 2.706752e-20, 8.501719e-21, -6.103012e-21, 
    6.979207e-21, -9.411827e-21, -1.709249e-20, 2.97328e-20, -1.189902e-20, 
    3.802729e-21, -2.671805e-20, 1.265136e-20, 2.978739e-20, 3.338187e-21, 
    -4.703792e-21, 5.015053e-21, 3.955365e-22, -3.954187e-20, 1.661074e-20, 
    3.007322e-20, 8.444046e-21, -1.253006e-20, -1.521121e-20, 2.557301e-20, 
    4.558466e-21, 2.000035e-21, 8.927218e-21, -1.506642e-20, 5.234201e-21, 
    1.636558e-20, 1.2739e-20, 2.609295e-20, -2.376438e-20, -3.730832e-20, 
    9.499193e-21, -1.901873e-20, 3.623816e-20, -1.127867e-20, -2.049543e-20, 
    -1.03259e-20, -1.024953e-20, -8.627791e-21, 8.045375e-21, -2.361001e-20, 
    1.791044e-20, 1.486202e-20, 3.609603e-21, -3.157002e-20, 9.914813e-21, 
    2.238097e-20, -8.85796e-21, 1.316338e-20, -7.932299e-21, -2.906468e-21, 
    1.247718e-20, 7.958587e-21, 1.143165e-20, -1.902695e-20, 1.91259e-20, 
    2.404338e-21, 3.20187e-20, -1.490811e-20, 1.42352e-20, -3.181484e-20, 
    3.010632e-20, -1.5392e-21, -5.026966e-21, -1.754627e-20, -4.085348e-20, 
    2.174456e-20, -2.869943e-20, -2.418648e-20, 1.651799e-20, -2.10168e-20, 
    -7.315926e-21, -1.475431e-20, 2.083498e-20, 1.73806e-20, 3.610331e-20, 
    1.115826e-20, 5.021863e-21, -2.39671e-20, -2.095744e-20, 1.873684e-20, 
    -2.250707e-20, -8.014579e-21, 1.939702e-20, -1.843377e-20, 2.339654e-20, 
    2.221416e-20, -3.544313e-20, -3.209136e-20, -1.67685e-20, 2.16501e-20, 
    1.372077e-21, -3.637335e-21, 6.752182e-21, 1.411902e-20, 7.736633e-21, 
    -8.425669e-21, -2.293088e-20, 1.586827e-20, 1.949089e-20, -3.87802e-20, 
    2.4163e-20, -2.421645e-20, -9.774566e-21, 1.131772e-20, -2.69236e-20, 
    -1.933315e-20, 2.63534e-21, -1.499594e-21, -5.581959e-21, -2.84512e-20, 
    4.261024e-21, -2.19252e-20, 6.221502e-21, -1.365504e-20, 3.150979e-20, 
    -3.820002e-20, 2.978908e-20, -1.545887e-20, 2.846534e-21, 1.03918e-20, 
    -2.631856e-20, 1.207063e-20, 4.086984e-20, 3.034352e-20, -3.183889e-20, 
    -3.527857e-20, -1.962913e-20, 3.81664e-20, 1.457705e-20, 3.187784e-21, 
    -1.889152e-20, 2.996012e-20, -1.42225e-20, -7.050726e-21, 2.025627e-20, 
    -2.840002e-20, -1.858247e-20, 1.527764e-20, -1.787394e-20, -1.554312e-20, 
    9.577504e-21, 2.292212e-20, 1.319618e-20, 1.149555e-20, -1.677017e-20, 
    -1.575715e-20, -1.786772e-20, 1.549846e-20, 2.648451e-20, -1.396181e-20, 
    7.28767e-21, -4.400704e-20, -5.735702e-20, 1.108586e-20, -2.928837e-20, 
    -3.800694e-20, -2.357268e-20, -1.667689e-20, 2.395293e-21, -5.601576e-20, 
    2.610565e-20, -5.884765e-21, -2.344975e-21, 7.280263e-22, -2.256181e-21, 
    -5.810102e-21, -3.154442e-21, -9.215818e-23, 5.340222e-21, -2.572903e-22, 
    -4.008414e-20, -5.756398e-21, -1.427903e-20, -6.747096e-21, 4.073897e-20, 
    2.709804e-20, -1.052805e-20, -1.477862e-20, -3.244322e-21, 2.923832e-20, 
    -8.564477e-21, -8.719421e-21, 2.122346e-20, -3.403035e-20, 3.547932e-20, 
    2.182259e-20, -2.832933e-20, 1.793445e-20, 1.611846e-21, 4.704131e-20, 
    -1.8492e-20, 6.548605e-21, 3.99493e-20, -1.699891e-20, 1.634606e-20, 
    -1.084641e-20, -4.416424e-20, -4.946374e-20, 7.617615e-21, 9.988594e-21, 
    3.83751e-21, -4.110058e-20, -2.987079e-20, 2.564735e-20, 1.763957e-20, 
    -1.896304e-20, 2.962792e-20, 4.489225e-21, 4.647134e-20, -1.578478e-21, 
    -6.23362e-20, -2.590387e-21, 3.152421e-20, -2.210094e-21, 2.367248e-20, 
    3.716579e-20, 1.600652e-20, 8.922928e-22, -2.819136e-20, 1.299232e-20, 
    1.925709e-20, 1.111785e-20, -1.288121e-20, 1.259339e-20, 1.722367e-20, 
    4.919404e-20, -4.270706e-20, -2.411893e-20, -1.523523e-20, 7.969888e-21, 
    3.024286e-20, 1.584844e-20, -1.521034e-20, -9.578582e-22, 4.67453e-20, 
    -5.408093e-21, 2.735426e-21, 2.627078e-20, -2.19631e-20, -5.212427e-21, 
    3.654294e-21, -1.639557e-20, 5.299238e-21, -2.655777e-20, 3.088889e-20, 
    1.114694e-20, -7.42252e-21, 2.283022e-20, 3.732159e-20, 1.722452e-20, 
    2.441946e-20, -6.155893e-21, -1.473479e-20, -1.424679e-21, 2.566924e-21, 
    2.625126e-20, 1.133949e-20, 2.119038e-20, 1.272848e-21, 6.38549e-21, 
    3.549739e-20, -1.040366e-22, -2.423935e-20, 6.967622e-21, 2.327449e-21, 
    -9.904346e-21, 1.036999e-20, 1.665623e-20, 3.276455e-20, -6.655454e-20, 
    1.321342e-20, 6.87205e-21, 1.43404e-20, -3.126042e-20, 3.506315e-20, 
    -1.975158e-20, -3.39868e-20, -2.310363e-20, -2.109228e-20, 4.794916e-20, 
    -3.611037e-20, 2.372964e-21, -2.851735e-20, 1.758003e-21, -9.74631e-21, 
    -7.639389e-21, -2.86361e-20, 1.974224e-20, 5.509558e-21, -1.46432e-20, 
    -2.042844e-20, 2.470728e-20, 2.904859e-20, -3.489472e-21, 5.637101e-21, 
    -3.617766e-20, 3.380443e-20, 4.305994e-21, -2.073888e-20, 6.970446e-21, 
    2.502743e-21, -2.901779e-20, -2.168064e-20, -2.362751e-20, 1.761412e-20, 
    -2.570955e-20, 6.502031e-23, -3.026464e-20, -4.718098e-20, -1.716486e-20, 
    1.357362e-20, -5.199645e-20, 6.955113e-23, -4.869697e-20, -2.032211e-20, 
    -2.016549e-20, -1.011217e-20, -3.15519e-20, 2.443332e-20, 2.4476e-20, 
    -1.953445e-20, -2.487298e-20, 4.985108e-21 ;

 NBP =
  -6.359163e-08, -6.387121e-08, -6.381686e-08, -6.404235e-08, -6.391726e-08, 
    -6.406492e-08, -6.364831e-08, -6.388231e-08, -6.373293e-08, -6.36168e-08, 
    -6.447997e-08, -6.405241e-08, -6.492405e-08, -6.465138e-08, 
    -6.533632e-08, -6.488163e-08, -6.542801e-08, -6.53232e-08, -6.563863e-08, 
    -6.554826e-08, -6.595173e-08, -6.568033e-08, -6.616087e-08, 
    -6.588692e-08, -6.592978e-08, -6.567138e-08, -6.413845e-08, 
    -6.442674e-08, -6.412137e-08, -6.416248e-08, -6.414403e-08, 
    -6.391985e-08, -6.380688e-08, -6.357025e-08, -6.361321e-08, -6.3787e-08, 
    -6.418097e-08, -6.404723e-08, -6.438426e-08, -6.437665e-08, 
    -6.475187e-08, -6.458269e-08, -6.521333e-08, -6.503409e-08, 
    -6.555204e-08, -6.542178e-08, -6.554592e-08, -6.550827e-08, 
    -6.554641e-08, -6.535537e-08, -6.543722e-08, -6.526912e-08, 
    -6.461438e-08, -6.480681e-08, -6.423289e-08, -6.38878e-08, -6.365858e-08, 
    -6.349591e-08, -6.351891e-08, -6.356274e-08, -6.378801e-08, 
    -6.399981e-08, -6.416121e-08, -6.426918e-08, -6.437556e-08, 
    -6.469757e-08, -6.486799e-08, -6.524958e-08, -6.518071e-08, 
    -6.529738e-08, -6.540882e-08, -6.559594e-08, -6.556514e-08, 
    -6.564758e-08, -6.529429e-08, -6.552909e-08, -6.514148e-08, -6.52475e-08, 
    -6.44045e-08, -6.40833e-08, -6.394681e-08, -6.38273e-08, -6.353659e-08, 
    -6.373735e-08, -6.365821e-08, -6.384649e-08, -6.396612e-08, 
    -6.390695e-08, -6.427213e-08, -6.413016e-08, -6.487809e-08, 
    -6.455593e-08, -6.539582e-08, -6.519484e-08, -6.544399e-08, 
    -6.531685e-08, -6.55347e-08, -6.533864e-08, -6.567826e-08, -6.575221e-08, 
    -6.570168e-08, -6.58958e-08, -6.532778e-08, -6.554592e-08, -6.39053e-08, 
    -6.391495e-08, -6.39599e-08, -6.376228e-08, -6.375019e-08, -6.356908e-08, 
    -6.373023e-08, -6.379886e-08, -6.397305e-08, -6.40761e-08, -6.417405e-08, 
    -6.438941e-08, -6.462994e-08, -6.496626e-08, -6.520787e-08, 
    -6.536983e-08, -6.527052e-08, -6.53582e-08, -6.526018e-08, -6.521424e-08, 
    -6.572451e-08, -6.543799e-08, -6.586788e-08, -6.584409e-08, 
    -6.564954e-08, -6.584677e-08, -6.392172e-08, -6.386619e-08, 
    -6.367338e-08, -6.382427e-08, -6.354936e-08, -6.370324e-08, 
    -6.379173e-08, -6.413313e-08, -6.420814e-08, -6.427769e-08, 
    -6.441505e-08, -6.459135e-08, -6.49006e-08, -6.516968e-08, -6.54153e-08, 
    -6.539731e-08, -6.540364e-08, -6.545852e-08, -6.53226e-08, -6.548083e-08, 
    -6.550739e-08, -6.543795e-08, -6.58409e-08, -6.572579e-08, -6.584358e-08, 
    -6.576862e-08, -6.388424e-08, -6.397768e-08, -6.392719e-08, 
    -6.402214e-08, -6.395525e-08, -6.425269e-08, -6.434187e-08, 
    -6.475913e-08, -6.458788e-08, -6.486043e-08, -6.461556e-08, 
    -6.465896e-08, -6.486933e-08, -6.462879e-08, -6.515485e-08, 
    -6.479821e-08, -6.546065e-08, -6.510453e-08, -6.548296e-08, 
    -6.541424e-08, -6.552803e-08, -6.562993e-08, -6.575814e-08, -6.59947e-08, 
    -6.593991e-08, -6.613774e-08, -6.411698e-08, -6.423819e-08, 
    -6.422751e-08, -6.435434e-08, -6.444814e-08, -6.465145e-08, 
    -6.497752e-08, -6.485489e-08, -6.508e-08, -6.512519e-08, -6.47832e-08, 
    -6.499319e-08, -6.431929e-08, -6.442818e-08, -6.436335e-08, 
    -6.412655e-08, -6.488316e-08, -6.449487e-08, -6.521186e-08, 
    -6.500152e-08, -6.56154e-08, -6.531011e-08, -6.590976e-08, -6.616612e-08, 
    -6.640736e-08, -6.668932e-08, -6.430432e-08, -6.422197e-08, 
    -6.436942e-08, -6.457343e-08, -6.476271e-08, -6.501435e-08, 
    -6.504009e-08, -6.508724e-08, -6.520934e-08, -6.531201e-08, 
    -6.510215e-08, -6.533775e-08, -6.445345e-08, -6.491686e-08, 
    -6.419084e-08, -6.440948e-08, -6.456141e-08, -6.449476e-08, 
    -6.484088e-08, -6.492246e-08, -6.525397e-08, -6.50826e-08, -6.610285e-08, 
    -6.565147e-08, -6.690398e-08, -6.655396e-08, -6.41932e-08, -6.430404e-08, 
    -6.46898e-08, -6.450625e-08, -6.503114e-08, -6.516034e-08, -6.526538e-08, 
    -6.539964e-08, -6.541413e-08, -6.549368e-08, -6.536332e-08, 
    -6.548853e-08, -6.501489e-08, -6.522654e-08, -6.46457e-08, -6.478708e-08, 
    -6.472204e-08, -6.46507e-08, -6.487087e-08, -6.510545e-08, -6.511046e-08, 
    -6.518567e-08, -6.539766e-08, -6.503327e-08, -6.616113e-08, 
    -6.546461e-08, -6.44249e-08, -6.463841e-08, -6.466889e-08, -6.458619e-08, 
    -6.514739e-08, -6.494405e-08, -6.549174e-08, -6.534372e-08, 
    -6.558625e-08, -6.546573e-08, -6.5448e-08, -6.529321e-08, -6.519684e-08, 
    -6.495338e-08, -6.475528e-08, -6.459818e-08, -6.463471e-08, 
    -6.480727e-08, -6.51198e-08, -6.541545e-08, -6.535068e-08, -6.556781e-08, 
    -6.499309e-08, -6.523408e-08, -6.514095e-08, -6.538381e-08, 
    -6.485164e-08, -6.530484e-08, -6.47358e-08, -6.47857e-08, -6.494002e-08, 
    -6.525044e-08, -6.53191e-08, -6.539243e-08, -6.534718e-08, -6.512773e-08, 
    -6.509178e-08, -6.493626e-08, -6.489333e-08, -6.477483e-08, 
    -6.467673e-08, -6.476636e-08, -6.486049e-08, -6.512782e-08, 
    -6.536873e-08, -6.563138e-08, -6.569566e-08, -6.600256e-08, 
    -6.575274e-08, -6.616501e-08, -6.581453e-08, -6.642122e-08, 
    -6.533109e-08, -6.58042e-08, -6.494704e-08, -6.503938e-08, -6.520641e-08, 
    -6.558949e-08, -6.538266e-08, -6.562454e-08, -6.509037e-08, 
    -6.481324e-08, -6.474151e-08, -6.460773e-08, -6.474458e-08, 
    -6.473344e-08, -6.486439e-08, -6.482231e-08, -6.51367e-08, -6.496782e-08, 
    -6.544756e-08, -6.562262e-08, -6.611701e-08, -6.642009e-08, 
    -6.672858e-08, -6.686479e-08, -6.690624e-08, -6.692357e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.359163e-08, 6.387121e-08, 6.381686e-08, 6.404235e-08, 6.391726e-08, 
    6.406492e-08, 6.364831e-08, 6.388231e-08, 6.373293e-08, 6.36168e-08, 
    6.447997e-08, 6.405241e-08, 6.492405e-08, 6.465138e-08, 6.533632e-08, 
    6.488163e-08, 6.542801e-08, 6.53232e-08, 6.563863e-08, 6.554826e-08, 
    6.595173e-08, 6.568033e-08, 6.616087e-08, 6.588692e-08, 6.592978e-08, 
    6.567138e-08, 6.413845e-08, 6.442674e-08, 6.412137e-08, 6.416248e-08, 
    6.414403e-08, 6.391985e-08, 6.380688e-08, 6.357025e-08, 6.361321e-08, 
    6.3787e-08, 6.418097e-08, 6.404723e-08, 6.438426e-08, 6.437665e-08, 
    6.475187e-08, 6.458269e-08, 6.521333e-08, 6.503409e-08, 6.555204e-08, 
    6.542178e-08, 6.554592e-08, 6.550827e-08, 6.554641e-08, 6.535537e-08, 
    6.543722e-08, 6.526912e-08, 6.461438e-08, 6.480681e-08, 6.423289e-08, 
    6.38878e-08, 6.365858e-08, 6.349591e-08, 6.351891e-08, 6.356274e-08, 
    6.378801e-08, 6.399981e-08, 6.416121e-08, 6.426918e-08, 6.437556e-08, 
    6.469757e-08, 6.486799e-08, 6.524958e-08, 6.518071e-08, 6.529738e-08, 
    6.540882e-08, 6.559594e-08, 6.556514e-08, 6.564758e-08, 6.529429e-08, 
    6.552909e-08, 6.514148e-08, 6.52475e-08, 6.44045e-08, 6.40833e-08, 
    6.394681e-08, 6.38273e-08, 6.353659e-08, 6.373735e-08, 6.365821e-08, 
    6.384649e-08, 6.396612e-08, 6.390695e-08, 6.427213e-08, 6.413016e-08, 
    6.487809e-08, 6.455593e-08, 6.539582e-08, 6.519484e-08, 6.544399e-08, 
    6.531685e-08, 6.55347e-08, 6.533864e-08, 6.567826e-08, 6.575221e-08, 
    6.570168e-08, 6.58958e-08, 6.532778e-08, 6.554592e-08, 6.39053e-08, 
    6.391495e-08, 6.39599e-08, 6.376228e-08, 6.375019e-08, 6.356908e-08, 
    6.373023e-08, 6.379886e-08, 6.397305e-08, 6.40761e-08, 6.417405e-08, 
    6.438941e-08, 6.462994e-08, 6.496626e-08, 6.520787e-08, 6.536983e-08, 
    6.527052e-08, 6.53582e-08, 6.526018e-08, 6.521424e-08, 6.572451e-08, 
    6.543799e-08, 6.586788e-08, 6.584409e-08, 6.564954e-08, 6.584677e-08, 
    6.392172e-08, 6.386619e-08, 6.367338e-08, 6.382427e-08, 6.354936e-08, 
    6.370324e-08, 6.379173e-08, 6.413313e-08, 6.420814e-08, 6.427769e-08, 
    6.441505e-08, 6.459135e-08, 6.49006e-08, 6.516968e-08, 6.54153e-08, 
    6.539731e-08, 6.540364e-08, 6.545852e-08, 6.53226e-08, 6.548083e-08, 
    6.550739e-08, 6.543795e-08, 6.58409e-08, 6.572579e-08, 6.584358e-08, 
    6.576862e-08, 6.388424e-08, 6.397768e-08, 6.392719e-08, 6.402214e-08, 
    6.395525e-08, 6.425269e-08, 6.434187e-08, 6.475913e-08, 6.458788e-08, 
    6.486043e-08, 6.461556e-08, 6.465896e-08, 6.486933e-08, 6.462879e-08, 
    6.515485e-08, 6.479821e-08, 6.546065e-08, 6.510453e-08, 6.548296e-08, 
    6.541424e-08, 6.552803e-08, 6.562993e-08, 6.575814e-08, 6.59947e-08, 
    6.593991e-08, 6.613774e-08, 6.411698e-08, 6.423819e-08, 6.422751e-08, 
    6.435434e-08, 6.444814e-08, 6.465145e-08, 6.497752e-08, 6.485489e-08, 
    6.508e-08, 6.512519e-08, 6.47832e-08, 6.499319e-08, 6.431929e-08, 
    6.442818e-08, 6.436335e-08, 6.412655e-08, 6.488316e-08, 6.449487e-08, 
    6.521186e-08, 6.500152e-08, 6.56154e-08, 6.531011e-08, 6.590976e-08, 
    6.616612e-08, 6.640736e-08, 6.668932e-08, 6.430432e-08, 6.422197e-08, 
    6.436942e-08, 6.457343e-08, 6.476271e-08, 6.501435e-08, 6.504009e-08, 
    6.508724e-08, 6.520934e-08, 6.531201e-08, 6.510215e-08, 6.533775e-08, 
    6.445345e-08, 6.491686e-08, 6.419084e-08, 6.440948e-08, 6.456141e-08, 
    6.449476e-08, 6.484088e-08, 6.492246e-08, 6.525397e-08, 6.50826e-08, 
    6.610285e-08, 6.565147e-08, 6.690398e-08, 6.655396e-08, 6.41932e-08, 
    6.430404e-08, 6.46898e-08, 6.450625e-08, 6.503114e-08, 6.516034e-08, 
    6.526538e-08, 6.539964e-08, 6.541413e-08, 6.549368e-08, 6.536332e-08, 
    6.548853e-08, 6.501489e-08, 6.522654e-08, 6.46457e-08, 6.478708e-08, 
    6.472204e-08, 6.46507e-08, 6.487087e-08, 6.510545e-08, 6.511046e-08, 
    6.518567e-08, 6.539766e-08, 6.503327e-08, 6.616113e-08, 6.546461e-08, 
    6.44249e-08, 6.463841e-08, 6.466889e-08, 6.458619e-08, 6.514739e-08, 
    6.494405e-08, 6.549174e-08, 6.534372e-08, 6.558625e-08, 6.546573e-08, 
    6.5448e-08, 6.529321e-08, 6.519684e-08, 6.495338e-08, 6.475528e-08, 
    6.459818e-08, 6.463471e-08, 6.480727e-08, 6.51198e-08, 6.541545e-08, 
    6.535068e-08, 6.556781e-08, 6.499309e-08, 6.523408e-08, 6.514095e-08, 
    6.538381e-08, 6.485164e-08, 6.530484e-08, 6.47358e-08, 6.47857e-08, 
    6.494002e-08, 6.525044e-08, 6.53191e-08, 6.539243e-08, 6.534718e-08, 
    6.512773e-08, 6.509178e-08, 6.493626e-08, 6.489333e-08, 6.477483e-08, 
    6.467673e-08, 6.476636e-08, 6.486049e-08, 6.512782e-08, 6.536873e-08, 
    6.563138e-08, 6.569566e-08, 6.600256e-08, 6.575274e-08, 6.616501e-08, 
    6.581453e-08, 6.642122e-08, 6.533109e-08, 6.58042e-08, 6.494704e-08, 
    6.503938e-08, 6.520641e-08, 6.558949e-08, 6.538266e-08, 6.562454e-08, 
    6.509037e-08, 6.481324e-08, 6.474151e-08, 6.460773e-08, 6.474458e-08, 
    6.473344e-08, 6.486439e-08, 6.482231e-08, 6.51367e-08, 6.496782e-08, 
    6.544756e-08, 6.562262e-08, 6.611701e-08, 6.642009e-08, 6.672858e-08, 
    6.686479e-08, 6.690624e-08, 6.692357e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.359163e-08, -6.387121e-08, -6.381686e-08, -6.404235e-08, -6.391726e-08, 
    -6.406492e-08, -6.364831e-08, -6.388231e-08, -6.373293e-08, -6.36168e-08, 
    -6.447997e-08, -6.405241e-08, -6.492405e-08, -6.465138e-08, 
    -6.533632e-08, -6.488163e-08, -6.542801e-08, -6.53232e-08, -6.563863e-08, 
    -6.554826e-08, -6.595173e-08, -6.568033e-08, -6.616087e-08, 
    -6.588692e-08, -6.592978e-08, -6.567138e-08, -6.413845e-08, 
    -6.442674e-08, -6.412137e-08, -6.416248e-08, -6.414403e-08, 
    -6.391985e-08, -6.380688e-08, -6.357025e-08, -6.361321e-08, -6.3787e-08, 
    -6.418097e-08, -6.404723e-08, -6.438426e-08, -6.437665e-08, 
    -6.475187e-08, -6.458269e-08, -6.521333e-08, -6.503409e-08, 
    -6.555204e-08, -6.542178e-08, -6.554592e-08, -6.550827e-08, 
    -6.554641e-08, -6.535537e-08, -6.543722e-08, -6.526912e-08, 
    -6.461438e-08, -6.480681e-08, -6.423289e-08, -6.38878e-08, -6.365858e-08, 
    -6.349591e-08, -6.351891e-08, -6.356274e-08, -6.378801e-08, 
    -6.399981e-08, -6.416121e-08, -6.426918e-08, -6.437556e-08, 
    -6.469757e-08, -6.486799e-08, -6.524958e-08, -6.518071e-08, 
    -6.529738e-08, -6.540882e-08, -6.559594e-08, -6.556514e-08, 
    -6.564758e-08, -6.529429e-08, -6.552909e-08, -6.514148e-08, -6.52475e-08, 
    -6.44045e-08, -6.40833e-08, -6.394681e-08, -6.38273e-08, -6.353659e-08, 
    -6.373735e-08, -6.365821e-08, -6.384649e-08, -6.396612e-08, 
    -6.390695e-08, -6.427213e-08, -6.413016e-08, -6.487809e-08, 
    -6.455593e-08, -6.539582e-08, -6.519484e-08, -6.544399e-08, 
    -6.531685e-08, -6.55347e-08, -6.533864e-08, -6.567826e-08, -6.575221e-08, 
    -6.570168e-08, -6.58958e-08, -6.532778e-08, -6.554592e-08, -6.39053e-08, 
    -6.391495e-08, -6.39599e-08, -6.376228e-08, -6.375019e-08, -6.356908e-08, 
    -6.373023e-08, -6.379886e-08, -6.397305e-08, -6.40761e-08, -6.417405e-08, 
    -6.438941e-08, -6.462994e-08, -6.496626e-08, -6.520787e-08, 
    -6.536983e-08, -6.527052e-08, -6.53582e-08, -6.526018e-08, -6.521424e-08, 
    -6.572451e-08, -6.543799e-08, -6.586788e-08, -6.584409e-08, 
    -6.564954e-08, -6.584677e-08, -6.392172e-08, -6.386619e-08, 
    -6.367338e-08, -6.382427e-08, -6.354936e-08, -6.370324e-08, 
    -6.379173e-08, -6.413313e-08, -6.420814e-08, -6.427769e-08, 
    -6.441505e-08, -6.459135e-08, -6.49006e-08, -6.516968e-08, -6.54153e-08, 
    -6.539731e-08, -6.540364e-08, -6.545852e-08, -6.53226e-08, -6.548083e-08, 
    -6.550739e-08, -6.543795e-08, -6.58409e-08, -6.572579e-08, -6.584358e-08, 
    -6.576862e-08, -6.388424e-08, -6.397768e-08, -6.392719e-08, 
    -6.402214e-08, -6.395525e-08, -6.425269e-08, -6.434187e-08, 
    -6.475913e-08, -6.458788e-08, -6.486043e-08, -6.461556e-08, 
    -6.465896e-08, -6.486933e-08, -6.462879e-08, -6.515485e-08, 
    -6.479821e-08, -6.546065e-08, -6.510453e-08, -6.548296e-08, 
    -6.541424e-08, -6.552803e-08, -6.562993e-08, -6.575814e-08, -6.59947e-08, 
    -6.593991e-08, -6.613774e-08, -6.411698e-08, -6.423819e-08, 
    -6.422751e-08, -6.435434e-08, -6.444814e-08, -6.465145e-08, 
    -6.497752e-08, -6.485489e-08, -6.508e-08, -6.512519e-08, -6.47832e-08, 
    -6.499319e-08, -6.431929e-08, -6.442818e-08, -6.436335e-08, 
    -6.412655e-08, -6.488316e-08, -6.449487e-08, -6.521186e-08, 
    -6.500152e-08, -6.56154e-08, -6.531011e-08, -6.590976e-08, -6.616612e-08, 
    -6.640736e-08, -6.668932e-08, -6.430432e-08, -6.422197e-08, 
    -6.436942e-08, -6.457343e-08, -6.476271e-08, -6.501435e-08, 
    -6.504009e-08, -6.508724e-08, -6.520934e-08, -6.531201e-08, 
    -6.510215e-08, -6.533775e-08, -6.445345e-08, -6.491686e-08, 
    -6.419084e-08, -6.440948e-08, -6.456141e-08, -6.449476e-08, 
    -6.484088e-08, -6.492246e-08, -6.525397e-08, -6.50826e-08, -6.610285e-08, 
    -6.565147e-08, -6.690398e-08, -6.655396e-08, -6.41932e-08, -6.430404e-08, 
    -6.46898e-08, -6.450625e-08, -6.503114e-08, -6.516034e-08, -6.526538e-08, 
    -6.539964e-08, -6.541413e-08, -6.549368e-08, -6.536332e-08, 
    -6.548853e-08, -6.501489e-08, -6.522654e-08, -6.46457e-08, -6.478708e-08, 
    -6.472204e-08, -6.46507e-08, -6.487087e-08, -6.510545e-08, -6.511046e-08, 
    -6.518567e-08, -6.539766e-08, -6.503327e-08, -6.616113e-08, 
    -6.546461e-08, -6.44249e-08, -6.463841e-08, -6.466889e-08, -6.458619e-08, 
    -6.514739e-08, -6.494405e-08, -6.549174e-08, -6.534372e-08, 
    -6.558625e-08, -6.546573e-08, -6.5448e-08, -6.529321e-08, -6.519684e-08, 
    -6.495338e-08, -6.475528e-08, -6.459818e-08, -6.463471e-08, 
    -6.480727e-08, -6.51198e-08, -6.541545e-08, -6.535068e-08, -6.556781e-08, 
    -6.499309e-08, -6.523408e-08, -6.514095e-08, -6.538381e-08, 
    -6.485164e-08, -6.530484e-08, -6.47358e-08, -6.47857e-08, -6.494002e-08, 
    -6.525044e-08, -6.53191e-08, -6.539243e-08, -6.534718e-08, -6.512773e-08, 
    -6.509178e-08, -6.493626e-08, -6.489333e-08, -6.477483e-08, 
    -6.467673e-08, -6.476636e-08, -6.486049e-08, -6.512782e-08, 
    -6.536873e-08, -6.563138e-08, -6.569566e-08, -6.600256e-08, 
    -6.575274e-08, -6.616501e-08, -6.581453e-08, -6.642122e-08, 
    -6.533109e-08, -6.58042e-08, -6.494704e-08, -6.503938e-08, -6.520641e-08, 
    -6.558949e-08, -6.538266e-08, -6.562454e-08, -6.509037e-08, 
    -6.481324e-08, -6.474151e-08, -6.460773e-08, -6.474458e-08, 
    -6.473344e-08, -6.486439e-08, -6.482231e-08, -6.51367e-08, -6.496782e-08, 
    -6.544756e-08, -6.562262e-08, -6.611701e-08, -6.642009e-08, 
    -6.672858e-08, -6.686479e-08, -6.690624e-08, -6.692357e-08 ;

 NET_NMIN =
  8.958641e-09, 8.998025e-09, 8.990368e-09, 9.022133e-09, 9.004512e-09, 
    9.025312e-09, 8.966625e-09, 8.999589e-09, 8.978545e-09, 8.962186e-09, 
    9.08378e-09, 9.02355e-09, 9.146336e-09, 9.107925e-09, 9.204411e-09, 
    9.14036e-09, 9.217326e-09, 9.202562e-09, 9.246996e-09, 9.234267e-09, 
    9.291101e-09, 9.252871e-09, 9.320561e-09, 9.281971e-09, 9.288009e-09, 
    9.25161e-09, 9.03567e-09, 9.076282e-09, 9.033264e-09, 9.039055e-09, 
    9.036456e-09, 9.004876e-09, 8.988962e-09, 8.95563e-09, 8.961681e-09, 
    8.986163e-09, 9.041659e-09, 9.02282e-09, 9.070297e-09, 9.069225e-09, 
    9.122081e-09, 9.098249e-09, 9.187086e-09, 9.161837e-09, 9.234798e-09, 
    9.216449e-09, 9.233936e-09, 9.228634e-09, 9.234006e-09, 9.207095e-09, 
    9.218625e-09, 9.194944e-09, 9.102713e-09, 9.12982e-09, 9.048974e-09, 
    9.000362e-09, 8.968071e-09, 8.945158e-09, 8.948397e-09, 8.954572e-09, 
    8.986306e-09, 9.016141e-09, 9.038876e-09, 9.054085e-09, 9.069071e-09, 
    9.114433e-09, 9.138438e-09, 9.192192e-09, 9.18249e-09, 9.198925e-09, 
    9.214624e-09, 9.240982e-09, 9.236643e-09, 9.248257e-09, 9.19849e-09, 
    9.231566e-09, 9.176964e-09, 9.191899e-09, 9.073149e-09, 9.027902e-09, 
    9.008674e-09, 8.991839e-09, 8.950887e-09, 8.979169e-09, 8.96802e-09, 
    8.994542e-09, 9.011395e-09, 9.00306e-09, 9.054501e-09, 9.034503e-09, 
    9.139861e-09, 9.094481e-09, 9.212792e-09, 9.184482e-09, 9.219578e-09, 
    9.201669e-09, 9.232356e-09, 9.204738e-09, 9.252578e-09, 9.262997e-09, 
    9.255877e-09, 9.283222e-09, 9.203207e-09, 9.233936e-09, 9.002826e-09, 
    9.004186e-09, 9.010519e-09, 8.98268e-09, 8.980977e-09, 8.955464e-09, 
    8.978165e-09, 8.987833e-09, 9.012371e-09, 9.026887e-09, 9.040686e-09, 
    9.071023e-09, 9.104904e-09, 9.152282e-09, 9.186317e-09, 9.209131e-09, 
    9.195142e-09, 9.207493e-09, 9.193686e-09, 9.187214e-09, 9.259093e-09, 
    9.218732e-09, 9.279289e-09, 9.275938e-09, 9.248533e-09, 9.276316e-09, 
    9.005141e-09, 8.997318e-09, 8.970157e-09, 8.991412e-09, 8.952686e-09, 
    8.974363e-09, 8.986828e-09, 9.034921e-09, 9.045487e-09, 9.055285e-09, 
    9.074635e-09, 9.09947e-09, 9.143033e-09, 9.180937e-09, 9.215537e-09, 
    9.213002e-09, 9.213895e-09, 9.221624e-09, 9.202477e-09, 9.224768e-09, 
    9.228509e-09, 9.218727e-09, 9.27549e-09, 9.259273e-09, 9.275867e-09, 
    9.265309e-09, 8.99986e-09, 9.013023e-09, 9.005911e-09, 9.019286e-09, 
    9.009863e-09, 9.051763e-09, 9.064325e-09, 9.123105e-09, 9.09898e-09, 
    9.137374e-09, 9.10288e-09, 9.108993e-09, 9.138628e-09, 9.104744e-09, 
    9.178848e-09, 9.12861e-09, 9.221925e-09, 9.171759e-09, 9.225069e-09, 
    9.215388e-09, 9.231416e-09, 9.245771e-09, 9.263831e-09, 9.297153e-09, 
    9.289437e-09, 9.317304e-09, 9.032646e-09, 9.04972e-09, 9.048216e-09, 
    9.066082e-09, 9.079296e-09, 9.107935e-09, 9.153868e-09, 9.136595e-09, 
    9.168304e-09, 9.17467e-09, 9.126495e-09, 9.156075e-09, 9.061146e-09, 
    9.076484e-09, 9.06735e-09, 9.033993e-09, 9.140576e-09, 9.085879e-09, 
    9.186879e-09, 9.157248e-09, 9.243725e-09, 9.200719e-09, 9.28519e-09, 
    9.321301e-09, 9.355284e-09, 9.395001e-09, 9.059037e-09, 9.047436e-09, 
    9.068207e-09, 9.096946e-09, 9.123609e-09, 9.159057e-09, 9.162682e-09, 
    9.169323e-09, 9.186524e-09, 9.200987e-09, 9.171425e-09, 9.204612e-09, 
    9.080042e-09, 9.145324e-09, 9.043051e-09, 9.073849e-09, 9.095252e-09, 
    9.085862e-09, 9.13462e-09, 9.146112e-09, 9.192811e-09, 9.16867e-09, 
    9.312389e-09, 9.248804e-09, 9.42524e-09, 9.375935e-09, 9.043383e-09, 
    9.058996e-09, 9.113338e-09, 9.087482e-09, 9.161422e-09, 9.179622e-09, 
    9.194417e-09, 9.213331e-09, 9.215372e-09, 9.226578e-09, 9.208215e-09, 
    9.225852e-09, 9.159131e-09, 9.188947e-09, 9.107126e-09, 9.127041e-09, 
    9.117879e-09, 9.107829e-09, 9.138845e-09, 9.171889e-09, 9.172594e-09, 
    9.18319e-09, 9.213051e-09, 9.161721e-09, 9.320599e-09, 9.222483e-09, 
    9.076023e-09, 9.106098e-09, 9.110392e-09, 9.098742e-09, 9.177797e-09, 
    9.149153e-09, 9.226304e-09, 9.205453e-09, 9.239617e-09, 9.22264e-09, 
    9.220143e-09, 9.198338e-09, 9.184763e-09, 9.150467e-09, 9.122561e-09, 
    9.100432e-09, 9.105577e-09, 9.129886e-09, 9.173911e-09, 9.215557e-09, 
    9.206435e-09, 9.237021e-09, 9.156061e-09, 9.19001e-09, 9.176889e-09, 
    9.2111e-09, 9.136135e-09, 9.199977e-09, 9.119818e-09, 9.126846e-09, 
    9.148585e-09, 9.192314e-09, 9.201986e-09, 9.212315e-09, 9.205941e-09, 
    9.175028e-09, 9.169963e-09, 9.148056e-09, 9.142008e-09, 9.125316e-09, 
    9.111496e-09, 9.124123e-09, 9.137383e-09, 9.17504e-09, 9.208977e-09, 
    9.245976e-09, 9.25503e-09, 9.298263e-09, 9.263071e-09, 9.321146e-09, 
    9.271774e-09, 9.357237e-09, 9.203674e-09, 9.27032e-09, 9.149574e-09, 
    9.162582e-09, 9.186111e-09, 9.240074e-09, 9.21094e-09, 9.245011e-09, 
    9.169765e-09, 9.130726e-09, 9.120622e-09, 9.101777e-09, 9.121054e-09, 
    9.119486e-09, 9.137931e-09, 9.132004e-09, 9.176291e-09, 9.152502e-09, 
    9.220081e-09, 9.244742e-09, 9.314384e-09, 9.357077e-09, 9.400534e-09, 
    9.419719e-09, 9.425558e-09, 9.428e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14 ;

 O_SCALAR =
  0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8 ;

 PCH4 =
  0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993 ;

 PCO2 =
  29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  4.726044e-14, 4.73878e-14, 4.736306e-14, 4.746568e-14, 4.740878e-14, 
    4.747595e-14, 4.728629e-14, 4.739284e-14, 4.732484e-14, 4.727194e-14, 
    4.766455e-14, 4.747026e-14, 4.786618e-14, 4.774249e-14, 4.805298e-14, 
    4.784692e-14, 4.809449e-14, 4.804707e-14, 4.818983e-14, 4.814895e-14, 
    4.833127e-14, 4.820869e-14, 4.842573e-14, 4.830203e-14, 4.832137e-14, 
    4.820464e-14, 4.750942e-14, 4.764037e-14, 4.750165e-14, 4.752034e-14, 
    4.751196e-14, 4.740994e-14, 4.735847e-14, 4.725073e-14, 4.72703e-14, 
    4.734945e-14, 4.752874e-14, 4.746793e-14, 4.76212e-14, 4.761774e-14, 
    4.77881e-14, 4.771132e-14, 4.799731e-14, 4.791613e-14, 4.815066e-14, 
    4.809171e-14, 4.814788e-14, 4.813086e-14, 4.814811e-14, 4.806164e-14, 
    4.809869e-14, 4.802259e-14, 4.77257e-14, 4.781302e-14, 4.755236e-14, 
    4.73953e-14, 4.729096e-14, 4.721684e-14, 4.722731e-14, 4.724729e-14, 
    4.734991e-14, 4.744636e-14, 4.751979e-14, 4.756888e-14, 4.761724e-14, 
    4.776339e-14, 4.784075e-14, 4.801371e-14, 4.798254e-14, 4.803536e-14, 
    4.808584e-14, 4.817051e-14, 4.815658e-14, 4.819386e-14, 4.803399e-14, 
    4.814025e-14, 4.796478e-14, 4.80128e-14, 4.763025e-14, 4.748435e-14, 
    4.742217e-14, 4.736781e-14, 4.723537e-14, 4.732684e-14, 4.729079e-14, 
    4.737657e-14, 4.743102e-14, 4.74041e-14, 4.757022e-14, 4.750566e-14, 
    4.784534e-14, 4.769915e-14, 4.807996e-14, 4.798894e-14, 4.810177e-14, 
    4.804421e-14, 4.81428e-14, 4.805408e-14, 4.820774e-14, 4.824116e-14, 
    4.821832e-14, 4.830607e-14, 4.804915e-14, 4.814787e-14, 4.740334e-14, 
    4.740773e-14, 4.74282e-14, 4.733819e-14, 4.733269e-14, 4.725018e-14, 
    4.732361e-14, 4.735486e-14, 4.743419e-14, 4.748107e-14, 4.752562e-14, 
    4.762352e-14, 4.773274e-14, 4.788534e-14, 4.799484e-14, 4.80682e-14, 
    4.802323e-14, 4.806293e-14, 4.801855e-14, 4.799774e-14, 4.822863e-14, 
    4.809903e-14, 4.829345e-14, 4.828271e-14, 4.819474e-14, 4.828392e-14, 
    4.741081e-14, 4.738554e-14, 4.729771e-14, 4.736645e-14, 4.72412e-14, 
    4.731131e-14, 4.735159e-14, 4.750698e-14, 4.754113e-14, 4.757274e-14, 
    4.763518e-14, 4.771525e-14, 4.785557e-14, 4.797753e-14, 4.808878e-14, 
    4.808064e-14, 4.808351e-14, 4.810833e-14, 4.804681e-14, 4.811843e-14, 
    4.813044e-14, 4.809903e-14, 4.828127e-14, 4.822924e-14, 4.828248e-14, 
    4.824861e-14, 4.739376e-14, 4.743628e-14, 4.741331e-14, 4.745651e-14, 
    4.742606e-14, 4.756134e-14, 4.760187e-14, 4.779137e-14, 4.771367e-14, 
    4.783734e-14, 4.772625e-14, 4.774593e-14, 4.784132e-14, 4.773226e-14, 
    4.797078e-14, 4.780908e-14, 4.81093e-14, 4.794797e-14, 4.81194e-14, 
    4.80883e-14, 4.81398e-14, 4.818588e-14, 4.824386e-14, 4.835071e-14, 
    4.832598e-14, 4.841531e-14, 4.749967e-14, 4.755476e-14, 4.754994e-14, 
    4.760759e-14, 4.76502e-14, 4.774254e-14, 4.789046e-14, 4.783487e-14, 
    4.793694e-14, 4.795738e-14, 4.780235e-14, 4.789755e-14, 4.759164e-14, 
    4.76411e-14, 4.761167e-14, 4.7504e-14, 4.784765e-14, 4.76714e-14, 
    4.799665e-14, 4.790135e-14, 4.817931e-14, 4.804112e-14, 4.831236e-14, 
    4.842806e-14, 4.853695e-14, 4.866394e-14, 4.758485e-14, 4.754742e-14, 
    4.761445e-14, 4.770708e-14, 4.779303e-14, 4.790716e-14, 4.791885e-14, 
    4.794021e-14, 4.799552e-14, 4.804202e-14, 4.794694e-14, 4.805368e-14, 
    4.765251e-14, 4.786295e-14, 4.753325e-14, 4.763259e-14, 4.770163e-14, 
    4.767138e-14, 4.782852e-14, 4.786551e-14, 4.801571e-14, 4.793812e-14, 
    4.839949e-14, 4.819558e-14, 4.876061e-14, 4.860298e-14, 4.753434e-14, 
    4.758473e-14, 4.775992e-14, 4.76766e-14, 4.791479e-14, 4.797331e-14, 
    4.80209e-14, 4.808167e-14, 4.808825e-14, 4.812424e-14, 4.806525e-14, 
    4.812192e-14, 4.79074e-14, 4.800331e-14, 4.773994e-14, 4.780409e-14, 
    4.777459e-14, 4.774221e-14, 4.784212e-14, 4.79484e-14, 4.795071e-14, 
    4.798477e-14, 4.808063e-14, 4.791576e-14, 4.842571e-14, 4.811095e-14, 
    4.763966e-14, 4.773657e-14, 4.775045e-14, 4.771292e-14, 4.796744e-14, 
    4.787529e-14, 4.812337e-14, 4.805638e-14, 4.816614e-14, 4.81116e-14, 
    4.810358e-14, 4.803351e-14, 4.798985e-14, 4.787951e-14, 4.778965e-14, 
    4.771837e-14, 4.773495e-14, 4.781324e-14, 4.795491e-14, 4.808883e-14, 
    4.80595e-14, 4.81578e-14, 4.789753e-14, 4.80067e-14, 4.79645e-14, 
    4.807452e-14, 4.783338e-14, 4.803863e-14, 4.778084e-14, 4.780347e-14, 
    4.787346e-14, 4.801408e-14, 4.804523e-14, 4.807841e-14, 4.805795e-14, 
    4.795851e-14, 4.794226e-14, 4.787177e-14, 4.785228e-14, 4.779855e-14, 
    4.775402e-14, 4.779469e-14, 4.783738e-14, 4.795857e-14, 4.806768e-14, 
    4.818653e-14, 4.821562e-14, 4.835419e-14, 4.824134e-14, 4.842745e-14, 
    4.826916e-14, 4.854308e-14, 4.805057e-14, 4.826458e-14, 4.787666e-14, 
    4.791852e-14, 4.799414e-14, 4.816754e-14, 4.8074e-14, 4.81834e-14, 
    4.794162e-14, 4.781592e-14, 4.778343e-14, 4.77227e-14, 4.778481e-14, 
    4.777977e-14, 4.783918e-14, 4.782009e-14, 4.796259e-14, 4.788608e-14, 
    4.810336e-14, 4.818255e-14, 4.840594e-14, 4.854264e-14, 4.868169e-14, 
    4.8743e-14, 4.876165e-14, 4.876945e-14 ;

 POT_F_DENIT =
  4.592699e-13, 4.603734e-13, 4.601579e-13, 4.610479e-13, 4.605535e-13, 
    4.611356e-13, 4.594913e-13, 4.604144e-13, 4.598244e-13, 4.593652e-13, 
    4.627707e-13, 4.610841e-13, 4.64519e-13, 4.63444e-13, 4.661405e-13, 
    4.64351e-13, 4.665006e-13, 4.660873e-13, 4.673277e-13, 4.669717e-13, 
    4.685577e-13, 4.674905e-13, 4.693781e-13, 4.683019e-13, 4.684699e-13, 
    4.674532e-13, 4.614263e-13, 4.625641e-13, 4.613581e-13, 4.615204e-13, 
    4.61447e-13, 4.60562e-13, 4.601164e-13, 4.591812e-13, 4.593503e-13, 
    4.600366e-13, 4.615902e-13, 4.610619e-13, 4.623902e-13, 4.623603e-13, 
    4.638381e-13, 4.631716e-13, 4.656545e-13, 4.649483e-13, 4.66986e-13, 
    4.664731e-13, 4.669612e-13, 4.668124e-13, 4.669619e-13, 4.662106e-13, 
    4.665316e-13, 4.658703e-13, 4.633017e-13, 4.640592e-13, 4.617972e-13, 
    4.604358e-13, 4.5953e-13, 4.588878e-13, 4.589776e-13, 4.591509e-13, 
    4.600397e-13, 4.608744e-13, 4.615109e-13, 4.619359e-13, 4.623547e-13, 
    4.636247e-13, 4.642951e-13, 4.657964e-13, 4.655249e-13, 4.659836e-13, 
    4.664216e-13, 4.671569e-13, 4.670356e-13, 4.673592e-13, 4.659689e-13, 
    4.668929e-13, 4.653666e-13, 4.65784e-13, 4.624745e-13, 4.612061e-13, 
    4.60668e-13, 4.601954e-13, 4.590472e-13, 4.5984e-13, 4.59527e-13, 
    4.602692e-13, 4.607411e-13, 4.605069e-13, 4.619471e-13, 4.613866e-13, 
    4.643341e-13, 4.630649e-13, 4.663711e-13, 4.655796e-13, 4.665592e-13, 
    4.660592e-13, 4.669153e-13, 4.661441e-13, 4.674788e-13, 4.677698e-13, 
    4.675701e-13, 4.683331e-13, 4.660986e-13, 4.669569e-13, 4.60503e-13, 
    4.605412e-13, 4.607179e-13, 4.599377e-13, 4.598897e-13, 4.59174e-13, 
    4.598096e-13, 4.600806e-13, 4.607672e-13, 4.611731e-13, 4.615589e-13, 
    4.624081e-13, 4.633557e-13, 4.646797e-13, 4.656304e-13, 4.662669e-13, 
    4.658759e-13, 4.662203e-13, 4.658345e-13, 4.656529e-13, 4.676597e-13, 
    4.66533e-13, 4.682221e-13, 4.681287e-13, 4.673635e-13, 4.68138e-13, 
    4.60567e-13, 4.603471e-13, 4.595862e-13, 4.601809e-13, 4.590952e-13, 
    4.59703e-13, 4.600518e-13, 4.61398e-13, 4.616929e-13, 4.619674e-13, 
    4.625083e-13, 4.632024e-13, 4.644207e-13, 4.654792e-13, 4.664453e-13, 
    4.663738e-13, 4.663986e-13, 4.666138e-13, 4.660789e-13, 4.667007e-13, 
    4.668047e-13, 4.665315e-13, 4.681149e-13, 4.676625e-13, 4.681249e-13, 
    4.678296e-13, 4.604179e-13, 4.60786e-13, 4.605862e-13, 4.60961e-13, 
    4.606962e-13, 4.618696e-13, 4.622208e-13, 4.638644e-13, 4.631888e-13, 
    4.642627e-13, 4.632969e-13, 4.634681e-13, 4.642969e-13, 4.633478e-13, 
    4.654197e-13, 4.640151e-13, 4.666217e-13, 4.652204e-13, 4.667086e-13, 
    4.664375e-13, 4.668845e-13, 4.672854e-13, 4.677884e-13, 4.687184e-13, 
    4.685021e-13, 4.692792e-13, 4.61335e-13, 4.618124e-13, 4.617699e-13, 
    4.622693e-13, 4.626386e-13, 4.634398e-13, 4.647236e-13, 4.6424e-13, 
    4.651257e-13, 4.653037e-13, 4.639561e-13, 4.647834e-13, 4.621277e-13, 
    4.625565e-13, 4.623004e-13, 4.613661e-13, 4.64348e-13, 4.628177e-13, 
    4.656409e-13, 4.648122e-13, 4.672271e-13, 4.660266e-13, 4.683833e-13, 
    4.69391e-13, 4.703369e-13, 4.714431e-13, 4.620726e-13, 4.617471e-13, 
    4.623279e-13, 4.631325e-13, 4.63877e-13, 4.648681e-13, 4.649687e-13, 
    4.651537e-13, 4.656336e-13, 4.660377e-13, 4.652116e-13, 4.661377e-13, 
    4.626562e-13, 4.644805e-13, 4.616188e-13, 4.624812e-13, 4.630788e-13, 
    4.628161e-13, 4.64179e-13, 4.644997e-13, 4.658043e-13, 4.651297e-13, 
    4.691413e-13, 4.673672e-13, 4.722836e-13, 4.709111e-13, 4.616332e-13, 
    4.620695e-13, 4.635896e-13, 4.628663e-13, 4.649328e-13, 4.654415e-13, 
    4.658538e-13, 4.663824e-13, 4.664382e-13, 4.667513e-13, 4.662375e-13, 
    4.667301e-13, 4.648655e-13, 4.656986e-13, 4.634107e-13, 4.639672e-13, 
    4.637106e-13, 4.634289e-13, 4.642956e-13, 4.652197e-13, 4.652385e-13, 
    4.655341e-13, 4.663692e-13, 4.649331e-13, 4.693692e-13, 4.666309e-13, 
    4.625455e-13, 4.633867e-13, 4.635059e-13, 4.6318e-13, 4.653893e-13, 
    4.645889e-13, 4.667436e-13, 4.661606e-13, 4.67114e-13, 4.666401e-13, 
    4.665694e-13, 4.659605e-13, 4.655804e-13, 4.646223e-13, 4.638411e-13, 
    4.632221e-13, 4.63365e-13, 4.640451e-13, 4.652749e-13, 4.664382e-13, 
    4.661829e-13, 4.67036e-13, 4.647741e-13, 4.657229e-13, 4.653555e-13, 
    4.66311e-13, 4.642254e-13, 4.660107e-13, 4.637686e-13, 4.639644e-13, 
    4.645717e-13, 4.657942e-13, 4.660629e-13, 4.663517e-13, 4.661725e-13, 
    4.653093e-13, 4.65167e-13, 4.64554e-13, 4.643845e-13, 4.639177e-13, 
    4.635303e-13, 4.638835e-13, 4.642535e-13, 4.65306e-13, 4.662536e-13, 
    4.672858e-13, 4.675382e-13, 4.687446e-13, 4.677624e-13, 4.693824e-13, 
    4.680053e-13, 4.70387e-13, 4.661122e-13, 4.679729e-13, 4.645993e-13, 
    4.649622e-13, 4.656199e-13, 4.671263e-13, 4.663118e-13, 4.672636e-13, 
    4.651612e-13, 4.640695e-13, 4.637861e-13, 4.632592e-13, 4.637973e-13, 
    4.637535e-13, 4.642687e-13, 4.641023e-13, 4.653397e-13, 4.646748e-13, 
    4.66562e-13, 4.672507e-13, 4.69193e-13, 4.703825e-13, 4.715922e-13, 
    4.721256e-13, 4.72288e-13, 4.723554e-13 ;

 POT_F_NIT =
  4.024307e-11, 4.05898e-11, 4.052226e-11, 4.080281e-11, 4.064705e-11, 
    4.083092e-11, 4.031322e-11, 4.060357e-11, 4.041808e-11, 4.027418e-11, 
    4.135007e-11, 4.081531e-11, 4.19093e-11, 4.156545e-11, 4.243196e-11, 
    4.18557e-11, 4.254865e-11, 4.241526e-11, 4.281734e-11, 4.270194e-11, 
    4.321838e-11, 4.287063e-11, 4.348734e-11, 4.313519e-11, 4.319018e-11, 
    4.285917e-11, 4.092265e-11, 4.128333e-11, 4.090133e-11, 4.095265e-11, 
    4.092961e-11, 4.065025e-11, 4.050985e-11, 4.021659e-11, 4.026974e-11, 
    4.048516e-11, 4.09757e-11, 4.080883e-11, 4.123003e-11, 4.122049e-11, 
    4.169198e-11, 4.147905e-11, 4.227567e-11, 4.204844e-11, 4.270675e-11, 
    4.254069e-11, 4.269893e-11, 4.265091e-11, 4.269955e-11, 4.245615e-11, 
    4.256033e-11, 4.234648e-11, 4.151894e-11, 4.17613e-11, 4.104061e-11, 
    4.06104e-11, 4.032591e-11, 4.012468e-11, 4.015309e-11, 4.020729e-11, 
    4.048642e-11, 4.074975e-11, 4.095102e-11, 4.108594e-11, 4.12191e-11, 
    4.162358e-11, 4.183846e-11, 4.232168e-11, 4.223425e-11, 4.23824e-11, 
    4.252418e-11, 4.276277e-11, 4.272345e-11, 4.282874e-11, 4.237846e-11, 
    4.267744e-11, 4.218445e-11, 4.2319e-11, 4.125543e-11, 4.085383e-11, 
    4.068378e-11, 4.05352e-11, 4.017494e-11, 4.042355e-11, 4.032545e-11, 
    4.055901e-11, 4.070779e-11, 4.063417e-11, 4.108963e-11, 4.091224e-11, 
    4.18512e-11, 4.144541e-11, 4.250764e-11, 4.225217e-11, 4.256897e-11, 
    4.240716e-11, 4.26846e-11, 4.243486e-11, 4.286795e-11, 4.296256e-11, 
    4.289788e-11, 4.314655e-11, 4.242101e-11, 4.269889e-11, 4.063213e-11, 
    4.064414e-11, 4.070007e-11, 4.045447e-11, 4.043947e-11, 4.021511e-11, 
    4.04147e-11, 4.049985e-11, 4.071641e-11, 4.08448e-11, 4.096703e-11, 
    4.123646e-11, 4.153843e-11, 4.19626e-11, 4.226871e-11, 4.247454e-11, 
    4.234825e-11, 4.245973e-11, 4.233511e-11, 4.227677e-11, 4.292709e-11, 
    4.256129e-11, 4.311072e-11, 4.308023e-11, 4.283121e-11, 4.308365e-11, 
    4.065255e-11, 4.05835e-11, 4.034424e-11, 4.053141e-11, 4.01907e-11, 
    4.038123e-11, 4.049099e-11, 4.091595e-11, 4.100961e-11, 4.109657e-11, 
    4.126859e-11, 4.14899e-11, 4.187962e-11, 4.222023e-11, 4.253242e-11, 
    4.25095e-11, 4.251756e-11, 4.258745e-11, 4.241443e-11, 4.261588e-11, 
    4.264973e-11, 4.256123e-11, 4.307613e-11, 4.29287e-11, 4.307956e-11, 
    4.298352e-11, 4.060593e-11, 4.072218e-11, 4.065933e-11, 4.077754e-11, 
    4.069424e-11, 4.106531e-11, 4.117689e-11, 4.170111e-11, 4.148554e-11, 
    4.182888e-11, 4.152034e-11, 4.157492e-11, 4.184011e-11, 4.153696e-11, 
    4.220141e-11, 4.175035e-11, 4.259016e-11, 4.21376e-11, 4.26186e-11, 
    4.253103e-11, 4.267604e-11, 4.280614e-11, 4.297009e-11, 4.327349e-11, 
    4.320312e-11, 4.345747e-11, 4.08958e-11, 4.104717e-11, 4.103382e-11, 
    4.119251e-11, 4.131008e-11, 4.156549e-11, 4.197684e-11, 4.18219e-11, 
    4.210655e-11, 4.216381e-11, 4.173143e-11, 4.199664e-11, 4.114859e-11, 
    4.1285e-11, 4.120375e-11, 4.090767e-11, 4.185755e-11, 4.136866e-11, 
    4.227372e-11, 4.200714e-11, 4.278757e-11, 4.239853e-11, 4.316442e-11, 
    4.349402e-11, 4.380537e-11, 4.417072e-11, 4.11299e-11, 4.102689e-11, 
    4.12114e-11, 4.146739e-11, 4.170561e-11, 4.202343e-11, 4.205601e-11, 
    4.211571e-11, 4.227055e-11, 4.240098e-11, 4.213459e-11, 4.243369e-11, 
    4.131668e-11, 4.190012e-11, 4.098794e-11, 4.126154e-11, 4.145221e-11, 
    4.13685e-11, 4.180415e-11, 4.190717e-11, 4.232717e-11, 4.210978e-11, 
    4.341254e-11, 4.283363e-11, 4.444993e-11, 4.399513e-11, 4.099094e-11, 
    4.112952e-11, 4.161375e-11, 4.138299e-11, 4.204468e-11, 4.220839e-11, 
    4.23417e-11, 4.251246e-11, 4.25309e-11, 4.263226e-11, 4.246622e-11, 
    4.262568e-11, 4.202406e-11, 4.229236e-11, 4.15582e-11, 4.173627e-11, 
    4.165429e-11, 4.156447e-11, 4.1842e-11, 4.213873e-11, 4.214506e-11, 
    4.224044e-11, 4.250986e-11, 4.204729e-11, 4.348756e-11, 4.259513e-11, 
    4.128092e-11, 4.154906e-11, 4.158742e-11, 4.148339e-11, 4.219195e-11, 
    4.193449e-11, 4.262979e-11, 4.244128e-11, 4.275035e-11, 4.259662e-11, 
    4.257402e-11, 4.237705e-11, 4.225464e-11, 4.194625e-11, 4.169617e-11, 
    4.149842e-11, 4.154434e-11, 4.176173e-11, 4.21569e-11, 4.253252e-11, 
    4.245009e-11, 4.272676e-11, 4.199643e-11, 4.230188e-11, 4.218368e-11, 
    4.249221e-11, 4.181777e-11, 4.239186e-11, 4.167167e-11, 4.173455e-11, 
    4.192938e-11, 4.232271e-11, 4.240996e-11, 4.250326e-11, 4.244567e-11, 
    4.216699e-11, 4.212141e-11, 4.192461e-11, 4.187035e-11, 4.172082e-11, 
    4.159722e-11, 4.171013e-11, 4.182888e-11, 4.216706e-11, 4.247305e-11, 
    4.280794e-11, 4.28901e-11, 4.328354e-11, 4.296314e-11, 4.349254e-11, 
    4.304225e-11, 4.382324e-11, 4.242522e-11, 4.302911e-11, 4.193825e-11, 
    4.205507e-11, 4.22668e-11, 4.275448e-11, 4.249082e-11, 4.279924e-11, 
    4.211963e-11, 4.176925e-11, 4.167882e-11, 4.151042e-11, 4.168267e-11, 
    4.166864e-11, 4.183379e-11, 4.178068e-11, 4.217831e-11, 4.196447e-11, 
    4.257339e-11, 4.279674e-11, 4.343073e-11, 4.382178e-11, 4.422169e-11, 
    4.439884e-11, 4.445283e-11, 4.447541e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.001212904, 0.001212831, 0.001212845, 0.001212786, 0.001212818, 
    0.00121278, 0.001212888, 0.001212828, 0.001212866, 0.001212896, 
    0.001212676, 0.001212784, 0.001212558, 0.001212628, 0.001212449, 
    0.00121257, 0.001212425, 0.001212451, 0.001212369, 0.001212393, 
    0.00121229, 0.001212358, 0.001212235, 0.001212306, 0.001212295, 
    0.001212361, 0.001212761, 0.00121269, 0.001212765, 0.001212755, 
    0.001212759, 0.001212818, 0.001212848, 0.001212908, 0.001212897, 
    0.001212853, 0.00121275, 0.001212784, 0.001212696, 0.001212698, 
    0.001212601, 0.001212645, 0.00121248, 0.001212528, 0.001212392, 
    0.001212426, 0.001212393, 0.001212403, 0.001212393, 0.001212443, 
    0.001212422, 0.001212465, 0.001212637, 0.001212587, 0.001212736, 
    0.001212828, 0.001212886, 0.001212928, 0.001212922, 0.001212911, 
    0.001212853, 0.001212796, 0.001212754, 0.001212726, 0.001212698, 
    0.001212618, 0.001212572, 0.001212471, 0.001212488, 0.001212459, 
    0.001212429, 0.001212381, 0.001212388, 0.001212367, 0.001212458, 
    0.001212398, 0.001212498, 0.001212471, 0.001212696, 0.001212775, 
    0.001212812, 0.001212842, 0.001212918, 0.001212866, 0.001212886, 
    0.001212836, 0.001212805, 0.00121282, 0.001212725, 0.001212763, 
    0.00121257, 0.001212653, 0.001212432, 0.001212484, 0.00121242, 
    0.001212452, 0.001212397, 0.001212447, 0.001212359, 0.001212341, 
    0.001212353, 0.001212303, 0.00121245, 0.001212394, 0.001212821, 
    0.001212819, 0.001212807, 0.001212859, 0.001212862, 0.001212909, 
    0.001212867, 0.001212849, 0.001212803, 0.001212777, 0.001212751, 
    0.001212695, 0.001212634, 0.001212546, 0.001212481, 0.001212439, 
    0.001212464, 0.001212442, 0.001212467, 0.001212479, 0.001212348, 
    0.001212422, 0.00121231, 0.001212316, 0.001212367, 0.001212315, 
    0.001212817, 0.001212831, 0.001212882, 0.001212842, 0.001212914, 
    0.001212874, 0.001212852, 0.001212763, 0.001212742, 0.001212724, 
    0.001212688, 0.001212643, 0.001212563, 0.001212491, 0.001212427, 
    0.001212432, 0.00121243, 0.001212416, 0.001212451, 0.00121241, 
    0.001212404, 0.001212421, 0.001212317, 0.001212347, 0.001212316, 
    0.001212335, 0.001212826, 0.001212802, 0.001212815, 0.001212791, 
    0.001212809, 0.001212732, 0.001212709, 0.001212601, 0.001212644, 
    0.001212574, 0.001212636, 0.001212626, 0.001212573, 0.001212633, 
    0.001212496, 0.001212591, 0.001212416, 0.001212512, 0.00121241, 
    0.001212427, 0.001212398, 0.001212372, 0.001212338, 0.001212278, 
    0.001212292, 0.001212241, 0.001212766, 0.001212735, 0.001212737, 
    0.001212704, 0.00121268, 0.001212627, 0.001212543, 0.001212574, 
    0.001212516, 0.001212502, 0.001212592, 0.001212539, 0.001212714, 
    0.001212687, 0.001212702, 0.001212764, 0.001212568, 0.001212669, 
    0.00121248, 0.001212536, 0.001212376, 0.001212456, 0.0012123, 
    0.001212235, 0.001212171, 0.0012121, 0.001212717, 0.001212738, 0.0012127, 
    0.001212649, 0.001212598, 0.001212533, 0.001212526, 0.001212514, 
    0.00121248, 0.001212454, 0.001212511, 0.001212447, 0.001212682, 
    0.001212559, 0.001212747, 0.001212692, 0.001212651, 0.001212668, 
    0.001212577, 0.001212556, 0.00121247, 0.001212515, 0.001212252, 
    0.001212368, 0.001212044, 0.001212134, 0.001212746, 0.001212717, 
    0.001212618, 0.001212665, 0.001212528, 0.001212493, 0.001212466, 
    0.001212432, 0.001212427, 0.001212407, 0.00121244, 0.001212408, 
    0.001212533, 0.001212476, 0.001212628, 0.001212592, 0.001212608, 
    0.001212627, 0.00121257, 0.001212509, 0.001212506, 0.001212487, 
    0.001212437, 0.001212528, 0.00121224, 0.001212419, 0.001212686, 
    0.001212632, 0.001212623, 0.001212644, 0.001212497, 0.001212551, 
    0.001212407, 0.001212446, 0.001212383, 0.001212414, 0.001212419, 
    0.001212459, 0.001212484, 0.001212549, 0.001212601, 0.00121264, 
    0.001212631, 0.001212587, 0.001212505, 0.001212428, 0.001212445, 
    0.001212387, 0.001212538, 0.001212475, 0.001212499, 0.001212435, 
    0.001212575, 0.00121246, 0.001212605, 0.001212592, 0.001212552, 
    0.001212472, 0.001212452, 0.001212434, 0.001212445, 0.001212502, 
    0.001212513, 0.001212553, 0.001212565, 0.001212595, 0.00121262, 
    0.001212597, 0.001212573, 0.001212502, 0.00121244, 0.001212372, 
    0.001212354, 0.001212278, 0.001212342, 0.001212239, 0.00121233, 
    0.001212171, 0.001212451, 0.001212329, 0.00121255, 0.001212526, 
    0.001212483, 0.001212384, 0.001212436, 0.001212374, 0.001212513, 
    0.001212586, 0.001212603, 0.001212638, 0.001212603, 0.001212605, 
    0.001212571, 0.001212582, 0.0012125, 0.001212545, 0.001212419, 
    0.001212375, 0.001212246, 0.001212169, 0.001212088, 0.001212053, 
    0.001212042, 0.001212038 ;

 QBOT =
  0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_NODYNLNDUSE =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_R =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  3.284727e-06, 3.290784e-06, 3.289606e-06, 3.294489e-06, 3.291784e-06, 
    3.294977e-06, 3.285955e-06, 3.291024e-06, 3.287787e-06, 3.285273e-06, 
    3.303962e-06, 3.294707e-06, 3.313613e-06, 3.307686e-06, 3.323243e-06, 
    3.312689e-06, 3.32525e-06, 3.322958e-06, 3.329868e-06, 3.327887e-06, 
    3.336739e-06, 3.330783e-06, 3.341345e-06, 3.335317e-06, 3.336258e-06, 
    3.330586e-06, 3.296568e-06, 3.302808e-06, 3.296199e-06, 3.297088e-06, 
    3.296689e-06, 3.291839e-06, 3.289387e-06, 3.284266e-06, 3.285196e-06, 
    3.288958e-06, 3.297488e-06, 3.294596e-06, 3.301894e-06, 3.301729e-06, 
    3.30987e-06, 3.306195e-06, 3.320556e-06, 3.316013e-06, 3.32797e-06, 
    3.325116e-06, 3.327835e-06, 3.327011e-06, 3.327846e-06, 3.323662e-06, 
    3.325453e-06, 3.321776e-06, 3.306883e-06, 3.311064e-06, 3.298612e-06, 
    3.291141e-06, 3.286177e-06, 3.282659e-06, 3.283156e-06, 3.284103e-06, 
    3.28898e-06, 3.293571e-06, 3.297062e-06, 3.299399e-06, 3.301705e-06, 
    3.308686e-06, 3.312393e-06, 3.321347e-06, 3.319844e-06, 3.322392e-06, 
    3.324832e-06, 3.328931e-06, 3.328256e-06, 3.330063e-06, 3.322326e-06, 
    3.327465e-06, 3.318988e-06, 3.321303e-06, 3.302326e-06, 3.295376e-06, 
    3.292421e-06, 3.289832e-06, 3.283538e-06, 3.287882e-06, 3.286169e-06, 
    3.290249e-06, 3.292843e-06, 3.29156e-06, 3.299463e-06, 3.296389e-06, 
    3.312613e-06, 3.305614e-06, 3.324548e-06, 3.320153e-06, 3.325603e-06, 
    3.32282e-06, 3.327588e-06, 3.323297e-06, 3.330737e-06, 3.332359e-06, 
    3.33125e-06, 3.335515e-06, 3.323059e-06, 3.327834e-06, 3.291524e-06, 
    3.291733e-06, 3.292709e-06, 3.288422e-06, 3.288161e-06, 3.284241e-06, 
    3.287729e-06, 3.289215e-06, 3.292993e-06, 3.29522e-06, 3.297339e-06, 
    3.302005e-06, 3.307219e-06, 3.314534e-06, 3.320437e-06, 3.323979e-06, 
    3.321807e-06, 3.323725e-06, 3.321581e-06, 3.320577e-06, 3.33175e-06, 
    3.325469e-06, 3.3349e-06, 3.334378e-06, 3.330106e-06, 3.334437e-06, 
    3.291881e-06, 3.290676e-06, 3.286497e-06, 3.289767e-06, 3.283814e-06, 
    3.287144e-06, 3.28906e-06, 3.296453e-06, 3.298077e-06, 3.299583e-06, 
    3.302561e-06, 3.306383e-06, 3.313105e-06, 3.319602e-06, 3.324975e-06, 
    3.324581e-06, 3.324719e-06, 3.32592e-06, 3.322945e-06, 3.326409e-06, 
    3.32699e-06, 3.32547e-06, 3.334308e-06, 3.33178e-06, 3.334367e-06, 
    3.332721e-06, 3.291068e-06, 3.293093e-06, 3.291999e-06, 3.294053e-06, 
    3.292607e-06, 3.29904e-06, 3.300972e-06, 3.310026e-06, 3.306308e-06, 
    3.31223e-06, 3.306909e-06, 3.307851e-06, 3.31242e-06, 3.307197e-06, 
    3.319277e-06, 3.310874e-06, 3.325967e-06, 3.317543e-06, 3.326456e-06, 
    3.324951e-06, 3.327443e-06, 3.329676e-06, 3.33249e-06, 3.337687e-06, 
    3.336483e-06, 3.340837e-06, 3.296105e-06, 3.298727e-06, 3.298497e-06, 
    3.301245e-06, 3.303277e-06, 3.307689e-06, 3.31478e-06, 3.312111e-06, 
    3.317014e-06, 3.318632e-06, 3.310552e-06, 3.31512e-06, 3.300484e-06, 
    3.302843e-06, 3.301439e-06, 3.29631e-06, 3.312724e-06, 3.304288e-06, 
    3.320524e-06, 3.315303e-06, 3.329358e-06, 3.32267e-06, 3.33582e-06, 
    3.341457e-06, 3.346782e-06, 3.353009e-06, 3.30016e-06, 3.298377e-06, 
    3.301572e-06, 3.305993e-06, 3.310106e-06, 3.315582e-06, 3.316144e-06, 
    3.317171e-06, 3.32047e-06, 3.322714e-06, 3.317494e-06, 3.323277e-06, 
    3.303387e-06, 3.313459e-06, 3.297702e-06, 3.302437e-06, 3.305733e-06, 
    3.304288e-06, 3.311807e-06, 3.313582e-06, 3.321443e-06, 3.31707e-06, 
    3.340063e-06, 3.330146e-06, 3.357767e-06, 3.350017e-06, 3.297754e-06, 
    3.300155e-06, 3.30852e-06, 3.304537e-06, 3.315949e-06, 3.319399e-06, 
    3.321695e-06, 3.32463e-06, 3.324948e-06, 3.32669e-06, 3.323837e-06, 
    3.326578e-06, 3.315594e-06, 3.320846e-06, 3.307564e-06, 3.310636e-06, 
    3.309223e-06, 3.307673e-06, 3.312459e-06, 3.318198e-06, 3.31831e-06, 
    3.319952e-06, 3.324577e-06, 3.315995e-06, 3.34134e-06, 3.326044e-06, 
    3.302774e-06, 3.307403e-06, 3.308067e-06, 3.306272e-06, 3.319116e-06, 
    3.314051e-06, 3.326648e-06, 3.323408e-06, 3.328719e-06, 3.326078e-06, 
    3.32569e-06, 3.322303e-06, 3.320197e-06, 3.314254e-06, 3.309944e-06, 
    3.306532e-06, 3.307325e-06, 3.311074e-06, 3.318512e-06, 3.324976e-06, 
    3.323558e-06, 3.328315e-06, 3.31512e-06, 3.321009e-06, 3.318974e-06, 
    3.324285e-06, 3.31204e-06, 3.322548e-06, 3.309522e-06, 3.310606e-06, 
    3.313963e-06, 3.321365e-06, 3.322869e-06, 3.324473e-06, 3.323484e-06, 
    3.318686e-06, 3.31727e-06, 3.313882e-06, 3.312947e-06, 3.31037e-06, 
    3.308238e-06, 3.310186e-06, 3.312232e-06, 3.318689e-06, 3.323953e-06, 
    3.329708e-06, 3.331119e-06, 3.337855e-06, 3.332366e-06, 3.341424e-06, 
    3.333715e-06, 3.347079e-06, 3.323126e-06, 3.333495e-06, 3.314117e-06, 
    3.316128e-06, 3.320403e-06, 3.328786e-06, 3.32426e-06, 3.329556e-06, 
    3.317239e-06, 3.311203e-06, 3.309646e-06, 3.306739e-06, 3.309712e-06, 
    3.30947e-06, 3.312318e-06, 3.311403e-06, 3.318883e-06, 3.31457e-06, 
    3.325679e-06, 3.329514e-06, 3.340379e-06, 3.34706e-06, 3.353884e-06, 
    3.356899e-06, 3.357819e-06, 3.358203e-06 ;

 QVEGE =
  -7.794849e-07, -7.790419e-07, -7.79126e-07, -7.787725e-07, -7.789653e-07, 
    -7.787362e-07, -7.793911e-07, -7.790279e-07, -7.792576e-07, 
    -7.794395e-07, -7.780956e-07, -7.787557e-07, -7.773741e-07, 
    -7.778003e-07, -7.767163e-07, -7.77446e-07, -7.765662e-07, -7.767281e-07, 
    -7.762169e-07, -7.763631e-07, -7.757253e-07, -7.761492e-07, 
    -7.753773e-07, -7.758217e-07, -7.757559e-07, -7.761647e-07, 
    -7.786142e-07, -7.781803e-07, -7.786419e-07, -7.785796e-07, 
    -7.786055e-07, -7.789646e-07, -7.79151e-07, -7.795124e-07, -7.794452e-07, 
    -7.791763e-07, -7.785514e-07, -7.787579e-07, -7.782185e-07, 
    -7.782305e-07, -7.776397e-07, -7.779063e-07, -7.769048e-07, 
    -7.771869e-07, -7.763568e-07, -7.765684e-07, -7.763684e-07, 
    -7.764279e-07, -7.763676e-07, -7.76677e-07, -7.765451e-07, -7.768139e-07, 
    -7.778582e-07, -7.775546e-07, -7.784658e-07, -7.790281e-07, 
    -7.793769e-07, -7.796305e-07, -7.795947e-07, -7.795283e-07, 
    -7.791749e-07, -7.788333e-07, -7.785751e-07, -7.784033e-07, 
    -7.782324e-07, -7.777431e-07, -7.774633e-07, -7.768516e-07, 
    -7.769549e-07, -7.767737e-07, -7.76589e-07, -7.762885e-07, -7.763369e-07, 
    -7.762062e-07, -7.767728e-07, -7.763995e-07, -7.770155e-07, 
    -7.768485e-07, -7.782173e-07, -7.787008e-07, -7.789324e-07, -7.79111e-07, 
    -7.795678e-07, -7.792543e-07, -7.793788e-07, -7.790758e-07, 
    -7.788873e-07, -7.789793e-07, -7.783985e-07, -7.78626e-07, -7.774467e-07, 
    -7.779536e-07, -7.766105e-07, -7.769331e-07, -7.765319e-07, 
    -7.767353e-07, -7.76389e-07, -7.767006e-07, -7.761549e-07, -7.760391e-07, 
    -7.76119e-07, -7.758013e-07, -7.767187e-07, -7.763714e-07, -7.789833e-07, 
    -7.789685e-07, -7.788958e-07, -7.792155e-07, -7.792332e-07, 
    -7.795157e-07, -7.792616e-07, -7.791557e-07, -7.788738e-07, 
    -7.787127e-07, -7.78557e-07, -7.782134e-07, -7.778379e-07, -7.773021e-07, 
    -7.769125e-07, -7.766503e-07, -7.768091e-07, -7.766691e-07, 
    -7.768268e-07, -7.768992e-07, -7.760846e-07, -7.765458e-07, 
    -7.758471e-07, -7.758848e-07, -7.762043e-07, -7.758805e-07, 
    -7.789576e-07, -7.790438e-07, -7.793524e-07, -7.791109e-07, -7.79546e-07, 
    -7.793067e-07, -7.79171e-07, -7.786281e-07, -7.785008e-07, -7.783925e-07, 
    -7.781711e-07, -7.778929e-07, -7.774056e-07, -7.769769e-07, 
    -7.765769e-07, -7.766056e-07, -7.765958e-07, -7.765095e-07, 
    -7.767276e-07, -7.764733e-07, -7.764336e-07, -7.765422e-07, -7.7589e-07, 
    -7.760765e-07, -7.758857e-07, -7.760063e-07, -7.79015e-07, -7.788684e-07, 
    -7.789481e-07, -7.787999e-07, -7.789068e-07, -7.784393e-07, 
    -7.782988e-07, -7.77636e-07, -7.779001e-07, -7.774709e-07, -7.778542e-07, 
    -7.777882e-07, -7.774701e-07, -7.778314e-07, -7.770067e-07, 
    -7.775776e-07, -7.765061e-07, -7.770924e-07, -7.764698e-07, 
    -7.765786e-07, -7.763952e-07, -7.762339e-07, -7.760246e-07, 
    -7.756464e-07, -7.757328e-07, -7.754102e-07, -7.786466e-07, 
    -7.784585e-07, -7.784693e-07, -7.782679e-07, -7.781209e-07, 
    -7.777961e-07, -7.772804e-07, -7.774726e-07, -7.771129e-07, 
    -7.770446e-07, -7.775856e-07, -7.772582e-07, -7.783279e-07, 
    -7.781606e-07, -7.782557e-07, -7.786352e-07, -7.774364e-07, 
    -7.780541e-07, -7.769072e-07, -7.772407e-07, -7.762577e-07, 
    -7.767553e-07, -7.757818e-07, -7.753774e-07, -7.749671e-07, 
    -7.745174e-07, -7.783493e-07, -7.78478e-07, -7.782422e-07, -7.779291e-07, 
    -7.776218e-07, -7.772214e-07, -7.771771e-07, -7.771036e-07, 
    -7.769075e-07, -7.767435e-07, -7.77086e-07, -7.767018e-07, -7.781338e-07, 
    -7.7738e-07, -7.78532e-07, -7.781916e-07, -7.779449e-07, -7.780471e-07, 
    -7.774931e-07, -7.773643e-07, -7.768429e-07, -7.771085e-07, 
    -7.754827e-07, -7.762081e-07, -7.741532e-07, -7.747368e-07, 
    -7.785243e-07, -7.783469e-07, -7.777414e-07, -7.78028e-07, -7.771915e-07, 
    -7.769891e-07, -7.768174e-07, -7.76607e-07, -7.765798e-07, -7.76454e-07, 
    -7.766607e-07, -7.7646e-07, -7.772206e-07, -7.768818e-07, -7.778036e-07, 
    -7.775829e-07, -7.776824e-07, -7.777959e-07, -7.774461e-07, 
    -7.770842e-07, -7.770669e-07, -7.769514e-07, -7.766418e-07, 
    -7.771879e-07, -7.754062e-07, -7.765294e-07, -7.781543e-07, 
    -7.778282e-07, -7.7777e-07, -7.778985e-07, -7.7701e-07, -7.773327e-07, 
    -7.764558e-07, -7.766923e-07, -7.763019e-07, -7.76497e-07, -7.765261e-07, 
    -7.767737e-07, -7.769299e-07, -7.773197e-07, -7.776345e-07, 
    -7.778787e-07, -7.778212e-07, -7.775525e-07, -7.770597e-07, 
    -7.765817e-07, -7.76688e-07, -7.763315e-07, -7.772527e-07, -7.768739e-07, 
    -7.770245e-07, -7.766296e-07, -7.774798e-07, -7.767855e-07, 
    -7.776604e-07, -7.775819e-07, -7.77339e-07, -7.768544e-07, -7.767321e-07, 
    -7.766185e-07, -7.766866e-07, -7.770453e-07, -7.770975e-07, 
    -7.773426e-07, -7.774149e-07, -7.775982e-07, -7.777544e-07, 
    -7.776141e-07, -7.774686e-07, -7.770412e-07, -7.766573e-07, -7.76233e-07, 
    -7.761251e-07, -7.756498e-07, -7.760502e-07, -7.754019e-07, 
    -7.759733e-07, -7.749715e-07, -7.767309e-07, -7.759706e-07, 
    -7.773248e-07, -7.771776e-07, -7.769228e-07, -7.763097e-07, 
    -7.766313e-07, -7.762504e-07, -7.770989e-07, -7.775479e-07, 
    -7.776521e-07, -7.778656e-07, -7.776472e-07, -7.776646e-07, 
    -7.774559e-07, -7.775224e-07, -7.770267e-07, -7.77292e-07, -7.765294e-07, 
    -7.762511e-07, -7.754476e-07, -7.74957e-07, -7.744388e-07, -7.742142e-07, 
    -7.741448e-07, -7.741164e-07 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  84.8408, 84.8404, 84.84048, 84.84018, 84.84034, 84.84015, 84.84071, 
    84.84039, 84.84059, 84.84076, 84.83964, 84.84016, 84.83916, 84.83945, 
    84.83832, 84.83921, 84.83823, 84.83833, 84.83804, 84.83812, 84.83775, 
    84.838, 84.83757, 84.83781, 84.83778, 84.83801, 84.84005, 84.8397, 
    84.84007, 84.84002, 84.84004, 84.84034, 84.84049, 84.84082, 84.84076, 
    84.84052, 84.84, 84.84016, 84.83974, 84.83975, 84.83934, 84.83952, 
    84.83844, 84.83906, 84.83812, 84.83824, 84.83812, 84.83816, 84.83812, 
    84.8383, 84.83823, 84.83839, 84.83949, 84.83929, 84.83993, 84.84039, 
    84.8407, 84.84093, 84.8409, 84.84084, 84.84052, 84.84023, 84.84002, 
    84.83988, 84.83975, 84.8394, 84.83923, 84.8384, 84.83847, 84.83836, 
    84.83825, 84.83807, 84.8381, 84.83803, 84.83836, 84.83813, 84.83851, 
    84.8384, 84.83972, 84.84012, 84.8403, 84.84046, 84.84087, 84.84059, 
    84.8407, 84.84044, 84.84027, 84.84035, 84.83988, 84.84006, 84.83921, 
    84.83955, 84.83826, 84.83846, 84.83822, 84.83834, 84.83813, 84.83832, 
    84.838, 84.83794, 84.83798, 84.83781, 84.83833, 84.83812, 84.84035, 
    84.84034, 84.84028, 84.84055, 84.84057, 84.84083, 84.8406, 84.8405, 
    84.84026, 84.84013, 84.84, 84.83974, 84.83947, 84.83913, 84.83845, 
    84.83829, 84.83839, 84.83829, 84.83839, 84.83844, 84.83796, 84.83823, 
    84.83783, 84.83785, 84.83803, 84.83784, 84.84033, 84.84041, 84.84068, 
    84.84047, 84.84085, 84.84064, 84.84052, 84.84006, 84.83996, 84.83987, 
    84.83971, 84.83951, 84.83919, 84.83848, 84.83824, 84.83826, 84.83826, 
    84.8382, 84.83833, 84.83818, 84.83816, 84.83823, 84.83785, 84.83796, 
    84.83785, 84.83792, 84.84039, 84.84026, 84.84032, 84.8402, 84.84029, 
    84.8399, 84.8398, 84.83933, 84.83952, 84.83923, 84.83949, 84.83944, 
    84.83923, 84.83947, 84.83849, 84.83929, 84.8382, 84.83899, 84.83818, 
    84.83824, 84.83813, 84.83804, 84.83793, 84.83772, 84.83777, 84.83759, 
    84.84008, 84.83993, 84.83994, 84.83978, 84.83967, 84.83945, 84.83911, 
    84.83923, 84.83901, 84.83852, 84.83931, 84.8391, 84.83982, 84.83969, 
    84.83977, 84.84007, 84.8392, 84.83961, 84.83844, 84.83909, 84.83806, 
    84.83835, 84.83779, 84.83757, 84.83736, 84.83714, 84.83984, 84.83994, 
    84.83976, 84.83953, 84.83933, 84.83907, 84.83905, 84.839, 84.83844, 
    84.83834, 84.83899, 84.83832, 84.83967, 84.83917, 84.83998, 84.83971, 
    84.83955, 84.83961, 84.83925, 84.83916, 84.8384, 84.839, 84.83762, 
    84.83803, 84.83698, 84.83725, 84.83998, 84.83984, 84.83941, 84.8396, 
    84.83906, 84.83849, 84.83839, 84.83826, 84.83825, 84.83817, 84.83829, 
    84.83817, 84.83907, 84.83842, 84.83945, 84.8393, 84.83937, 84.83945, 
    84.83922, 84.83855, 84.83854, 84.83846, 84.83826, 84.83906, 84.83758, 
    84.8382, 84.83969, 84.83946, 84.83943, 84.83952, 84.8385, 84.83914, 
    84.83817, 84.83831, 84.83808, 84.8382, 84.83821, 84.83836, 84.83846, 
    84.83913, 84.83934, 84.8395, 84.83946, 84.83929, 84.83853, 84.83824, 
    84.83831, 84.8381, 84.8391, 84.83842, 84.83851, 84.83827, 84.83924, 
    84.83836, 84.83936, 84.8393, 84.83915, 84.8384, 84.83833, 84.83826, 
    84.83831, 84.83852, 84.839, 84.83915, 84.8392, 84.83932, 84.83942, 
    84.83932, 84.83923, 84.83852, 84.83829, 84.83804, 84.83798, 84.83772, 
    84.83794, 84.83758, 84.83788, 84.83736, 84.83833, 84.83789, 84.83914, 
    84.83905, 84.83845, 84.83808, 84.83827, 84.83805, 84.839, 84.83928, 
    84.83935, 84.83949, 84.83935, 84.83936, 84.83923, 84.83926, 84.83852, 
    84.83912, 84.83821, 84.83805, 84.83761, 84.83736, 84.8371, 84.837, 
    84.83697, 84.83696 ;

 RH2M_R =
  84.8408, 84.8404, 84.84048, 84.84018, 84.84034, 84.84015, 84.84071, 
    84.84039, 84.84059, 84.84076, 84.83964, 84.84016, 84.83916, 84.83945, 
    84.83832, 84.83921, 84.83823, 84.83833, 84.83804, 84.83812, 84.83775, 
    84.838, 84.83757, 84.83781, 84.83778, 84.83801, 84.84005, 84.8397, 
    84.84007, 84.84002, 84.84004, 84.84034, 84.84049, 84.84082, 84.84076, 
    84.84052, 84.84, 84.84016, 84.83974, 84.83975, 84.83934, 84.83952, 
    84.83844, 84.83906, 84.83812, 84.83824, 84.83812, 84.83816, 84.83812, 
    84.8383, 84.83823, 84.83839, 84.83949, 84.83929, 84.83993, 84.84039, 
    84.8407, 84.84093, 84.8409, 84.84084, 84.84052, 84.84023, 84.84002, 
    84.83988, 84.83975, 84.8394, 84.83923, 84.8384, 84.83847, 84.83836, 
    84.83825, 84.83807, 84.8381, 84.83803, 84.83836, 84.83813, 84.83851, 
    84.8384, 84.83972, 84.84012, 84.8403, 84.84046, 84.84087, 84.84059, 
    84.8407, 84.84044, 84.84027, 84.84035, 84.83988, 84.84006, 84.83921, 
    84.83955, 84.83826, 84.83846, 84.83822, 84.83834, 84.83813, 84.83832, 
    84.838, 84.83794, 84.83798, 84.83781, 84.83833, 84.83812, 84.84035, 
    84.84034, 84.84028, 84.84055, 84.84057, 84.84083, 84.8406, 84.8405, 
    84.84026, 84.84013, 84.84, 84.83974, 84.83947, 84.83913, 84.83845, 
    84.83829, 84.83839, 84.83829, 84.83839, 84.83844, 84.83796, 84.83823, 
    84.83783, 84.83785, 84.83803, 84.83784, 84.84033, 84.84041, 84.84068, 
    84.84047, 84.84085, 84.84064, 84.84052, 84.84006, 84.83996, 84.83987, 
    84.83971, 84.83951, 84.83919, 84.83848, 84.83824, 84.83826, 84.83826, 
    84.8382, 84.83833, 84.83818, 84.83816, 84.83823, 84.83785, 84.83796, 
    84.83785, 84.83792, 84.84039, 84.84026, 84.84032, 84.8402, 84.84029, 
    84.8399, 84.8398, 84.83933, 84.83952, 84.83923, 84.83949, 84.83944, 
    84.83923, 84.83947, 84.83849, 84.83929, 84.8382, 84.83899, 84.83818, 
    84.83824, 84.83813, 84.83804, 84.83793, 84.83772, 84.83777, 84.83759, 
    84.84008, 84.83993, 84.83994, 84.83978, 84.83967, 84.83945, 84.83911, 
    84.83923, 84.83901, 84.83852, 84.83931, 84.8391, 84.83982, 84.83969, 
    84.83977, 84.84007, 84.8392, 84.83961, 84.83844, 84.83909, 84.83806, 
    84.83835, 84.83779, 84.83757, 84.83736, 84.83714, 84.83984, 84.83994, 
    84.83976, 84.83953, 84.83933, 84.83907, 84.83905, 84.839, 84.83844, 
    84.83834, 84.83899, 84.83832, 84.83967, 84.83917, 84.83998, 84.83971, 
    84.83955, 84.83961, 84.83925, 84.83916, 84.8384, 84.839, 84.83762, 
    84.83803, 84.83698, 84.83725, 84.83998, 84.83984, 84.83941, 84.8396, 
    84.83906, 84.83849, 84.83839, 84.83826, 84.83825, 84.83817, 84.83829, 
    84.83817, 84.83907, 84.83842, 84.83945, 84.8393, 84.83937, 84.83945, 
    84.83922, 84.83855, 84.83854, 84.83846, 84.83826, 84.83906, 84.83758, 
    84.8382, 84.83969, 84.83946, 84.83943, 84.83952, 84.8385, 84.83914, 
    84.83817, 84.83831, 84.83808, 84.8382, 84.83821, 84.83836, 84.83846, 
    84.83913, 84.83934, 84.8395, 84.83946, 84.83929, 84.83853, 84.83824, 
    84.83831, 84.8381, 84.8391, 84.83842, 84.83851, 84.83827, 84.83924, 
    84.83836, 84.83936, 84.8393, 84.83915, 84.8384, 84.83833, 84.83826, 
    84.83831, 84.83852, 84.839, 84.83915, 84.8392, 84.83932, 84.83942, 
    84.83932, 84.83923, 84.83852, 84.83829, 84.83804, 84.83798, 84.83772, 
    84.83794, 84.83758, 84.83788, 84.83736, 84.83833, 84.83789, 84.83914, 
    84.83905, 84.83845, 84.83808, 84.83827, 84.83805, 84.839, 84.83928, 
    84.83935, 84.83949, 84.83935, 84.83936, 84.83923, 84.83926, 84.83852, 
    84.83912, 84.83821, 84.83805, 84.83761, 84.83736, 84.8371, 84.837, 
    84.83697, 84.83696 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.00046391, 0.0004658502, 0.0004654728, 0.0004670377, 0.0004661695, 
    0.0004671942, 0.000464303, 0.0004659269, 0.0004648901, 0.000464084, 
    0.0004700741, 0.000467107, 0.0004731544, 0.0004712626, 0.0004760139, 
    0.00047286, 0.0004766496, 0.0004759225, 0.00047811, 0.0004774832, 
    0.0004802814, 0.0004783991, 0.0004817312, 0.0004798316, 0.0004801288, 
    0.0004783367, 0.0004677043, 0.0004697052, 0.0004675857, 0.0004678711, 
    0.0004677429, 0.0004661873, 0.0004654035, 0.000463761, 0.000464059, 
    0.0004652652, 0.000467999, 0.0004670708, 0.0004694092, 0.0004693564, 
    0.0004719595, 0.0004707858, 0.0004751604, 0.000473917, 0.0004775093, 
    0.0004766059, 0.0004774668, 0.0004772056, 0.0004774701, 0.0004761452, 
    0.0004767128, 0.0004755468, 0.0004710064, 0.0004723413, 0.0004683595, 
    0.0004659651, 0.000464374, 0.0004632451, 0.0004634045, 0.0004637089, 
    0.0004652722, 0.0004667417, 0.0004678616, 0.0004686106, 0.0004693486, 
    0.0004715832, 0.0004727651, 0.0004754118, 0.0004749339, 0.0004757432, 
    0.000476516, 0.0004778136, 0.0004776, 0.0004781717, 0.0004757213, 
    0.0004773499, 0.0004746613, 0.0004753967, 0.0004695507, 0.0004673214, 
    0.0004663744, 0.0004655449, 0.0004635272, 0.0004649206, 0.0004643713, 
    0.0004656777, 0.0004665079, 0.0004660971, 0.000468631, 0.0004676459, 
    0.0004728351, 0.0004706001, 0.0004764259, 0.0004750319, 0.0004767598, 
    0.000475878, 0.0004773889, 0.000476029, 0.0004783843, 0.0004788972, 
    0.0004785466, 0.0004798927, 0.0004759533, 0.0004774664, 0.000466086, 
    0.000466153, 0.0004664649, 0.0004650935, 0.0004650096, 0.0004637525, 
    0.0004648708, 0.0004653471, 0.0004665558, 0.0004672708, 0.0004679504, 
    0.0004694447, 0.0004711134, 0.0004734464, 0.0004751222, 0.0004762454, 
    0.0004755565, 0.0004761646, 0.0004754847, 0.000475166, 0.0004787049, 
    0.0004767179, 0.0004796989, 0.0004795339, 0.0004781848, 0.0004795523, 
    0.0004661999, 0.0004658144, 0.0004644764, 0.0004655234, 0.0004636155, 
    0.0004646835, 0.0004652976, 0.0004676666, 0.0004681868, 0.0004686695, 
    0.0004696224, 0.0004708455, 0.0004729909, 0.0004748572, 0.0004765607, 
    0.0004764358, 0.0004764797, 0.0004768602, 0.0004759175, 0.0004770149, 
    0.000477199, 0.0004767174, 0.0004795117, 0.0004787134, 0.0004795302, 
    0.0004790103, 0.0004659396, 0.000466588, 0.0004662375, 0.0004668965, 
    0.0004664322, 0.0004684962, 0.0004691149, 0.0004720097, 0.0004708214, 
    0.0004727122, 0.0004710133, 0.0004713144, 0.0004727741, 0.0004711049, 
    0.0004747543, 0.0004722804, 0.0004768749, 0.0004744052, 0.0004770296, 
    0.0004765528, 0.0004773419, 0.0004780487, 0.0004789376, 0.000480578, 
    0.000480198, 0.0004815697, 0.0004675545, 0.0004683955, 0.0004683213, 
    0.0004692012, 0.000469852, 0.0004712624, 0.0004735244, 0.0004726737, 
    0.000474235, 0.0004745485, 0.0004721761, 0.0004736329, 0.0004689577, 
    0.0004697132, 0.0004692632, 0.0004676201, 0.0004728694, 0.0004701756, 
    0.0004751492, 0.0004736901, 0.0004779478, 0.0004758306, 0.0004799889, 
    0.0004817667, 0.0004834389, 0.0004853937, 0.0004688543, 0.0004682827, 
    0.0004693057, 0.0004707214, 0.0004720342, 0.0004737798, 0.0004739582, 
    0.0004742852, 0.000475132, 0.0004758441, 0.0004743886, 0.0004760225, 
    0.0004698886, 0.0004731031, 0.0004680661, 0.0004695832, 0.0004706371, 
    0.0004701746, 0.0004725757, 0.0004731415, 0.000475441, 0.0004742522, 
    0.0004813279, 0.0004781978, 0.0004868813, 0.0004844552, 0.000468083, 
    0.000468852, 0.0004715284, 0.000470255, 0.0004738961, 0.0004747923, 
    0.0004755206, 0.0004764519, 0.0004765522, 0.000477104, 0.0004761997, 
    0.0004770681, 0.0004737829, 0.000475251, 0.0004712217, 0.0004722025, 
    0.0004717512, 0.0004712562, 0.0004727835, 0.0004744109, 0.0004744454, 
    0.0004749671, 0.000476438, 0.0004739098, 0.0004817322, 0.000476902, 
    0.0004696905, 0.0004711719, 0.0004713831, 0.0004708093, 0.0004747023, 
    0.0004732918, 0.0004770905, 0.0004760638, 0.0004777457, 0.00047691, 
    0.0004767869, 0.0004757133, 0.0004750449, 0.0004733561, 0.0004719818, 
    0.0004708919, 0.0004711451, 0.0004723424, 0.0004745102, 0.0004765608, 
    0.0004761115, 0.0004776172, 0.0004736309, 0.0004753027, 0.0004746565, 
    0.0004763409, 0.0004726509, 0.000475795, 0.0004718472, 0.0004721932, 
    0.0004732637, 0.0004754171, 0.000475893, 0.0004764017, 0.0004760876, 
    0.0004745657, 0.0004743161, 0.0004732372, 0.0004729394, 0.0004721173, 
    0.0004714366, 0.0004720585, 0.0004727115, 0.0004745657, 0.0004762367, 
    0.0004780581, 0.0004785037, 0.0004806323, 0.0004788998, 0.0004817588, 
    0.0004793286, 0.0004835348, 0.0004759766, 0.0004792578, 0.0004733123, 
    0.0004739528, 0.0004751115, 0.0004777684, 0.0004763337, 0.0004780113, 
    0.0004743063, 0.0004723839, 0.0004718862, 0.0004709581, 0.0004719073, 
    0.00047183, 0.0004727383, 0.0004724464, 0.0004746271, 0.0004734557, 
    0.0004767831, 0.0004779973, 0.0004814254, 0.0004835267, 0.000485665, 
    0.000486609, 0.0004868963, 0.0004870164 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.280768e-14, 3.289606e-14, 3.287889e-14, 3.295011e-14, 3.291062e-14, 
    3.295724e-14, 3.282561e-14, 3.289956e-14, 3.285237e-14, 3.281565e-14, 
    3.308812e-14, 3.295329e-14, 3.322804e-14, 3.314221e-14, 3.335767e-14, 
    3.321467e-14, 3.338648e-14, 3.335358e-14, 3.345264e-14, 3.342428e-14, 
    3.35508e-14, 3.346573e-14, 3.361635e-14, 3.353051e-14, 3.354393e-14, 
    3.346292e-14, 3.298046e-14, 3.307133e-14, 3.297507e-14, 3.298804e-14, 
    3.298223e-14, 3.291142e-14, 3.287571e-14, 3.280093e-14, 3.281452e-14, 
    3.286945e-14, 3.299387e-14, 3.295167e-14, 3.305803e-14, 3.305563e-14, 
    3.317386e-14, 3.312057e-14, 3.331904e-14, 3.32627e-14, 3.342546e-14, 
    3.338455e-14, 3.342354e-14, 3.341172e-14, 3.342369e-14, 3.336368e-14, 
    3.33894e-14, 3.333658e-14, 3.313055e-14, 3.319115e-14, 3.301026e-14, 
    3.290126e-14, 3.282885e-14, 3.277741e-14, 3.278469e-14, 3.279855e-14, 
    3.286977e-14, 3.29367e-14, 3.298766e-14, 3.302173e-14, 3.305528e-14, 
    3.315671e-14, 3.32104e-14, 3.333042e-14, 3.330879e-14, 3.334545e-14, 
    3.338048e-14, 3.343924e-14, 3.342957e-14, 3.345544e-14, 3.33445e-14, 
    3.341824e-14, 3.329647e-14, 3.332979e-14, 3.306431e-14, 3.296306e-14, 
    3.291991e-14, 3.288218e-14, 3.279028e-14, 3.285376e-14, 3.282873e-14, 
    3.288826e-14, 3.292605e-14, 3.290737e-14, 3.302266e-14, 3.297785e-14, 
    3.321358e-14, 3.311213e-14, 3.33764e-14, 3.331324e-14, 3.339153e-14, 
    3.335159e-14, 3.342001e-14, 3.335844e-14, 3.346508e-14, 3.348826e-14, 
    3.347241e-14, 3.353331e-14, 3.335502e-14, 3.342353e-14, 3.290684e-14, 
    3.290989e-14, 3.29241e-14, 3.286163e-14, 3.285781e-14, 3.280056e-14, 
    3.285152e-14, 3.28732e-14, 3.292825e-14, 3.296078e-14, 3.29917e-14, 
    3.305965e-14, 3.313544e-14, 3.324134e-14, 3.331733e-14, 3.336824e-14, 
    3.333703e-14, 3.336458e-14, 3.333378e-14, 3.331934e-14, 3.347957e-14, 
    3.338963e-14, 3.352455e-14, 3.35171e-14, 3.345605e-14, 3.351794e-14, 
    3.291203e-14, 3.289449e-14, 3.283354e-14, 3.288124e-14, 3.279432e-14, 
    3.284298e-14, 3.287093e-14, 3.297877e-14, 3.300246e-14, 3.30244e-14, 
    3.306774e-14, 3.31233e-14, 3.322068e-14, 3.330531e-14, 3.338252e-14, 
    3.337687e-14, 3.337886e-14, 3.339609e-14, 3.335339e-14, 3.34031e-14, 
    3.341143e-14, 3.338963e-14, 3.35161e-14, 3.347999e-14, 3.351694e-14, 
    3.349343e-14, 3.29002e-14, 3.292971e-14, 3.291376e-14, 3.294374e-14, 
    3.292261e-14, 3.301649e-14, 3.304462e-14, 3.317613e-14, 3.31222e-14, 
    3.320803e-14, 3.313093e-14, 3.314459e-14, 3.321079e-14, 3.313511e-14, 
    3.330063e-14, 3.318842e-14, 3.339676e-14, 3.32848e-14, 3.340377e-14, 
    3.338219e-14, 3.341792e-14, 3.344991e-14, 3.349014e-14, 3.356429e-14, 
    3.354713e-14, 3.360912e-14, 3.297369e-14, 3.301193e-14, 3.300858e-14, 
    3.304859e-14, 3.307816e-14, 3.314224e-14, 3.324489e-14, 3.320631e-14, 
    3.327715e-14, 3.329134e-14, 3.318374e-14, 3.324981e-14, 3.303752e-14, 
    3.307184e-14, 3.305142e-14, 3.29767e-14, 3.321518e-14, 3.309287e-14, 
    3.331858e-14, 3.325245e-14, 3.344534e-14, 3.334945e-14, 3.353768e-14, 
    3.361797e-14, 3.369354e-14, 3.378166e-14, 3.303281e-14, 3.300683e-14, 
    3.305335e-14, 3.311763e-14, 3.317728e-14, 3.325648e-14, 3.326459e-14, 
    3.327942e-14, 3.33178e-14, 3.335007e-14, 3.328409e-14, 3.335816e-14, 
    3.307976e-14, 3.32258e-14, 3.2997e-14, 3.306594e-14, 3.311385e-14, 
    3.309286e-14, 3.320191e-14, 3.322758e-14, 3.333181e-14, 3.327796e-14, 
    3.359814e-14, 3.345664e-14, 3.384875e-14, 3.373936e-14, 3.299775e-14, 
    3.303273e-14, 3.31543e-14, 3.309648e-14, 3.326178e-14, 3.330239e-14, 
    3.333542e-14, 3.337759e-14, 3.338215e-14, 3.340713e-14, 3.336619e-14, 
    3.340552e-14, 3.325665e-14, 3.33232e-14, 3.314044e-14, 3.318495e-14, 
    3.316448e-14, 3.314201e-14, 3.321135e-14, 3.32851e-14, 3.32867e-14, 
    3.331034e-14, 3.337686e-14, 3.326245e-14, 3.361634e-14, 3.339791e-14, 
    3.307084e-14, 3.31381e-14, 3.314773e-14, 3.312168e-14, 3.329832e-14, 
    3.323436e-14, 3.340653e-14, 3.336003e-14, 3.34362e-14, 3.339836e-14, 
    3.339279e-14, 3.334416e-14, 3.331386e-14, 3.32373e-14, 3.317493e-14, 
    3.312547e-14, 3.313697e-14, 3.31913e-14, 3.328962e-14, 3.338255e-14, 
    3.33622e-14, 3.343042e-14, 3.32498e-14, 3.332556e-14, 3.329627e-14, 
    3.337262e-14, 3.320528e-14, 3.334772e-14, 3.316882e-14, 3.318452e-14, 
    3.32331e-14, 3.333068e-14, 3.33523e-14, 3.337532e-14, 3.336112e-14, 
    3.329212e-14, 3.328084e-14, 3.323192e-14, 3.32184e-14, 3.318111e-14, 
    3.315021e-14, 3.317843e-14, 3.320806e-14, 3.329216e-14, 3.336788e-14, 
    3.345036e-14, 3.347054e-14, 3.356671e-14, 3.348839e-14, 3.361755e-14, 
    3.35077e-14, 3.369778e-14, 3.3356e-14, 3.350452e-14, 3.323531e-14, 
    3.326437e-14, 3.331684e-14, 3.343718e-14, 3.337226e-14, 3.344819e-14, 
    3.32804e-14, 3.319316e-14, 3.317062e-14, 3.312847e-14, 3.317158e-14, 
    3.316808e-14, 3.320931e-14, 3.319606e-14, 3.329495e-14, 3.324186e-14, 
    3.339264e-14, 3.344759e-14, 3.360262e-14, 3.369748e-14, 3.379398e-14, 
    3.383652e-14, 3.384947e-14, 3.385488e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.090895e-14, 1.093837e-14, 1.093265e-14, 1.095636e-14, 1.094321e-14, 
    1.095873e-14, 1.091492e-14, 1.093953e-14, 1.092382e-14, 1.09116e-14, 
    1.100229e-14, 1.095742e-14, 1.104887e-14, 1.10203e-14, 1.109202e-14, 
    1.104442e-14, 1.110161e-14, 1.109065e-14, 1.112363e-14, 1.111419e-14, 
    1.11563e-14, 1.112799e-14, 1.117812e-14, 1.114955e-14, 1.115402e-14, 
    1.112705e-14, 1.096646e-14, 1.099671e-14, 1.096467e-14, 1.096898e-14, 
    1.096705e-14, 1.094348e-14, 1.093159e-14, 1.090671e-14, 1.091123e-14, 
    1.092951e-14, 1.097092e-14, 1.095688e-14, 1.099228e-14, 1.099148e-14, 
    1.103083e-14, 1.10131e-14, 1.107916e-14, 1.106041e-14, 1.111458e-14, 
    1.110096e-14, 1.111394e-14, 1.111001e-14, 1.111399e-14, 1.109402e-14, 
    1.110258e-14, 1.1085e-14, 1.101642e-14, 1.103659e-14, 1.097638e-14, 
    1.09401e-14, 1.0916e-14, 1.089888e-14, 1.09013e-14, 1.090591e-14, 
    1.092962e-14, 1.095189e-14, 1.096886e-14, 1.09802e-14, 1.099137e-14, 
    1.102512e-14, 1.104299e-14, 1.108295e-14, 1.107575e-14, 1.108795e-14, 
    1.109961e-14, 1.111917e-14, 1.111595e-14, 1.112456e-14, 1.108763e-14, 
    1.111218e-14, 1.107164e-14, 1.108273e-14, 1.099437e-14, 1.096067e-14, 
    1.094631e-14, 1.093375e-14, 1.090316e-14, 1.092429e-14, 1.091596e-14, 
    1.093577e-14, 1.094835e-14, 1.094213e-14, 1.098051e-14, 1.096559e-14, 
    1.104405e-14, 1.101029e-14, 1.109825e-14, 1.107723e-14, 1.110329e-14, 
    1.108999e-14, 1.111276e-14, 1.109227e-14, 1.112777e-14, 1.113549e-14, 
    1.113021e-14, 1.115048e-14, 1.109113e-14, 1.111394e-14, 1.094196e-14, 
    1.094297e-14, 1.09477e-14, 1.092691e-14, 1.092564e-14, 1.090658e-14, 
    1.092354e-14, 1.093076e-14, 1.094908e-14, 1.095991e-14, 1.09702e-14, 
    1.099282e-14, 1.101805e-14, 1.105329e-14, 1.107859e-14, 1.109553e-14, 
    1.108515e-14, 1.109432e-14, 1.108406e-14, 1.107926e-14, 1.113259e-14, 
    1.110265e-14, 1.114757e-14, 1.114508e-14, 1.112476e-14, 1.114536e-14, 
    1.094368e-14, 1.093785e-14, 1.091756e-14, 1.093344e-14, 1.09045e-14, 
    1.09207e-14, 1.093e-14, 1.09659e-14, 1.097378e-14, 1.098109e-14, 
    1.099551e-14, 1.1014e-14, 1.104642e-14, 1.107459e-14, 1.110029e-14, 
    1.109841e-14, 1.109907e-14, 1.11048e-14, 1.109059e-14, 1.110714e-14, 
    1.110991e-14, 1.110265e-14, 1.114475e-14, 1.113273e-14, 1.114503e-14, 
    1.113721e-14, 1.093974e-14, 1.094957e-14, 1.094426e-14, 1.095424e-14, 
    1.094721e-14, 1.097845e-14, 1.098782e-14, 1.103159e-14, 1.101364e-14, 
    1.104221e-14, 1.101655e-14, 1.102109e-14, 1.104313e-14, 1.101793e-14, 
    1.107303e-14, 1.103568e-14, 1.110503e-14, 1.106776e-14, 1.110736e-14, 
    1.110018e-14, 1.111207e-14, 1.112272e-14, 1.113611e-14, 1.116079e-14, 
    1.115508e-14, 1.117571e-14, 1.096421e-14, 1.097693e-14, 1.097582e-14, 
    1.098914e-14, 1.099898e-14, 1.102031e-14, 1.105448e-14, 1.104164e-14, 
    1.106521e-14, 1.106994e-14, 1.103412e-14, 1.105612e-14, 1.098545e-14, 
    1.099688e-14, 1.099008e-14, 1.096521e-14, 1.104459e-14, 1.100388e-14, 
    1.107901e-14, 1.105699e-14, 1.11212e-14, 1.108928e-14, 1.115193e-14, 
    1.117866e-14, 1.120381e-14, 1.123315e-14, 1.098388e-14, 1.097524e-14, 
    1.099072e-14, 1.101212e-14, 1.103197e-14, 1.105834e-14, 1.106103e-14, 
    1.106597e-14, 1.107875e-14, 1.108949e-14, 1.106752e-14, 1.109218e-14, 
    1.099951e-14, 1.104812e-14, 1.097196e-14, 1.099491e-14, 1.101086e-14, 
    1.100387e-14, 1.104017e-14, 1.104871e-14, 1.108341e-14, 1.106549e-14, 
    1.117206e-14, 1.112496e-14, 1.125548e-14, 1.121906e-14, 1.097222e-14, 
    1.098386e-14, 1.102432e-14, 1.100508e-14, 1.10601e-14, 1.107361e-14, 
    1.108461e-14, 1.109865e-14, 1.110017e-14, 1.110848e-14, 1.109485e-14, 
    1.110794e-14, 1.105839e-14, 1.108054e-14, 1.101971e-14, 1.103453e-14, 
    1.102771e-14, 1.102023e-14, 1.104331e-14, 1.106786e-14, 1.106839e-14, 
    1.107626e-14, 1.10984e-14, 1.106032e-14, 1.117812e-14, 1.110541e-14, 
    1.099655e-14, 1.101893e-14, 1.102214e-14, 1.101347e-14, 1.107226e-14, 
    1.105097e-14, 1.110828e-14, 1.10928e-14, 1.111816e-14, 1.110556e-14, 
    1.110371e-14, 1.108752e-14, 1.107744e-14, 1.105195e-14, 1.103119e-14, 
    1.101473e-14, 1.101856e-14, 1.103664e-14, 1.106936e-14, 1.11003e-14, 
    1.109352e-14, 1.111623e-14, 1.105611e-14, 1.108133e-14, 1.107158e-14, 
    1.109699e-14, 1.104129e-14, 1.10887e-14, 1.102916e-14, 1.103438e-14, 
    1.105055e-14, 1.108303e-14, 1.109023e-14, 1.109789e-14, 1.109317e-14, 
    1.10702e-14, 1.106644e-14, 1.105016e-14, 1.104566e-14, 1.103325e-14, 
    1.102296e-14, 1.103236e-14, 1.104222e-14, 1.107021e-14, 1.109541e-14, 
    1.112287e-14, 1.112959e-14, 1.11616e-14, 1.113553e-14, 1.117852e-14, 
    1.114195e-14, 1.120523e-14, 1.109146e-14, 1.11409e-14, 1.105129e-14, 
    1.106096e-14, 1.107843e-14, 1.111848e-14, 1.109687e-14, 1.112215e-14, 
    1.10663e-14, 1.103726e-14, 1.102975e-14, 1.101573e-14, 1.103007e-14, 
    1.102891e-14, 1.104263e-14, 1.103822e-14, 1.107114e-14, 1.105347e-14, 
    1.110366e-14, 1.112195e-14, 1.117355e-14, 1.120513e-14, 1.123725e-14, 
    1.125141e-14, 1.125572e-14, 1.125752e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.3676e-11, -8.404414e-11, -8.397257e-11, -8.426951e-11, -8.410479e-11, 
    -8.429922e-11, -8.375063e-11, -8.405876e-11, -8.386206e-11, 
    -8.370913e-11, -8.484577e-11, -8.428275e-11, -8.543054e-11, 
    -8.507148e-11, -8.597343e-11, -8.537467e-11, -8.609416e-11, 
    -8.595614e-11, -8.637151e-11, -8.625251e-11, -8.678381e-11, 
    -8.642643e-11, -8.705921e-11, -8.669845e-11, -8.675489e-11, 
    -8.641464e-11, -8.439605e-11, -8.477568e-11, -8.437356e-11, 
    -8.442769e-11, -8.44034e-11, -8.410819e-11, -8.395944e-11, -8.364785e-11, 
    -8.370442e-11, -8.393326e-11, -8.445204e-11, -8.427593e-11, 
    -8.471974e-11, -8.470971e-11, -8.52038e-11, -8.498103e-11, -8.581147e-11, 
    -8.557544e-11, -8.625748e-11, -8.608596e-11, -8.624942e-11, 
    -8.619985e-11, -8.625007e-11, -8.599851e-11, -8.610629e-11, 
    -8.588493e-11, -8.502275e-11, -8.527615e-11, -8.45204e-11, -8.4066e-11, 
    -8.376415e-11, -8.354995e-11, -8.358023e-11, -8.363796e-11, -8.39346e-11, 
    -8.421349e-11, -8.442602e-11, -8.456819e-11, -8.470828e-11, 
    -8.513231e-11, -8.535671e-11, -8.58592e-11, -8.57685e-11, -8.592214e-11, 
    -8.606889e-11, -8.63153e-11, -8.627474e-11, -8.63833e-11, -8.591808e-11, 
    -8.622727e-11, -8.571685e-11, -8.585645e-11, -8.47464e-11, -8.432344e-11, 
    -8.414369e-11, -8.398633e-11, -8.360352e-11, -8.386788e-11, 
    -8.376367e-11, -8.401159e-11, -8.416913e-11, -8.409121e-11, 
    -8.457208e-11, -8.438513e-11, -8.537002e-11, -8.494579e-11, 
    -8.605178e-11, -8.578712e-11, -8.611521e-11, -8.594779e-11, 
    -8.623465e-11, -8.597648e-11, -8.642369e-11, -8.652108e-11, 
    -8.645453e-11, -8.671015e-11, -8.596217e-11, -8.624942e-11, 
    -8.408903e-11, -8.410174e-11, -8.416094e-11, -8.390071e-11, 
    -8.388479e-11, -8.36463e-11, -8.38585e-11, -8.394887e-11, -8.417825e-11, 
    -8.431394e-11, -8.444292e-11, -8.472652e-11, -8.504324e-11, 
    -8.548612e-11, -8.580427e-11, -8.601755e-11, -8.588677e-11, 
    -8.600223e-11, -8.587316e-11, -8.581266e-11, -8.648459e-11, -8.61073e-11, 
    -8.667339e-11, -8.664206e-11, -8.638588e-11, -8.664559e-11, 
    -8.411066e-11, -8.403753e-11, -8.378365e-11, -8.398233e-11, 
    -8.362033e-11, -8.382297e-11, -8.393949e-11, -8.438905e-11, 
    -8.448781e-11, -8.457941e-11, -8.476029e-11, -8.499243e-11, 
    -8.539967e-11, -8.575398e-11, -8.607743e-11, -8.605373e-11, 
    -8.606207e-11, -8.613433e-11, -8.595535e-11, -8.616372e-11, 
    -8.619869e-11, -8.610725e-11, -8.663787e-11, -8.648628e-11, -8.66414e-11, 
    -8.654269e-11, -8.40613e-11, -8.418435e-11, -8.411786e-11, -8.424289e-11, 
    -8.415481e-11, -8.454648e-11, -8.466391e-11, -8.521338e-11, 
    -8.498786e-11, -8.534676e-11, -8.502432e-11, -8.508146e-11, 
    -8.535848e-11, -8.504174e-11, -8.573445e-11, -8.526483e-11, 
    -8.613714e-11, -8.566819e-11, -8.616653e-11, -8.607603e-11, 
    -8.622586e-11, -8.636006e-11, -8.652887e-11, -8.684038e-11, 
    -8.676825e-11, -8.702875e-11, -8.436778e-11, -8.452738e-11, 
    -8.451332e-11, -8.468034e-11, -8.480386e-11, -8.507157e-11, 
    -8.550094e-11, -8.533948e-11, -8.563589e-11, -8.56954e-11, -8.524507e-11, 
    -8.552158e-11, -8.463419e-11, -8.477757e-11, -8.469219e-11, 
    -8.438037e-11, -8.53767e-11, -8.486539e-11, -8.580953e-11, -8.553255e-11, 
    -8.634093e-11, -8.593892e-11, -8.672854e-11, -8.706612e-11, 
    -8.738379e-11, -8.775508e-11, -8.461448e-11, -8.450603e-11, -8.47002e-11, 
    -8.496884e-11, -8.521808e-11, -8.554945e-11, -8.558335e-11, 
    -8.564543e-11, -8.580622e-11, -8.594141e-11, -8.566506e-11, -8.59753e-11, 
    -8.481083e-11, -8.542107e-11, -8.446504e-11, -8.475293e-11, -8.4953e-11, 
    -8.486523e-11, -8.532102e-11, -8.542845e-11, -8.586498e-11, 
    -8.563932e-11, -8.698281e-11, -8.638842e-11, -8.803776e-11, 
    -8.757684e-11, -8.446814e-11, -8.46141e-11, -8.512208e-11, -8.488038e-11, 
    -8.557156e-11, -8.57417e-11, -8.588e-11, -8.60568e-11, -8.607588e-11, 
    -8.618064e-11, -8.600898e-11, -8.617385e-11, -8.555015e-11, 
    -8.582887e-11, -8.5064e-11, -8.525017e-11, -8.516452e-11, -8.507058e-11, 
    -8.536052e-11, -8.566941e-11, -8.567599e-11, -8.577505e-11, 
    -8.605419e-11, -8.557436e-11, -8.705955e-11, -8.614236e-11, 
    -8.477325e-11, -8.50544e-11, -8.509454e-11, -8.498564e-11, -8.572464e-11, 
    -8.545688e-11, -8.617808e-11, -8.598317e-11, -8.630253e-11, 
    -8.614383e-11, -8.612049e-11, -8.591666e-11, -8.578976e-11, 
    -8.546915e-11, -8.520829e-11, -8.500143e-11, -8.504953e-11, 
    -8.527676e-11, -8.56883e-11, -8.607762e-11, -8.599234e-11, -8.627826e-11, 
    -8.552144e-11, -8.58388e-11, -8.571614e-11, -8.603596e-11, -8.533519e-11, 
    -8.593197e-11, -8.518265e-11, -8.524834e-11, -8.545156e-11, 
    -8.586033e-11, -8.595075e-11, -8.604732e-11, -8.598772e-11, 
    -8.569875e-11, -8.56514e-11, -8.544662e-11, -8.539008e-11, -8.523404e-11, 
    -8.510486e-11, -8.522289e-11, -8.534685e-11, -8.569886e-11, -8.60161e-11, 
    -8.636197e-11, -8.644661e-11, -8.685075e-11, -8.652178e-11, 
    -8.706466e-11, -8.660313e-11, -8.740205e-11, -8.596653e-11, 
    -8.658953e-11, -8.546081e-11, -8.55824e-11, -8.580235e-11, -8.63068e-11, 
    -8.603445e-11, -8.635295e-11, -8.564954e-11, -8.528461e-11, 
    -8.519017e-11, -8.501401e-11, -8.51942e-11, -8.517954e-11, -8.535198e-11, 
    -8.529656e-11, -8.571055e-11, -8.548818e-11, -8.61199e-11, -8.635043e-11, 
    -8.700145e-11, -8.740056e-11, -8.78068e-11, -8.798615e-11, -8.804073e-11, 
    -8.806356e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -2.01674e-12, -2.025611e-12, -2.023886e-12, -2.031042e-12, -2.027072e-12, 
    -2.031758e-12, -2.018538e-12, -2.025963e-12, -2.021223e-12, 
    -2.017538e-12, -2.044927e-12, -2.031361e-12, -2.059018e-12, 
    -2.050366e-12, -2.0721e-12, -2.057672e-12, -2.075009e-12, -2.071683e-12, 
    -2.081692e-12, -2.078825e-12, -2.091627e-12, -2.083015e-12, 
    -2.098263e-12, -2.08957e-12, -2.09093e-12, -2.082731e-12, -2.034091e-12, 
    -2.043238e-12, -2.033549e-12, -2.034853e-12, -2.034268e-12, 
    -2.027154e-12, -2.02357e-12, -2.016062e-12, -2.017425e-12, -2.022939e-12, 
    -2.03544e-12, -2.031196e-12, -2.04189e-12, -2.041649e-12, -2.053555e-12, 
    -2.048187e-12, -2.068197e-12, -2.06251e-12, -2.078944e-12, -2.074811e-12, 
    -2.07875e-12, -2.077556e-12, -2.078766e-12, -2.072704e-12, -2.075301e-12, 
    -2.069967e-12, -2.049192e-12, -2.055298e-12, -2.037087e-12, 
    -2.026138e-12, -2.018864e-12, -2.013703e-12, -2.014432e-12, 
    -2.015823e-12, -2.022971e-12, -2.029692e-12, -2.034813e-12, 
    -2.038239e-12, -2.041614e-12, -2.051832e-12, -2.057239e-12, 
    -2.069347e-12, -2.067162e-12, -2.070864e-12, -2.0744e-12, -2.080337e-12, 
    -2.07936e-12, -2.081976e-12, -2.070766e-12, -2.078216e-12, -2.065917e-12, 
    -2.069281e-12, -2.042533e-12, -2.032341e-12, -2.02801e-12, -2.024218e-12, 
    -2.014993e-12, -2.021364e-12, -2.018853e-12, -2.024827e-12, 
    -2.028623e-12, -2.026745e-12, -2.038332e-12, -2.033828e-12, -2.05756e-12, 
    -2.047338e-12, -2.073988e-12, -2.06761e-12, -2.075516e-12, -2.071482e-12, 
    -2.078394e-12, -2.072173e-12, -2.082949e-12, -2.085296e-12, 
    -2.083692e-12, -2.089852e-12, -2.071828e-12, -2.07875e-12, -2.026693e-12, 
    -2.026999e-12, -2.028425e-12, -2.022155e-12, -2.021771e-12, 
    -2.016025e-12, -2.021138e-12, -2.023315e-12, -2.028843e-12, 
    -2.032112e-12, -2.03522e-12, -2.042054e-12, -2.049686e-12, -2.060357e-12, 
    -2.068024e-12, -2.073163e-12, -2.070012e-12, -2.072794e-12, 
    -2.069684e-12, -2.068226e-12, -2.084417e-12, -2.075326e-12, 
    -2.088966e-12, -2.088211e-12, -2.082038e-12, -2.088296e-12, 
    -2.027214e-12, -2.025452e-12, -2.019334e-12, -2.024122e-12, 
    -2.015398e-12, -2.020282e-12, -2.023089e-12, -2.033922e-12, 
    -2.036302e-12, -2.038509e-12, -2.042868e-12, -2.048461e-12, 
    -2.058274e-12, -2.066812e-12, -2.074606e-12, -2.074035e-12, 
    -2.074236e-12, -2.075977e-12, -2.071664e-12, -2.076685e-12, 
    -2.077528e-12, -2.075324e-12, -2.08811e-12, -2.084457e-12, -2.088195e-12, 
    -2.085817e-12, -2.026025e-12, -2.028989e-12, -2.027387e-12, -2.0304e-12, 
    -2.028278e-12, -2.037715e-12, -2.040545e-12, -2.053785e-12, 
    -2.048351e-12, -2.056999e-12, -2.04923e-12, -2.050606e-12, -2.057282e-12, 
    -2.04965e-12, -2.066341e-12, -2.055025e-12, -2.076045e-12, -2.064745e-12, 
    -2.076753e-12, -2.074572e-12, -2.078182e-12, -2.081416e-12, 
    -2.085484e-12, -2.09299e-12, -2.091252e-12, -2.097529e-12, -2.033409e-12, 
    -2.037255e-12, -2.036916e-12, -2.040941e-12, -2.043917e-12, 
    -2.050368e-12, -2.060715e-12, -2.056824e-12, -2.063966e-12, -2.0654e-12, 
    -2.054549e-12, -2.061212e-12, -2.039829e-12, -2.043284e-12, 
    -2.041227e-12, -2.033713e-12, -2.057721e-12, -2.0454e-12, -2.068151e-12, 
    -2.061476e-12, -2.080955e-12, -2.071268e-12, -2.090295e-12, -2.09843e-12, 
    -2.106084e-12, -2.115031e-12, -2.039354e-12, -2.036741e-12, -2.04142e-12, 
    -2.047893e-12, -2.053899e-12, -2.061883e-12, -2.0627e-12, -2.064196e-12, 
    -2.068071e-12, -2.071328e-12, -2.064669e-12, -2.072145e-12, 
    -2.044086e-12, -2.05879e-12, -2.035753e-12, -2.04269e-12, -2.047511e-12, 
    -2.045396e-12, -2.056379e-12, -2.058968e-12, -2.069487e-12, 
    -2.064049e-12, -2.096422e-12, -2.082099e-12, -2.121842e-12, 
    -2.110736e-12, -2.035828e-12, -2.039345e-12, -2.051585e-12, 
    -2.045761e-12, -2.062416e-12, -2.066516e-12, -2.069848e-12, 
    -2.074109e-12, -2.074568e-12, -2.077093e-12, -2.072956e-12, 
    -2.076929e-12, -2.0619e-12, -2.068616e-12, -2.050186e-12, -2.054672e-12, 
    -2.052608e-12, -2.050344e-12, -2.057331e-12, -2.064774e-12, 
    -2.064933e-12, -2.06732e-12, -2.074046e-12, -2.062484e-12, -2.098271e-12, 
    -2.07617e-12, -2.04318e-12, -2.049955e-12, -2.050922e-12, -2.048298e-12, 
    -2.066105e-12, -2.059653e-12, -2.077031e-12, -2.072334e-12, -2.08003e-12, 
    -2.076206e-12, -2.075643e-12, -2.070732e-12, -2.067674e-12, 
    -2.059949e-12, -2.053663e-12, -2.048678e-12, -2.049837e-12, 
    -2.055313e-12, -2.065229e-12, -2.07461e-12, -2.072555e-12, -2.079445e-12, 
    -2.061209e-12, -2.068856e-12, -2.0659e-12, -2.073606e-12, -2.05672e-12, 
    -2.071101e-12, -2.053045e-12, -2.054628e-12, -2.059525e-12, 
    -2.069375e-12, -2.071553e-12, -2.07388e-12, -2.072444e-12, -2.065481e-12, 
    -2.06434e-12, -2.059406e-12, -2.058043e-12, -2.054283e-12, -2.05117e-12, 
    -2.054015e-12, -2.057001e-12, -2.065484e-12, -2.073128e-12, 
    -2.081462e-12, -2.083502e-12, -2.09324e-12, -2.085313e-12, -2.098394e-12, 
    -2.087273e-12, -2.106524e-12, -2.071934e-12, -2.086946e-12, 
    -2.059747e-12, -2.062678e-12, -2.067978e-12, -2.080133e-12, -2.07357e-12, 
    -2.081245e-12, -2.064295e-12, -2.055502e-12, -2.053226e-12, 
    -2.048981e-12, -2.053323e-12, -2.05297e-12, -2.057125e-12, -2.05579e-12, 
    -2.065765e-12, -2.060407e-12, -2.075629e-12, -2.081184e-12, 
    -2.096871e-12, -2.106488e-12, -2.116277e-12, -2.120598e-12, 
    -2.121914e-12, -2.122464e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.543816e-15, 3.553372e-15, 3.551516e-15, 3.559217e-15, 3.554947e-15, 
    3.559987e-15, 3.545755e-15, 3.55375e-15, 3.548648e-15, 3.544678e-15, 
    3.574139e-15, 3.55956e-15, 3.589269e-15, 3.579988e-15, 3.603286e-15, 
    3.587824e-15, 3.606401e-15, 3.602843e-15, 3.613555e-15, 3.610488e-15, 
    3.624169e-15, 3.614971e-15, 3.631257e-15, 3.621975e-15, 3.623426e-15, 
    3.614667e-15, 3.562499e-15, 3.572324e-15, 3.561916e-15, 3.563318e-15, 
    3.562689e-15, 3.555034e-15, 3.551172e-15, 3.543087e-15, 3.544556e-15, 
    3.550495e-15, 3.563948e-15, 3.559385e-15, 3.570886e-15, 3.570626e-15, 
    3.583411e-15, 3.577649e-15, 3.599109e-15, 3.593017e-15, 3.610616e-15, 
    3.606192e-15, 3.610408e-15, 3.60913e-15, 3.610425e-15, 3.603936e-15, 
    3.606716e-15, 3.601006e-15, 3.578727e-15, 3.58528e-15, 3.565721e-15, 
    3.553935e-15, 3.546106e-15, 3.540544e-15, 3.54133e-15, 3.542829e-15, 
    3.550529e-15, 3.557766e-15, 3.563277e-15, 3.56696e-15, 3.570589e-15, 
    3.581556e-15, 3.587361e-15, 3.600339e-15, 3.598001e-15, 3.601964e-15, 
    3.605752e-15, 3.612106e-15, 3.61106e-15, 3.613858e-15, 3.601861e-15, 
    3.609835e-15, 3.596668e-15, 3.600271e-15, 3.571566e-15, 3.560617e-15, 
    3.555951e-15, 3.551872e-15, 3.541935e-15, 3.548798e-15, 3.546093e-15, 
    3.552529e-15, 3.556616e-15, 3.554595e-15, 3.567061e-15, 3.562217e-15, 
    3.587705e-15, 3.576735e-15, 3.605311e-15, 3.598481e-15, 3.606947e-15, 
    3.602628e-15, 3.610026e-15, 3.603369e-15, 3.614899e-15, 3.617407e-15, 
    3.615693e-15, 3.622278e-15, 3.602999e-15, 3.610407e-15, 3.554538e-15, 
    3.554868e-15, 3.556404e-15, 3.54965e-15, 3.549237e-15, 3.543046e-15, 
    3.548556e-15, 3.5509e-15, 3.556854e-15, 3.560371e-15, 3.563714e-15, 
    3.57106e-15, 3.579256e-15, 3.590707e-15, 3.598924e-15, 3.604428e-15, 
    3.601054e-15, 3.604033e-15, 3.600702e-15, 3.599141e-15, 3.616467e-15, 
    3.606742e-15, 3.621331e-15, 3.620525e-15, 3.613924e-15, 3.620616e-15, 
    3.555099e-15, 3.553203e-15, 3.546612e-15, 3.551771e-15, 3.542372e-15, 
    3.547633e-15, 3.550655e-15, 3.562316e-15, 3.564878e-15, 3.56725e-15, 
    3.571935e-15, 3.577943e-15, 3.588473e-15, 3.597624e-15, 3.605973e-15, 
    3.605362e-15, 3.605577e-15, 3.60744e-15, 3.602823e-15, 3.608198e-15, 
    3.609099e-15, 3.606742e-15, 3.620417e-15, 3.616512e-15, 3.620508e-15, 
    3.617966e-15, 3.553819e-15, 3.557011e-15, 3.555286e-15, 3.558528e-15, 
    3.556244e-15, 3.566395e-15, 3.569436e-15, 3.583655e-15, 3.577825e-15, 
    3.587105e-15, 3.578769e-15, 3.580246e-15, 3.587403e-15, 3.57922e-15, 
    3.597118e-15, 3.584984e-15, 3.607512e-15, 3.595406e-15, 3.608271e-15, 
    3.605937e-15, 3.609801e-15, 3.613259e-15, 3.61761e-15, 3.625628e-15, 
    3.623773e-15, 3.630476e-15, 3.561767e-15, 3.565901e-15, 3.565539e-15, 
    3.569865e-15, 3.573063e-15, 3.579992e-15, 3.591091e-15, 3.586919e-15, 
    3.594579e-15, 3.596113e-15, 3.584479e-15, 3.591623e-15, 3.568668e-15, 
    3.572379e-15, 3.570171e-15, 3.562092e-15, 3.587878e-15, 3.574653e-15, 
    3.599059e-15, 3.591908e-15, 3.612766e-15, 3.602396e-15, 3.62275e-15, 
    3.631432e-15, 3.639603e-15, 3.649132e-15, 3.568158e-15, 3.56535e-15, 
    3.57038e-15, 3.577331e-15, 3.58378e-15, 3.592344e-15, 3.593221e-15, 
    3.594824e-15, 3.598975e-15, 3.602464e-15, 3.595329e-15, 3.603338e-15, 
    3.573236e-15, 3.589026e-15, 3.564286e-15, 3.571741e-15, 3.576922e-15, 
    3.574651e-15, 3.586443e-15, 3.589219e-15, 3.600489e-15, 3.594667e-15, 
    3.629288e-15, 3.613987e-15, 3.656387e-15, 3.644558e-15, 3.564368e-15, 
    3.56815e-15, 3.581296e-15, 3.575044e-15, 3.592917e-15, 3.597308e-15, 
    3.600879e-15, 3.605439e-15, 3.605933e-15, 3.608634e-15, 3.604207e-15, 
    3.608459e-15, 3.592362e-15, 3.599559e-15, 3.579796e-15, 3.58461e-15, 
    3.582396e-15, 3.579967e-15, 3.587464e-15, 3.595439e-15, 3.595612e-15, 
    3.598168e-15, 3.605361e-15, 3.592989e-15, 3.631256e-15, 3.607637e-15, 
    3.572271e-15, 3.579543e-15, 3.580585e-15, 3.577768e-15, 3.596867e-15, 
    3.589953e-15, 3.608568e-15, 3.603541e-15, 3.611777e-15, 3.607685e-15, 
    3.607083e-15, 3.601825e-15, 3.598549e-15, 3.590269e-15, 3.583527e-15, 
    3.578178e-15, 3.579422e-15, 3.585297e-15, 3.595927e-15, 3.605976e-15, 
    3.603775e-15, 3.611152e-15, 3.591622e-15, 3.599814e-15, 3.596647e-15, 
    3.604903e-15, 3.586808e-15, 3.60221e-15, 3.582865e-15, 3.584564e-15, 
    3.589815e-15, 3.600367e-15, 3.602705e-15, 3.605195e-15, 3.603659e-15, 
    3.596197e-15, 3.594978e-15, 3.589689e-15, 3.588226e-15, 3.584194e-15, 
    3.580853e-15, 3.583905e-15, 3.587108e-15, 3.596202e-15, 3.604389e-15, 
    3.613308e-15, 3.61549e-15, 3.625889e-15, 3.617421e-15, 3.631386e-15, 
    3.619508e-15, 3.640063e-15, 3.603106e-15, 3.619165e-15, 3.590056e-15, 
    3.593197e-15, 3.598871e-15, 3.611883e-15, 3.604864e-15, 3.613073e-15, 
    3.59493e-15, 3.585498e-15, 3.583059e-15, 3.578502e-15, 3.583164e-15, 
    3.582785e-15, 3.587243e-15, 3.585811e-15, 3.596504e-15, 3.590762e-15, 
    3.607067e-15, 3.613009e-15, 3.629772e-15, 3.64003e-15, 3.650464e-15, 
    3.655065e-15, 3.656465e-15, 3.65705e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.760421e-09, -8.798932e-09, -8.791446e-09, -8.822508e-09, -8.805277e-09, 
    -8.825616e-09, -8.768228e-09, -8.800462e-09, -8.779884e-09, 
    -8.763887e-09, -8.882789e-09, -8.823894e-09, -8.94396e-09, -8.9064e-09, 
    -9.00075e-09, -8.938116e-09, -9.013379e-09, -8.998942e-09, -9.042392e-09, 
    -9.029944e-09, -9.085521e-09, -9.048136e-09, -9.114328e-09, 
    -9.076592e-09, -9.082496e-09, -9.046904e-09, -8.835745e-09, 
    -8.875457e-09, -8.833392e-09, -8.839055e-09, -8.836514e-09, 
    -8.805633e-09, -8.790071e-09, -8.757477e-09, -8.763394e-09, 
    -8.787334e-09, -8.841601e-09, -8.823179e-09, -8.869605e-09, 
    -8.868557e-09, -8.920242e-09, -8.896938e-09, -8.983807e-09, 
    -8.959118e-09, -9.030463e-09, -9.012521e-09, -9.029621e-09, 
    -9.024435e-09, -9.029688e-09, -9.003374e-09, -9.014649e-09, 
    -8.991493e-09, -8.901303e-09, -8.92781e-09, -8.848754e-09, -8.801218e-09, 
    -8.769642e-09, -8.747236e-09, -8.750404e-09, -8.756443e-09, 
    -8.787473e-09, -8.816648e-09, -8.838881e-09, -8.853752e-09, 
    -8.868406e-09, -8.912764e-09, -8.936238e-09, -8.988801e-09, 
    -8.979314e-09, -8.995385e-09, -9.010736e-09, -9.036511e-09, 
    -9.032268e-09, -9.043625e-09, -8.99496e-09, -9.027303e-09, -8.973911e-09, 
    -8.988514e-09, -8.872394e-09, -8.828149e-09, -8.809346e-09, 
    -8.792885e-09, -8.752839e-09, -8.780495e-09, -8.769592e-09, 
    -8.795527e-09, -8.812007e-09, -8.803856e-09, -8.854159e-09, 
    -8.834603e-09, -8.937629e-09, -8.893253e-09, -9.008946e-09, 
    -8.981261e-09, -9.015581e-09, -8.998068e-09, -9.028076e-09, 
    -9.001069e-09, -9.04785e-09, -9.058038e-09, -9.051076e-09, -9.077816e-09, 
    -8.999572e-09, -9.029621e-09, -8.803628e-09, -8.804958e-09, -8.81115e-09, 
    -8.783928e-09, -8.782263e-09, -8.757315e-09, -8.779513e-09, 
    -8.788966e-09, -8.812962e-09, -8.827156e-09, -8.840649e-09, 
    -8.870315e-09, -8.903447e-09, -8.949774e-09, -8.983056e-09, 
    -9.005365e-09, -8.991685e-09, -9.003763e-09, -8.990262e-09, 
    -8.983933e-09, -9.05422e-09, -9.014753e-09, -9.07397e-09, -9.070693e-09, 
    -9.043895e-09, -9.071062e-09, -8.805891e-09, -8.798241e-09, 
    -8.771682e-09, -8.792467e-09, -8.754598e-09, -8.775796e-09, 
    -8.787985e-09, -8.835013e-09, -8.845344e-09, -8.854925e-09, 
    -8.873847e-09, -8.898131e-09, -8.940731e-09, -8.977795e-09, 
    -9.011629e-09, -9.00915e-09, -9.010023e-09, -9.017581e-09, -8.998859e-09, 
    -9.020655e-09, -9.024314e-09, -9.014749e-09, -9.070254e-09, 
    -9.054396e-09, -9.070623e-09, -9.060298e-09, -8.800727e-09, -8.8136e-09, 
    -8.806644e-09, -8.819724e-09, -8.810509e-09, -8.851481e-09, 
    -8.863766e-09, -8.921243e-09, -8.897653e-09, -8.935196e-09, 
    -8.901467e-09, -8.907444e-09, -8.936422e-09, -8.903289e-09, 
    -8.975752e-09, -8.926627e-09, -9.017875e-09, -8.96882e-09, -9.020949e-09, 
    -9.011483e-09, -9.027156e-09, -9.041194e-09, -9.058853e-09, 
    -9.091439e-09, -9.083893e-09, -9.111143e-09, -8.832788e-09, 
    -8.849483e-09, -8.848012e-09, -8.865483e-09, -8.878405e-09, 
    -8.906409e-09, -8.951325e-09, -8.934435e-09, -8.965442e-09, 
    -8.971667e-09, -8.924559e-09, -8.953483e-09, -8.860656e-09, 
    -8.875655e-09, -8.866724e-09, -8.834105e-09, -8.938328e-09, 
    -8.884841e-09, -8.983606e-09, -8.954632e-09, -9.039193e-09, -8.99714e-09, 
    -9.079739e-09, -9.115052e-09, -9.148282e-09, -9.18712e-09, -8.858594e-09, 
    -8.84725e-09, -8.867561e-09, -8.895664e-09, -8.921736e-09, -8.956399e-09, 
    -8.959945e-09, -8.966439e-09, -8.983259e-09, -8.997401e-09, 
    -8.968493e-09, -9.000946e-09, -8.879135e-09, -8.94297e-09, -8.842962e-09, 
    -8.873078e-09, -8.894007e-09, -8.884825e-09, -8.932504e-09, 
    -8.943742e-09, -8.989406e-09, -8.9658e-09, -9.106337e-09, -9.04416e-09, 
    -9.216689e-09, -9.168476e-09, -8.843287e-09, -8.858555e-09, 
    -8.911693e-09, -8.88641e-09, -8.958712e-09, -8.976509e-09, -8.990977e-09, 
    -9.009471e-09, -9.011467e-09, -9.022425e-09, -9.004469e-09, 
    -9.021716e-09, -8.956473e-09, -8.985628e-09, -8.905618e-09, 
    -8.925093e-09, -8.916134e-09, -8.906307e-09, -8.936635e-09, 
    -8.968948e-09, -8.969637e-09, -8.979998e-09, -9.009198e-09, 
    -8.959005e-09, -9.114364e-09, -9.018422e-09, -8.875204e-09, 
    -8.904613e-09, -8.908812e-09, -8.897421e-09, -8.974725e-09, 
    -8.946715e-09, -9.022158e-09, -9.001768e-09, -9.035176e-09, 
    -9.018575e-09, -9.016133e-09, -8.994811e-09, -8.981537e-09, -8.948e-09, 
    -8.920712e-09, -8.899073e-09, -8.904104e-09, -8.927874e-09, 
    -8.970924e-09, -9.011649e-09, -9.002728e-09, -9.032637e-09, -8.95347e-09, 
    -8.986667e-09, -8.973837e-09, -9.007291e-09, -8.933986e-09, 
    -8.996413e-09, -8.918029e-09, -8.924902e-09, -8.946159e-09, -8.98892e-09, 
    -8.998378e-09, -9.008479e-09, -9.002246e-09, -8.972017e-09, 
    -8.967064e-09, -8.945642e-09, -8.939728e-09, -8.923405e-09, 
    -8.909891e-09, -8.922239e-09, -8.935205e-09, -8.972029e-09, 
    -9.005214e-09, -9.041394e-09, -9.050248e-09, -9.092523e-09, 
    -9.058111e-09, -9.114899e-09, -9.066621e-09, -9.150191e-09, 
    -9.000029e-09, -9.065198e-09, -8.947127e-09, -8.959846e-09, 
    -8.982854e-09, -9.035623e-09, -9.007134e-09, -9.040451e-09, -8.96687e-09, 
    -8.928695e-09, -8.918817e-09, -8.900388e-09, -8.919238e-09, 
    -8.917705e-09, -8.935742e-09, -8.929946e-09, -8.973251e-09, -8.94999e-09, 
    -9.016072e-09, -9.040187e-09, -9.108287e-09, -9.150035e-09, 
    -9.192529e-09, -9.21129e-09, -9.217e-09, -9.219387e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.039521e-10, -1.044092e-10, -1.043203e-10, -1.046891e-10, -1.044845e-10, 
    -1.04726e-10, -1.040447e-10, -1.044274e-10, -1.041831e-10, -1.039932e-10, 
    -1.054047e-10, -1.047055e-10, -1.061308e-10, -1.056849e-10, -1.06805e-10, 
    -1.060614e-10, -1.069549e-10, -1.067835e-10, -1.072993e-10, 
    -1.071516e-10, -1.078113e-10, -1.073675e-10, -1.081533e-10, 
    -1.077053e-10, -1.077754e-10, -1.073529e-10, -1.048462e-10, 
    -1.053176e-10, -1.048183e-10, -1.048855e-10, -1.048553e-10, 
    -1.044887e-10, -1.04304e-10, -1.039171e-10, -1.039873e-10, -1.042715e-10, 
    -1.049157e-10, -1.04697e-10, -1.052482e-10, -1.052357e-10, -1.058493e-10, 
    -1.055726e-10, -1.066039e-10, -1.063108e-10, -1.071577e-10, 
    -1.069447e-10, -1.071477e-10, -1.070862e-10, -1.071485e-10, 
    -1.068361e-10, -1.0697e-10, -1.066951e-10, -1.056244e-10, -1.059391e-10, 
    -1.050006e-10, -1.044363e-10, -1.040615e-10, -1.037955e-10, 
    -1.038331e-10, -1.039048e-10, -1.042732e-10, -1.046195e-10, 
    -1.048834e-10, -1.0506e-10, -1.052339e-10, -1.057605e-10, -1.060391e-10, 
    -1.066631e-10, -1.065505e-10, -1.067413e-10, -1.069235e-10, 
    -1.072295e-10, -1.071792e-10, -1.07314e-10, -1.067362e-10, -1.071202e-10, 
    -1.064864e-10, -1.066597e-10, -1.052813e-10, -1.04756e-10, -1.045328e-10, 
    -1.043374e-10, -1.038621e-10, -1.041903e-10, -1.040609e-10, 
    -1.043688e-10, -1.045644e-10, -1.044677e-10, -1.050648e-10, 
    -1.048326e-10, -1.060557e-10, -1.055289e-10, -1.069023e-10, 
    -1.065736e-10, -1.06981e-10, -1.067731e-10, -1.071294e-10, -1.068088e-10, 
    -1.073641e-10, -1.074851e-10, -1.074024e-10, -1.077199e-10, -1.06791e-10, 
    -1.071477e-10, -1.04465e-10, -1.044807e-10, -1.045542e-10, -1.042311e-10, 
    -1.042113e-10, -1.039152e-10, -1.041787e-10, -1.042909e-10, 
    -1.045758e-10, -1.047442e-10, -1.049044e-10, -1.052566e-10, 
    -1.056499e-10, -1.061998e-10, -1.065949e-10, -1.068598e-10, 
    -1.066974e-10, -1.068408e-10, -1.066805e-10, -1.066053e-10, 
    -1.074398e-10, -1.069712e-10, -1.076742e-10, -1.076353e-10, 
    -1.073172e-10, -1.076397e-10, -1.044918e-10, -1.04401e-10, -1.040857e-10, 
    -1.043325e-10, -1.038829e-10, -1.041346e-10, -1.042793e-10, 
    -1.048375e-10, -1.049601e-10, -1.050739e-10, -1.052985e-10, 
    -1.055868e-10, -1.060925e-10, -1.065325e-10, -1.069341e-10, 
    -1.069047e-10, -1.069151e-10, -1.070048e-10, -1.067825e-10, 
    -1.070413e-10, -1.070847e-10, -1.069712e-10, -1.076301e-10, 
    -1.074418e-10, -1.076345e-10, -1.075119e-10, -1.044305e-10, 
    -1.045833e-10, -1.045007e-10, -1.04656e-10, -1.045466e-10, -1.05033e-10, 
    -1.051788e-10, -1.058611e-10, -1.055811e-10, -1.060268e-10, 
    -1.056264e-10, -1.056973e-10, -1.060413e-10, -1.05648e-10, -1.065082e-10, 
    -1.05925e-10, -1.070083e-10, -1.064259e-10, -1.070448e-10, -1.069324e-10, 
    -1.071185e-10, -1.072851e-10, -1.074947e-10, -1.078816e-10, -1.07792e-10, 
    -1.081155e-10, -1.048111e-10, -1.050093e-10, -1.049918e-10, 
    -1.051992e-10, -1.053526e-10, -1.05685e-10, -1.062182e-10, -1.060177e-10, 
    -1.063858e-10, -1.064597e-10, -1.059005e-10, -1.062439e-10, 
    -1.051419e-10, -1.0532e-10, -1.052139e-10, -1.048267e-10, -1.06064e-10, 
    -1.05429e-10, -1.066015e-10, -1.062575e-10, -1.072614e-10, -1.067621e-10, 
    -1.077427e-10, -1.081619e-10, -1.085564e-10, -1.090175e-10, 
    -1.051174e-10, -1.049828e-10, -1.052239e-10, -1.055575e-10, -1.05867e-10, 
    -1.062785e-10, -1.063206e-10, -1.063977e-10, -1.065973e-10, 
    -1.067652e-10, -1.064221e-10, -1.068073e-10, -1.053613e-10, 
    -1.061191e-10, -1.049319e-10, -1.052894e-10, -1.055378e-10, 
    -1.054288e-10, -1.059948e-10, -1.061282e-10, -1.066703e-10, 
    -1.063901e-10, -1.080585e-10, -1.073203e-10, -1.093685e-10, 
    -1.087962e-10, -1.049357e-10, -1.05117e-10, -1.057478e-10, -1.054476e-10, 
    -1.063059e-10, -1.065172e-10, -1.06689e-10, -1.069085e-10, -1.069322e-10, 
    -1.070623e-10, -1.068491e-10, -1.070539e-10, -1.062794e-10, 
    -1.066255e-10, -1.056757e-10, -1.059068e-10, -1.058005e-10, 
    -1.056838e-10, -1.060439e-10, -1.064275e-10, -1.064356e-10, 
    -1.065586e-10, -1.069053e-10, -1.063094e-10, -1.081538e-10, 
    -1.070148e-10, -1.053146e-10, -1.056637e-10, -1.057136e-10, 
    -1.055783e-10, -1.06496e-10, -1.061635e-10, -1.070591e-10, -1.068171e-10, 
    -1.072137e-10, -1.070166e-10, -1.069876e-10, -1.067345e-10, 
    -1.065769e-10, -1.061788e-10, -1.058548e-10, -1.055979e-10, 
    -1.056577e-10, -1.059399e-10, -1.064509e-10, -1.069344e-10, 
    -1.068285e-10, -1.071835e-10, -1.062437e-10, -1.066378e-10, 
    -1.064855e-10, -1.068826e-10, -1.060124e-10, -1.067535e-10, -1.05823e-10, 
    -1.059046e-10, -1.061569e-10, -1.066645e-10, -1.067768e-10, 
    -1.068967e-10, -1.068227e-10, -1.064639e-10, -1.064051e-10, 
    -1.061508e-10, -1.060806e-10, -1.058868e-10, -1.057264e-10, -1.05873e-10, 
    -1.060269e-10, -1.06464e-10, -1.06858e-10, -1.072875e-10, -1.073926e-10, 
    -1.078945e-10, -1.074859e-10, -1.081601e-10, -1.07587e-10, -1.085791e-10, 
    -1.067964e-10, -1.075701e-10, -1.061684e-10, -1.063194e-10, 
    -1.065925e-10, -1.07219e-10, -1.068808e-10, -1.072763e-10, -1.064028e-10, 
    -1.059496e-10, -1.058323e-10, -1.056136e-10, -1.058373e-10, 
    -1.058191e-10, -1.060333e-10, -1.059644e-10, -1.064785e-10, 
    -1.062024e-10, -1.069869e-10, -1.072732e-10, -1.080816e-10, 
    -1.085772e-10, -1.090817e-10, -1.093045e-10, -1.093722e-10, -1.094006e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.622351e-12, -8.660286e-12, -8.652911e-12, -8.683509e-12, -8.666535e-12, 
    -8.686571e-12, -8.630041e-12, -8.661793e-12, -8.641523e-12, 
    -8.625765e-12, -8.742889e-12, -8.684874e-12, -8.803147e-12, 
    -8.766148e-12, -8.859089e-12, -8.79739e-12, -8.871529e-12, -8.857307e-12, 
    -8.900108e-12, -8.887847e-12, -8.942594e-12, -8.905768e-12, 
    -8.970972e-12, -8.933799e-12, -8.939615e-12, -8.904553e-12, 
    -8.696548e-12, -8.735667e-12, -8.69423e-12, -8.699809e-12, -8.697306e-12, 
    -8.666887e-12, -8.651558e-12, -8.619451e-12, -8.625279e-12, -8.64886e-12, 
    -8.702318e-12, -8.684171e-12, -8.729902e-12, -8.72887e-12, -8.779783e-12, 
    -8.756828e-12, -8.842399e-12, -8.818078e-12, -8.888359e-12, 
    -8.870684e-12, -8.887529e-12, -8.882421e-12, -8.887595e-12, 
    -8.861674e-12, -8.872779e-12, -8.849969e-12, -8.761127e-12, 
    -8.787237e-12, -8.709363e-12, -8.662539e-12, -8.631434e-12, 
    -8.609363e-12, -8.612483e-12, -8.618431e-12, -8.648998e-12, 
    -8.677736e-12, -8.699637e-12, -8.714287e-12, -8.728721e-12, 
    -8.772416e-12, -8.79554e-12, -8.847318e-12, -8.837973e-12, -8.853803e-12, 
    -8.868926e-12, -8.894316e-12, -8.890137e-12, -8.901323e-12, 
    -8.853385e-12, -8.885245e-12, -8.83265e-12, -8.847035e-12, -8.73265e-12, 
    -8.689066e-12, -8.670544e-12, -8.654329e-12, -8.614882e-12, 
    -8.642123e-12, -8.631385e-12, -8.656932e-12, -8.673165e-12, 
    -8.665136e-12, -8.714687e-12, -8.695424e-12, -8.79691e-12, -8.753197e-12, 
    -8.867162e-12, -8.839891e-12, -8.873698e-12, -8.856447e-12, 
    -8.886007e-12, -8.859403e-12, -8.905486e-12, -8.915521e-12, 
    -8.908664e-12, -8.935005e-12, -8.857928e-12, -8.887529e-12, 
    -8.664912e-12, -8.666221e-12, -8.672322e-12, -8.645506e-12, 
    -8.643866e-12, -8.619291e-12, -8.641157e-12, -8.650469e-12, 
    -8.674106e-12, -8.688088e-12, -8.701379e-12, -8.730601e-12, 
    -8.763238e-12, -8.808874e-12, -8.841658e-12, -8.863635e-12, 
    -8.850159e-12, -8.862056e-12, -8.848757e-12, -8.842523e-12, 
    -8.911761e-12, -8.872883e-12, -8.931216e-12, -8.927988e-12, -8.90159e-12, 
    -8.928351e-12, -8.667141e-12, -8.659605e-12, -8.633444e-12, 
    -8.653917e-12, -8.616614e-12, -8.637495e-12, -8.649502e-12, 
    -8.695827e-12, -8.706004e-12, -8.715442e-12, -8.734081e-12, 
    -8.758002e-12, -8.799966e-12, -8.836476e-12, -8.869805e-12, 
    -8.867363e-12, -8.868223e-12, -8.875668e-12, -8.857226e-12, 
    -8.878696e-12, -8.8823e-12, -8.872878e-12, -8.927556e-12, -8.911935e-12, 
    -8.927919e-12, -8.917748e-12, -8.662055e-12, -8.674734e-12, 
    -8.667882e-12, -8.680766e-12, -8.67169e-12, -8.712049e-12, -8.72415e-12, 
    -8.78077e-12, -8.757532e-12, -8.794514e-12, -8.761288e-12, -8.767175e-12, 
    -8.795722e-12, -8.763083e-12, -8.834464e-12, -8.786072e-12, 
    -8.875958e-12, -8.827636e-12, -8.878986e-12, -8.869661e-12, -8.8851e-12, 
    -8.898928e-12, -8.916324e-12, -8.948424e-12, -8.94099e-12, -8.967834e-12, 
    -8.693635e-12, -8.710081e-12, -8.708633e-12, -8.725843e-12, 
    -8.738571e-12, -8.766157e-12, -8.810401e-12, -8.793763e-12, 
    -8.824308e-12, -8.830439e-12, -8.784035e-12, -8.812528e-12, 
    -8.721087e-12, -8.735862e-12, -8.727064e-12, -8.694933e-12, 
    -8.797599e-12, -8.744911e-12, -8.8422e-12, -8.813658e-12, -8.896957e-12, 
    -8.855532e-12, -8.936899e-12, -8.971685e-12, -9.00442e-12, -9.042678e-12, 
    -8.719056e-12, -8.707882e-12, -8.727889e-12, -8.755572e-12, 
    -8.781254e-12, -8.8154e-12, -8.818893e-12, -8.825289e-12, -8.841858e-12, 
    -8.855789e-12, -8.827313e-12, -8.859281e-12, -8.73929e-12, -8.802172e-12, 
    -8.703658e-12, -8.733324e-12, -8.753939e-12, -8.744895e-12, 
    -8.791861e-12, -8.802931e-12, -8.847914e-12, -8.824661e-12, -8.9631e-12, 
    -8.901851e-12, -9.071807e-12, -9.024312e-12, -8.703978e-12, 
    -8.719017e-12, -8.771361e-12, -8.746456e-12, -8.817678e-12, 
    -8.835209e-12, -8.849461e-12, -8.867679e-12, -8.869645e-12, -8.88044e-12, 
    -8.862752e-12, -8.879742e-12, -8.815473e-12, -8.844193e-12, 
    -8.765377e-12, -8.784561e-12, -8.775735e-12, -8.766056e-12, 
    -8.795931e-12, -8.827761e-12, -8.82844e-12, -8.838647e-12, -8.86741e-12, 
    -8.817967e-12, -8.971008e-12, -8.876496e-12, -8.735417e-12, 
    -8.764388e-12, -8.768524e-12, -8.757302e-12, -8.833452e-12, 
    -8.805861e-12, -8.880177e-12, -8.860091e-12, -8.893001e-12, 
    -8.876648e-12, -8.874242e-12, -8.853238e-12, -8.840162e-12, 
    -8.807126e-12, -8.780246e-12, -8.758929e-12, -8.763885e-12, 
    -8.787302e-12, -8.829708e-12, -8.869825e-12, -8.861037e-12, 
    -8.890499e-12, -8.812514e-12, -8.845215e-12, -8.832577e-12, 
    -8.865532e-12, -8.793321e-12, -8.854817e-12, -8.777603e-12, 
    -8.784373e-12, -8.805313e-12, -8.847435e-12, -8.856751e-12, 
    -8.866703e-12, -8.860562e-12, -8.830784e-12, -8.825905e-12, 
    -8.804804e-12, -8.798978e-12, -8.782899e-12, -8.769587e-12, -8.78175e-12, 
    -8.794523e-12, -8.830796e-12, -8.863486e-12, -8.899126e-12, 
    -8.907847e-12, -8.949492e-12, -8.915593e-12, -8.971534e-12, 
    -8.923976e-12, -9.0063e-12, -8.858378e-12, -8.922575e-12, -8.806266e-12, 
    -8.818796e-12, -8.84146e-12, -8.893441e-12, -8.865377e-12, -8.898196e-12, 
    -8.825714e-12, -8.78811e-12, -8.778379e-12, -8.760225e-12, -8.778794e-12, 
    -8.777284e-12, -8.795051e-12, -8.789342e-12, -8.832e-12, -8.809086e-12, 
    -8.874182e-12, -8.897937e-12, -8.965021e-12, -9.006147e-12, 
    -9.048007e-12, -9.066488e-12, -9.072113e-12, -9.074464e-12 ;

 SMIN_NH4 =
  0.0004625543, 0.0004644829, 0.0004641078, 0.0004656634, 0.0004648004, 
    0.0004658189, 0.0004629449, 0.0004645592, 0.0004635286, 0.0004627273, 
    0.0004686815, 0.0004657323, 0.0004717432, 0.0004698628, 0.0004745852, 
    0.0004714506, 0.0004752171, 0.0004744944, 0.0004766685, 0.0004760456, 
    0.0004788265, 0.0004769558, 0.0004802673, 0.0004783795, 0.0004786749, 
    0.0004768938, 0.000466326, 0.0004683149, 0.0004662081, 0.0004664917, 
    0.0004663644, 0.000464818, 0.0004640389, 0.0004624062, 0.0004627025, 
    0.0004639015, 0.0004666189, 0.0004656962, 0.0004680206, 0.0004679681, 
    0.0004705555, 0.0004693889, 0.000473737, 0.0004725011, 0.0004760715, 
    0.0004751736, 0.0004760292, 0.0004757697, 0.0004760325, 0.0004747158, 
    0.0004752798, 0.000474121, 0.0004696081, 0.000470935, 0.0004669772, 
    0.0004645972, 0.0004630156, 0.0004618934, 0.0004620519, 0.0004623544, 
    0.0004639084, 0.0004653691, 0.0004664823, 0.0004672269, 0.0004679604, 
    0.0004701815, 0.0004713562, 0.0004739868, 0.0004735118, 0.0004743162, 
    0.0004750842, 0.0004763739, 0.0004761616, 0.0004767297, 0.0004742945, 
    0.0004759131, 0.0004732409, 0.0004739718, 0.0004681613, 0.0004659453, 
    0.0004650041, 0.0004641795, 0.0004621738, 0.0004635589, 0.0004630129, 
    0.0004643115, 0.0004651367, 0.0004647284, 0.0004672472, 0.0004662679, 
    0.0004714258, 0.0004692043, 0.0004749947, 0.0004736092, 0.0004753266, 
    0.0004744502, 0.0004759517, 0.0004746003, 0.000476941, 0.0004774508, 
    0.0004771024, 0.0004784401, 0.000474525, 0.0004760288, 0.0004647174, 
    0.000464784, 0.000465094, 0.0004637308, 0.0004636474, 0.0004623978, 
    0.0004635094, 0.0004639829, 0.0004651843, 0.000465895, 0.0004665705, 
    0.0004680559, 0.0004697145, 0.0004720334, 0.000473699, 0.0004748153, 
    0.0004741306, 0.000474735, 0.0004740593, 0.0004737425, 0.0004772597, 
    0.0004752849, 0.0004782476, 0.0004780836, 0.0004767428, 0.0004781019, 
    0.0004648306, 0.0004644474, 0.0004631174, 0.0004641581, 0.0004622616, 
    0.0004633233, 0.0004639337, 0.0004662885, 0.0004668056, 0.0004672853, 
    0.0004682326, 0.0004694482, 0.0004715807, 0.0004734356, 0.0004751286, 
    0.0004750045, 0.0004750481, 0.0004754264, 0.0004744894, 0.00047558, 
    0.0004757631, 0.0004752844, 0.0004780615, 0.0004772681, 0.0004780799, 
    0.0004775632, 0.0004645718, 0.0004652163, 0.000464868, 0.000465523, 
    0.0004650615, 0.0004671131, 0.0004677281, 0.0004706054, 0.0004694243, 
    0.0004713037, 0.000469615, 0.0004699143, 0.0004713651, 0.0004697061, 
    0.0004733333, 0.0004708745, 0.000475441, 0.0004729863, 0.0004755947, 
    0.0004751208, 0.000475905, 0.0004766076, 0.0004774909, 0.0004791213, 
    0.0004787436, 0.0004801068, 0.0004661771, 0.000467013, 0.0004669392, 
    0.0004678139, 0.0004684608, 0.0004698627, 0.0004721109, 0.0004712653, 
    0.0004728172, 0.0004731288, 0.0004707708, 0.0004722187, 0.0004675718, 
    0.0004683227, 0.0004678754, 0.0004662422, 0.0004714599, 0.0004687824, 
    0.0004737258, 0.0004722756, 0.0004765072, 0.0004744031, 0.0004785358, 
    0.0004803026, 0.0004819644, 0.000483907, 0.000467469, 0.0004669009, 
    0.0004679178, 0.0004693249, 0.0004706297, 0.0004723648, 0.0004725421, 
    0.000472867, 0.0004737087, 0.0004744165, 0.0004729698, 0.0004745937, 
    0.0004684972, 0.0004716922, 0.0004666856, 0.0004681936, 0.0004692411, 
    0.0004687814, 0.0004711679, 0.0004717303, 0.0004740158, 0.0004728343, 
    0.0004798665, 0.0004767557, 0.0004853854, 0.0004829744, 0.0004667024, 
    0.0004674668, 0.0004701271, 0.0004688613, 0.0004724803, 0.0004733711, 
    0.0004740949, 0.0004750206, 0.0004751202, 0.0004756686, 0.0004747699, 
    0.000475633, 0.0004723678, 0.000473827, 0.0004698222, 0.000470797, 
    0.0004703485, 0.0004698565, 0.0004713745, 0.000472992, 0.0004730262, 
    0.0004735448, 0.0004750067, 0.0004724939, 0.0004802683, 0.0004754679, 
    0.0004683002, 0.0004697727, 0.0004699826, 0.0004694123, 0.0004732816, 
    0.0004718798, 0.0004756553, 0.0004746348, 0.0004763064, 0.0004754758, 
    0.0004753535, 0.0004742865, 0.0004736221, 0.0004719436, 0.0004705777, 
    0.0004694943, 0.0004697461, 0.0004709361, 0.0004730907, 0.0004751287, 
    0.0004746823, 0.0004761787, 0.0004722168, 0.0004738783, 0.0004732361, 
    0.0004749103, 0.0004712427, 0.0004743677, 0.0004704438, 0.0004707878, 
    0.0004718518, 0.0004739921, 0.000474465, 0.0004749706, 0.0004746585, 
    0.0004731458, 0.0004728978, 0.0004718255, 0.0004715295, 0.0004707123, 
    0.0004700358, 0.0004706539, 0.0004713029, 0.0004731459, 0.0004748066, 
    0.0004766169, 0.0004770597, 0.0004791752, 0.0004774534, 0.0004802948, 
    0.0004778796, 0.0004820597, 0.0004745482, 0.0004778092, 0.0004719001, 
    0.0004725367, 0.0004736884, 0.0004763289, 0.0004749031, 0.0004765704, 
    0.000472888, 0.0004709774, 0.0004704826, 0.0004695602, 0.0004705036, 
    0.0004704268, 0.0004713296, 0.0004710394, 0.0004732069, 0.0004720426, 
    0.0004753497, 0.0004765565, 0.0004799634, 0.0004820517, 0.0004841767, 
    0.0004851148, 0.0004854003, 0.0004855196 ;

 SMIN_NH4_vr =
  0.003061824, 0.003066965, 0.003065959, 0.003070103, 0.0030678, 0.003070507, 
    0.00306285, 0.003067148, 0.003064399, 0.003062258, 0.003078107, 
    0.003070261, 0.003086228, 0.003081233, 0.003093749, 0.003085444, 
    0.003095417, 0.003093499, 0.003099248, 0.003097596, 0.003104943, 
    0.003099999, 0.003108737, 0.003103756, 0.003104532, 0.003099821, 
    0.003071862, 0.003077156, 0.003071543, 0.003072298, 0.003071955, 
    0.003067834, 0.003065759, 0.0030614, 0.003062186, 0.003065384, 
    0.003072614, 0.003070153, 0.003076331, 0.003076193, 0.003083058, 
    0.003079962, 0.003091489, 0.00308821, 0.003097661, 0.003095282, 
    0.003097544, 0.003096852, 0.003097543, 0.003094061, 0.003095547, 
    0.00309248, 0.003080581, 0.003084098, 0.003073583, 0.003067246, 
    0.003063025, 0.003060032, 0.003060449, 0.003061257, 0.003065396, 
    0.003069281, 0.003072242, 0.003074217, 0.003076163, 0.003082067, 
    0.003085179, 0.003092145, 0.003090885, 0.003093011, 0.003095041, 
    0.003098448, 0.003097885, 0.003099383, 0.003092936, 0.003097221, 
    0.003090139, 0.003092076, 0.003076734, 0.00307083, 0.003068326, 
    0.003066123, 0.003060772, 0.003064466, 0.003063007, 0.003066462, 
    0.003068658, 0.003067566, 0.003074268, 0.003071658, 0.003085358, 
    0.003079462, 0.003094809, 0.003091136, 0.003095678, 0.003093359, 
    0.003097326, 0.00309375, 0.003099935, 0.003101284, 0.003100356, 
    0.00310389, 0.003093532, 0.003097512, 0.003067555, 0.003067733, 
    0.003068554, 0.003064919, 0.003064696, 0.003061359, 0.003064319, 
    0.003065581, 0.003068776, 0.003070664, 0.003072457, 0.003076408, 
    0.003080811, 0.003086959, 0.00309137, 0.00309432, 0.003092506, 
    0.003094102, 0.003092312, 0.003091468, 0.00310077, 0.003095548, 
    0.003103373, 0.00310294, 0.003099394, 0.00310298, 0.003067851, 
    0.003066825, 0.00306328, 0.003066049, 0.003060989, 0.003063821, 
    0.003065445, 0.00307171, 0.00307308, 0.003074357, 0.003076871, 
    0.003080096, 0.003085754, 0.003090666, 0.003095146, 0.003094813, 
    0.003094927, 0.003095923, 0.003093442, 0.003096324, 0.003096804, 
    0.003095538, 0.003102873, 0.003100778, 0.003102918, 0.003101548, 
    0.003067153, 0.003068865, 0.003067933, 0.003069678, 0.003068443, 
    0.003073904, 0.003075536, 0.003083173, 0.003080033, 0.003085022, 
    0.003080533, 0.003081328, 0.003085177, 0.003080766, 0.003090387, 
    0.003083864, 0.003095959, 0.003089458, 0.003096359, 0.0030951, 
    0.003097171, 0.00309903, 0.003101357, 0.003105665, 0.00310466, 
    0.003108258, 0.003071419, 0.003073639, 0.00307344, 0.003075761, 
    0.003077477, 0.003081201, 0.003087162, 0.003084914, 0.003089024, 
    0.003089851, 0.003083592, 0.003087434, 0.003075093, 0.003077085, 
    0.003075894, 0.003071545, 0.003085406, 0.003078294, 0.003091404, 
    0.003087557, 0.003098756, 0.00309319, 0.003104109, 0.003108775, 
    0.003113149, 0.003118261, 0.003074847, 0.003073331, 0.003076031, 
    0.003079772, 0.003083228, 0.00308783, 0.003088296, 0.003089153, 
    0.003091378, 0.003093253, 0.003089419, 0.003093713, 0.003077547, 
    0.003086021, 0.003072718, 0.00307673, 0.003079505, 0.003078284, 
    0.003084615, 0.003086102, 0.003092156, 0.003089025, 0.003107616, 
    0.0030994, 0.003122141, 0.0031158, 0.0030728, 0.003074828, 0.003081892, 
    0.003078531, 0.003088127, 0.003090489, 0.003092398, 0.00309485, 
    0.003095107, 0.003096559, 0.003094173, 0.003096458, 0.003087805, 
    0.003091672, 0.003081048, 0.003083631, 0.003082439, 0.003081128, 
    0.003085152, 0.003089443, 0.003089528, 0.003090898, 0.003094772, 
    0.003088106, 0.003108667, 0.003095981, 0.00307704, 0.003080948, 
    0.0030815, 0.003079986, 0.003090243, 0.003086528, 0.003096523, 
    0.003093818, 0.003098236, 0.00309604, 0.003095709, 0.003092886, 
    0.00309112, 0.003086673, 0.003083043, 0.003080167, 0.003080829, 
    0.003083989, 0.003089695, 0.003095092, 0.003093906, 0.003097859, 
    0.003087366, 0.00309177, 0.003090062, 0.003094495, 0.003084842, 
    0.003093128, 0.003082718, 0.003083626, 0.003086445, 0.003092119, 
    0.003093362, 0.003094702, 0.003093868, 0.003089864, 0.003089202, 
    0.003086354, 0.003085566, 0.003083398, 0.003081596, 0.003083237, 
    0.003084953, 0.003089839, 0.003094233, 0.003099017, 0.003100185, 
    0.003105771, 0.003101222, 0.003108722, 0.003102346, 0.003113366, 
    0.003093595, 0.00310222, 0.003086573, 0.003088256, 0.003091308, 
    0.003098291, 0.003094513, 0.003098926, 0.003089174, 0.003084104, 
    0.003082786, 0.003080338, 0.003082835, 0.003082632, 0.003085023, 
    0.003084249, 0.003089992, 0.003086906, 0.003095659, 0.003098852, 
    0.003107845, 0.003113346, 0.003118938, 0.0031214, 0.003122149, 0.003122459,
  0.001811062, 0.001817816, 0.001816503, 0.001821947, 0.001818927, 
    0.001822492, 0.001812431, 0.001818084, 0.001814476, 0.001811669, 
    0.0018325, 0.00182219, 0.001843187, 0.001836626, 0.001853092, 
    0.001842167, 0.001855292, 0.001852776, 0.001860343, 0.001858176, 
    0.001867847, 0.001861343, 0.001872851, 0.001866293, 0.00186732, 
    0.001861128, 0.001824265, 0.001831218, 0.001823853, 0.001824845, 
    0.0018244, 0.00181899, 0.001816263, 0.001810544, 0.001811583, 
    0.001815782, 0.001825291, 0.001822064, 0.001830191, 0.001830008, 
    0.001839044, 0.001834971, 0.001850138, 0.001845831, 0.001858267, 
    0.001855142, 0.00185812, 0.001857217, 0.001858132, 0.001853548, 
    0.001855512, 0.001851477, 0.001835735, 0.001840366, 0.001826543, 
    0.001818218, 0.001812679, 0.001808747, 0.001809303, 0.001810363, 
    0.001815807, 0.00182092, 0.001824814, 0.001827418, 0.001829982, 
    0.001837739, 0.001841838, 0.001851009, 0.001849354, 0.001852156, 
    0.001854831, 0.00185932, 0.001858581, 0.001860558, 0.001852082, 
    0.001857717, 0.001848411, 0.001850958, 0.001830682, 0.001822935, 
    0.001819642, 0.001816756, 0.001809731, 0.001814583, 0.001812671, 
    0.001817218, 0.001820107, 0.001818678, 0.001827489, 0.001824065, 
    0.001842081, 0.001834328, 0.001854519, 0.001849693, 0.001855675, 
    0.001852623, 0.001857851, 0.001853146, 0.001861293, 0.001863066, 
    0.001861855, 0.001866506, 0.001852885, 0.00185812, 0.001818639, 
    0.001818872, 0.001819957, 0.001815185, 0.001814893, 0.001810516, 
    0.001814411, 0.001816069, 0.001820274, 0.001822761, 0.001825124, 
    0.001830316, 0.00183611, 0.001844201, 0.001850006, 0.001853895, 
    0.00185151, 0.001853616, 0.001851262, 0.001850159, 0.001862402, 
    0.001855531, 0.001865837, 0.001865267, 0.001860605, 0.001865331, 
    0.001819035, 0.001817694, 0.001813037, 0.001816682, 0.001810039, 
    0.001813759, 0.001815897, 0.001824138, 0.001825946, 0.001827623, 
    0.001830934, 0.00183518, 0.001842622, 0.001849089, 0.001854986, 
    0.001854554, 0.001854706, 0.001856023, 0.001852761, 0.001856559, 
    0.001857196, 0.00185553, 0.001865191, 0.001862432, 0.001865255, 
    0.001863459, 0.00181813, 0.001820386, 0.001819167, 0.001821459, 
    0.001819845, 0.001827021, 0.001829171, 0.00183922, 0.001835097, 
    0.001841656, 0.001835763, 0.001836808, 0.001841871, 0.001836081, 
    0.001848734, 0.00184016, 0.001856075, 0.001847525, 0.00185661, 
    0.001854961, 0.001857691, 0.001860135, 0.001863208, 0.001868874, 
    0.001867562, 0.001872297, 0.001823747, 0.001826671, 0.001826413, 
    0.001829471, 0.001831731, 0.001836627, 0.001844471, 0.001841522, 
    0.001846934, 0.00184802, 0.001839797, 0.001844848, 0.001828626, 
    0.001831251, 0.001829688, 0.001823978, 0.001842203, 0.001832857, 
    0.001850102, 0.001845048, 0.001859787, 0.001852462, 0.00186684, 
    0.001872978, 0.001878744, 0.00188548, 0.001828265, 0.001826279, 
    0.001829834, 0.001834749, 0.001839305, 0.001845357, 0.001845975, 
    0.001847108, 0.001850041, 0.001852507, 0.001847467, 0.001853125, 
    0.001831861, 0.001843013, 0.001825529, 0.0018308, 0.001834459, 
    0.001832854, 0.001841185, 0.001843147, 0.001851114, 0.001846996, 
    0.001871464, 0.001860652, 0.0018906, 0.001882248, 0.001825585, 
    0.001828258, 0.001837551, 0.001833131, 0.00184576, 0.001848865, 
    0.001851387, 0.001854611, 0.001854958, 0.001856867, 0.001853739, 
    0.001856743, 0.001845369, 0.001850455, 0.001836488, 0.001839891, 
    0.001838326, 0.001836609, 0.001841906, 0.001847547, 0.001847666, 
    0.001849474, 0.001854566, 0.001845811, 0.00187286, 0.001856172, 
    0.001831171, 0.001836314, 0.001837047, 0.001835055, 0.001848554, 
    0.001843667, 0.00185682, 0.001853268, 0.001859087, 0.001856196, 
    0.001855771, 0.001852056, 0.001849742, 0.001843891, 0.001839126, 
    0.001835344, 0.001836224, 0.001840377, 0.001847891, 0.00185499, 
    0.001853436, 0.001858645, 0.001844845, 0.001850636, 0.001848399, 
    0.001854231, 0.001841444, 0.001852338, 0.001838657, 0.001839857, 
    0.001843569, 0.00185103, 0.001852677, 0.001854438, 0.001853351, 
    0.001848082, 0.001847217, 0.001843479, 0.001842447, 0.001839596, 
    0.001837235, 0.001839392, 0.001841657, 0.001848083, 0.001853869, 
    0.00186017, 0.00186171, 0.001869064, 0.00186308, 0.001872953, 
    0.001864563, 0.001879078, 0.001852967, 0.001864314, 0.001843738, 
    0.001845958, 0.001849972, 0.001859166, 0.001854203, 0.001860006, 
    0.001847183, 0.001840521, 0.001838794, 0.001835574, 0.001838868, 
    0.0018386, 0.00184175, 0.001840738, 0.001848297, 0.001844238, 
    0.001855761, 0.00185996, 0.001871802, 0.00187905, 0.001886416, 
    0.001889665, 0.001890654, 0.001891067,
  0.001646651, 0.001653856, 0.001652455, 0.001658264, 0.001655042, 
    0.001658845, 0.001648112, 0.001654142, 0.001650293, 0.001647299, 
    0.001669527, 0.001658523, 0.001680939, 0.001673932, 0.001691522, 
    0.00167985, 0.001693874, 0.001691185, 0.001699273, 0.001696957, 
    0.001707296, 0.001700342, 0.001712649, 0.001705635, 0.001706733, 
    0.001700113, 0.001660738, 0.001668158, 0.001660298, 0.001661357, 
    0.001660881, 0.001655109, 0.001652199, 0.001646099, 0.001647207, 
    0.001651686, 0.001661832, 0.001658389, 0.001667063, 0.001666867, 
    0.001676515, 0.001672166, 0.001688366, 0.001683764, 0.001697053, 
    0.001693713, 0.001696897, 0.001695931, 0.001696909, 0.00169201, 
    0.00169411, 0.001689797, 0.001672981, 0.001677927, 0.001663169, 
    0.001654284, 0.001648376, 0.001644183, 0.001644776, 0.001645906, 
    0.001651713, 0.001657168, 0.001661323, 0.001664102, 0.001666839, 
    0.001675121, 0.001679499, 0.001689296, 0.001687528, 0.001690522, 
    0.001693381, 0.001698179, 0.001697389, 0.001699503, 0.001690443, 
    0.001696466, 0.001686521, 0.001689242, 0.001667586, 0.001659318, 
    0.001655804, 0.001652725, 0.001645232, 0.001650407, 0.001648367, 
    0.001653219, 0.001656301, 0.001654776, 0.001664178, 0.001660524, 
    0.001679759, 0.001671479, 0.001693048, 0.001687891, 0.001694283, 
    0.001691022, 0.001696609, 0.001691581, 0.001700289, 0.001702184, 
    0.001700889, 0.001705862, 0.001691302, 0.001696897, 0.001654734, 
    0.001654982, 0.00165614, 0.001651049, 0.001650738, 0.001646069, 
    0.001650223, 0.001651992, 0.001656479, 0.001659133, 0.001661654, 
    0.001667196, 0.001673381, 0.001682023, 0.001688225, 0.001692381, 
    0.001689833, 0.001692083, 0.001689568, 0.001688389, 0.001701474, 
    0.001694129, 0.001705147, 0.001704538, 0.001699553, 0.001704606, 
    0.001655157, 0.001653726, 0.001648758, 0.001652646, 0.001645561, 
    0.001649528, 0.001651808, 0.001660601, 0.001662531, 0.001664322, 
    0.001667855, 0.001672389, 0.001680337, 0.001687245, 0.001693547, 
    0.001693086, 0.001693248, 0.001694656, 0.001691169, 0.001695228, 
    0.001695909, 0.001694128, 0.001704456, 0.001701507, 0.001704525, 
    0.001702604, 0.001654191, 0.001656598, 0.001655298, 0.001657743, 
    0.001656021, 0.001663679, 0.001665973, 0.001676702, 0.0016723, 
    0.001679305, 0.001673011, 0.001674127, 0.001679534, 0.001673352, 
    0.001686865, 0.001677707, 0.00169471, 0.001685574, 0.001695283, 
    0.00169352, 0.001696438, 0.001699051, 0.001702336, 0.001708395, 
    0.001706992, 0.001712057, 0.001660185, 0.001663305, 0.00166303, 
    0.001666293, 0.001668707, 0.001673934, 0.001682312, 0.001679162, 
    0.001684943, 0.001686103, 0.00167732, 0.001682714, 0.001665392, 
    0.001668193, 0.001666525, 0.001660431, 0.001679889, 0.001669909, 
    0.001688328, 0.001682928, 0.001698678, 0.001690849, 0.00170622, 
    0.001712784, 0.001718954, 0.001726162, 0.001665007, 0.001662887, 
    0.001666681, 0.001671929, 0.001676794, 0.001683258, 0.001683918, 
    0.001685129, 0.001688263, 0.001690898, 0.001685512, 0.001691558, 
    0.001668844, 0.001680754, 0.001662086, 0.001667712, 0.001671619, 
    0.001669905, 0.001678802, 0.001680898, 0.001689409, 0.00168501, 
    0.001711165, 0.001699603, 0.001731644, 0.001722703, 0.001662147, 
    0.001664999, 0.00167492, 0.001670201, 0.001683689, 0.001687006, 
    0.001689701, 0.001693146, 0.001693517, 0.001695557, 0.001692214, 
    0.001695425, 0.001683271, 0.001688705, 0.001673786, 0.00167742, 
    0.001675748, 0.001673914, 0.001679572, 0.001685597, 0.001685725, 
    0.001687656, 0.001693097, 0.001683743, 0.001712657, 0.001694814, 
    0.001668109, 0.001673599, 0.001674382, 0.001672256, 0.001686673, 
    0.001681452, 0.001695508, 0.001691711, 0.001697931, 0.00169484, 
    0.001694386, 0.001690415, 0.001687943, 0.001681692, 0.001676603, 
    0.001672564, 0.001673504, 0.001677939, 0.001685965, 0.001693551, 
    0.00169189, 0.001697458, 0.001682711, 0.001688898, 0.001686508, 
    0.00169274, 0.001679079, 0.001690715, 0.001676102, 0.001677384, 
    0.001681349, 0.001689318, 0.001691079, 0.001692961, 0.0016918, 
    0.001686169, 0.001685246, 0.001681252, 0.00168015, 0.001677105, 
    0.001674584, 0.001676887, 0.001679306, 0.001686171, 0.001692353, 
    0.001699088, 0.001700735, 0.001708598, 0.001702199, 0.001712757, 
    0.001703783, 0.00171931, 0.001691388, 0.001703517, 0.001681529, 
    0.0016839, 0.001688188, 0.001698014, 0.00169271, 0.001698913, 
    0.001685209, 0.001678092, 0.001676249, 0.00167281, 0.001676327, 
    0.001676041, 0.001679406, 0.001678325, 0.001686399, 0.001682063, 
    0.001694375, 0.001698863, 0.001711526, 0.00171928, 0.001727164, 
    0.001730643, 0.001731701, 0.001732144,
  0.001515203, 0.001522335, 0.001520949, 0.0015267, 0.001523509, 0.001527275, 
    0.001516649, 0.001522618, 0.001518808, 0.001515845, 0.001537858, 
    0.001526956, 0.001549174, 0.001542225, 0.001559675, 0.001548093, 
    0.00156201, 0.00155934, 0.001567372, 0.001565071, 0.001575342, 
    0.001568433, 0.001580663, 0.001573692, 0.001574783, 0.001568206, 
    0.00152915, 0.001536501, 0.001528714, 0.001529763, 0.001529292, 
    0.001523576, 0.001520695, 0.001514658, 0.001515754, 0.001520187, 
    0.001530234, 0.001526824, 0.001535417, 0.001535223, 0.001544786, 
    0.001540475, 0.001556542, 0.001551976, 0.001565167, 0.001561851, 
    0.001565011, 0.001564053, 0.001565024, 0.00156016, 0.001562244, 
    0.001557963, 0.001541282, 0.001546186, 0.001531558, 0.001522759, 
    0.001516911, 0.001512761, 0.001513348, 0.001514466, 0.001520213, 
    0.001525615, 0.00152973, 0.001532483, 0.001535195, 0.001543403, 
    0.001547745, 0.001557466, 0.001555711, 0.001558683, 0.001561521, 
    0.001566285, 0.001565501, 0.0015676, 0.001558604, 0.001564583, 
    0.001554712, 0.001557412, 0.001535934, 0.001527744, 0.001524264, 
    0.001521215, 0.001513799, 0.001518921, 0.001516902, 0.001521704, 
    0.001524755, 0.001523246, 0.001532558, 0.001528938, 0.001548003, 
    0.001539793, 0.00156119, 0.001556071, 0.001562416, 0.001559179, 
    0.001564726, 0.001559733, 0.001568381, 0.001570263, 0.001568977, 
    0.001573918, 0.001559457, 0.001565012, 0.001523204, 0.00152345, 
    0.001524597, 0.001519557, 0.001519248, 0.001514628, 0.001518739, 
    0.00152049, 0.001524932, 0.00152756, 0.001530058, 0.001535548, 
    0.001541679, 0.001550249, 0.001556403, 0.001560528, 0.001557998, 
    0.001560231, 0.001557735, 0.001556565, 0.001569558, 0.001562264, 
    0.001573207, 0.001572602, 0.00156765, 0.00157267, 0.001523623, 
    0.001522207, 0.001517289, 0.001521138, 0.001514125, 0.001518051, 
    0.001520308, 0.001529015, 0.001530927, 0.0015327, 0.001536202, 
    0.001540695, 0.001548576, 0.00155543, 0.001561686, 0.001561227, 
    0.001561389, 0.001562786, 0.001559325, 0.001563354, 0.001564031, 
    0.001562262, 0.001572521, 0.00156959, 0.001572589, 0.001570681, 
    0.001522667, 0.00152505, 0.001523762, 0.001526184, 0.001524478, 
    0.001532063, 0.001534337, 0.001544972, 0.001540607, 0.001547552, 
    0.001541312, 0.001542418, 0.00154778, 0.001541649, 0.001555053, 
    0.001545968, 0.00156284, 0.001553772, 0.001563409, 0.001561659, 
    0.001564556, 0.00156715, 0.001570414, 0.001576435, 0.001575041, 
    0.001580075, 0.001528602, 0.001531693, 0.00153142, 0.001534654, 
    0.001537045, 0.001542227, 0.001550535, 0.001547411, 0.001553146, 
    0.001554297, 0.001545584, 0.001550935, 0.001533761, 0.001536537, 
    0.001534884, 0.001528846, 0.001548132, 0.001538237, 0.001556505, 
    0.001551147, 0.001566781, 0.001559007, 0.001574273, 0.001580797, 
    0.001586934, 0.001594105, 0.001533379, 0.001531279, 0.001535038, 
    0.001540239, 0.001545062, 0.001551474, 0.001552129, 0.00155333, 
    0.00155644, 0.001559055, 0.001553711, 0.001559711, 0.001537182, 
    0.00154899, 0.001530486, 0.00153606, 0.001539932, 0.001538233, 
    0.001547054, 0.001549133, 0.001557578, 0.001553212, 0.001579188, 
    0.001567699, 0.001599562, 0.001590663, 0.001530546, 0.001533372, 
    0.001543205, 0.001538526, 0.001551901, 0.001555193, 0.001557868, 
    0.001561287, 0.001561656, 0.001563682, 0.001560362, 0.00156355, 
    0.001551487, 0.001556879, 0.00154208, 0.001545683, 0.001544026, 
    0.001542208, 0.001547818, 0.001553795, 0.001553922, 0.001555838, 
    0.001561238, 0.001551956, 0.001580672, 0.001562943, 0.001536453, 
    0.001541895, 0.001542671, 0.001540564, 0.001554863, 0.001549683, 
    0.001563632, 0.001559863, 0.001566038, 0.00156297, 0.001562518, 
    0.001558576, 0.001556122, 0.00154992, 0.001544873, 0.001540869, 
    0.0015418, 0.001546198, 0.00155416, 0.00156169, 0.001560041, 0.001565569, 
    0.001550932, 0.001557071, 0.001554699, 0.001560884, 0.001547328, 
    0.001558874, 0.001544376, 0.001545648, 0.00154958, 0.001557488, 
    0.001559236, 0.001561104, 0.001559951, 0.001554362, 0.001553446, 
    0.001549484, 0.001548391, 0.001545371, 0.001542871, 0.001545155, 
    0.001547554, 0.001554364, 0.0015605, 0.001567188, 0.001568824, 
    0.001576636, 0.001570278, 0.00158077, 0.001571851, 0.001587288, 
    0.001559542, 0.001571588, 0.001549759, 0.001552111, 0.001556366, 
    0.001566121, 0.001560855, 0.001567014, 0.00155341, 0.00154635, 
    0.001544522, 0.001541113, 0.0015446, 0.001544316, 0.001547653, 
    0.001546581, 0.00155459, 0.001550288, 0.001562507, 0.001566965, 
    0.001579547, 0.001587258, 0.001595103, 0.001598565, 0.001599619, 
    0.00160006,
  0.001379622, 0.001386014, 0.001384771, 0.001389929, 0.001387067, 
    0.001390446, 0.001380917, 0.001386268, 0.001382852, 0.001380197, 
    0.001399948, 0.001390159, 0.001410122, 0.001403872, 0.001419577, 
    0.001409149, 0.001421681, 0.001419275, 0.001426515, 0.00142444, 
    0.001433707, 0.001427472, 0.001438514, 0.001432218, 0.001433203, 
    0.001427267, 0.001392128, 0.001398729, 0.001391737, 0.001392678, 
    0.001392256, 0.001387127, 0.001384543, 0.001379133, 0.001380115, 
    0.001384089, 0.001393101, 0.00139004, 0.001397754, 0.00139758, 
    0.001406175, 0.001402299, 0.001416755, 0.001412644, 0.001424527, 
    0.001421537, 0.001424387, 0.001423522, 0.001424398, 0.001420013, 
    0.001421892, 0.001418034, 0.001403025, 0.001407434, 0.001394289, 
    0.001386394, 0.001381152, 0.001377434, 0.00137796, 0.001378962, 
    0.001384112, 0.001388956, 0.001392649, 0.00139512, 0.001397555, 
    0.001404932, 0.001408837, 0.001417586, 0.001416006, 0.001418683, 
    0.00142124, 0.001425535, 0.001424828, 0.001426721, 0.001418612, 0.001424, 
    0.001415106, 0.001417538, 0.001398219, 0.001390866, 0.001387744, 
    0.00138501, 0.001378364, 0.001382953, 0.001381144, 0.001385449, 
    0.001388185, 0.001386831, 0.001395187, 0.001391938, 0.001409068, 
    0.001401686, 0.001420942, 0.00141633, 0.001422047, 0.001419129, 
    0.001424129, 0.001419629, 0.001427425, 0.001429124, 0.001427963, 
    0.001432422, 0.00141938, 0.001424387, 0.001386794, 0.001387014, 
    0.001388043, 0.001383523, 0.001383247, 0.001379106, 0.00138279, 
    0.00138436, 0.001388344, 0.001390701, 0.001392943, 0.001397872, 
    0.001403381, 0.001411089, 0.001416629, 0.001420345, 0.001418066, 
    0.001420078, 0.001417829, 0.001416775, 0.001428487, 0.001421909, 
    0.00143178, 0.001431233, 0.001426766, 0.001431295, 0.001387169, 
    0.001385899, 0.001381491, 0.00138494, 0.001378656, 0.001382173, 
    0.001384197, 0.001392007, 0.001393722, 0.001395315, 0.00139846, 
    0.001402497, 0.001409584, 0.001415754, 0.001421388, 0.001420975, 
    0.001421121, 0.00142238, 0.001419261, 0.001422892, 0.001423502, 
    0.001421908, 0.00143116, 0.001428516, 0.001431222, 0.0014295, 
    0.001386312, 0.001388449, 0.001387294, 0.001389467, 0.001387936, 
    0.001394743, 0.001396784, 0.001406342, 0.001402418, 0.001408663, 
    0.001403052, 0.001404046, 0.001408868, 0.001403355, 0.001415414, 
    0.001407237, 0.001422429, 0.00141426, 0.001422941, 0.001421364, 
    0.001423976, 0.001426315, 0.001429259, 0.001434694, 0.001433435, 
    0.001437982, 0.001391636, 0.001394411, 0.001394166, 0.001397069, 
    0.001399217, 0.001403874, 0.001411347, 0.001408536, 0.001413696, 
    0.001414733, 0.001406893, 0.001411706, 0.001396267, 0.001398761, 
    0.001397276, 0.001391856, 0.001409184, 0.001400288, 0.001416721, 
    0.001411897, 0.001425982, 0.001418975, 0.001432742, 0.001438635, 
    0.001444181, 0.00145067, 0.001395924, 0.001394039, 0.001397415, 
    0.001402087, 0.001406423, 0.001412191, 0.001412781, 0.001413863, 
    0.001416663, 0.001419018, 0.001414205, 0.001419609, 0.00139934, 
    0.001409956, 0.001393327, 0.001398332, 0.001401811, 0.001400285, 
    0.001408214, 0.001410084, 0.001417687, 0.001413756, 0.001437181, 
    0.00142681, 0.001455612, 0.001447555, 0.001393381, 0.001395918, 
    0.001404753, 0.001400548, 0.001412576, 0.001415539, 0.001417948, 
    0.001421029, 0.001421362, 0.001423187, 0.001420196, 0.001423069, 
    0.001412204, 0.001417058, 0.001403742, 0.001406982, 0.001405491, 
    0.001403857, 0.001408902, 0.001414281, 0.001414395, 0.00141612, 
    0.001420985, 0.001412625, 0.001438521, 0.001422522, 0.001398685, 
    0.001403576, 0.001404273, 0.001402379, 0.001415242, 0.00141058, 
    0.001423143, 0.001419746, 0.001425312, 0.001422546, 0.001422139, 
    0.001418587, 0.001416376, 0.001410793, 0.001406253, 0.001402653, 
    0.00140349, 0.001407445, 0.00141461, 0.001421392, 0.001419906, 
    0.001424889, 0.001411704, 0.001417231, 0.001415094, 0.001420666, 
    0.001408461, 0.001418856, 0.001405806, 0.00140695, 0.001410487, 
    0.001417606, 0.001419181, 0.001420864, 0.001419825, 0.001414791, 
    0.001413967, 0.001410401, 0.001409417, 0.001406701, 0.001404453, 
    0.001406507, 0.001408664, 0.001414793, 0.00142032, 0.001426349, 
    0.001427824, 0.001434876, 0.001429136, 0.001438611, 0.001430557, 
    0.001444502, 0.001419457, 0.001430318, 0.001410648, 0.001412765, 
    0.001416596, 0.001425387, 0.00142064, 0.001426192, 0.001413934, 
    0.001407581, 0.001405937, 0.001402872, 0.001406007, 0.001405752, 
    0.001408753, 0.001407789, 0.001414997, 0.001411124, 0.001422129, 
    0.001426148, 0.001437505, 0.001444475, 0.001451573, 0.001454709, 
    0.001455664, 0.001456063,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.355651e-06, 1.367222e-06, 1.364968e-06, 1.374331e-06, 1.369132e-06, 
    1.375269e-06, 1.357991e-06, 1.367682e-06, 1.361491e-06, 1.356688e-06, 
    1.392593e-06, 1.374748e-06, 1.411247e-06, 1.399776e-06, 1.42868e-06, 
    1.409459e-06, 1.432571e-06, 1.428122e-06, 1.44153e-06, 1.437682e-06, 
    1.454904e-06, 1.443307e-06, 1.46387e-06, 1.452129e-06, 1.453963e-06, 
    1.442925e-06, 1.378329e-06, 1.390366e-06, 1.377618e-06, 1.379331e-06, 
    1.378561e-06, 1.369239e-06, 1.364555e-06, 1.354766e-06, 1.35654e-06, 
    1.36373e-06, 1.3801e-06, 1.374531e-06, 1.388585e-06, 1.388267e-06, 
    1.403997e-06, 1.396893e-06, 1.423466e-06, 1.415887e-06, 1.437843e-06, 
    1.432305e-06, 1.437582e-06, 1.43598e-06, 1.437602e-06, 1.429486e-06, 
    1.43296e-06, 1.425828e-06, 1.398224e-06, 1.40631e-06, 1.382265e-06, 
    1.367911e-06, 1.358415e-06, 1.351699e-06, 1.352647e-06, 1.354456e-06, 
    1.363772e-06, 1.372559e-06, 1.379276e-06, 1.383778e-06, 1.38822e-06, 
    1.401717e-06, 1.408884e-06, 1.425002e-06, 1.422085e-06, 1.427027e-06, 
    1.431754e-06, 1.439711e-06, 1.4384e-06, 1.441911e-06, 1.426894e-06, 
    1.436866e-06, 1.420424e-06, 1.424911e-06, 1.389435e-06, 1.376033e-06, 
    1.370359e-06, 1.3654e-06, 1.353376e-06, 1.361674e-06, 1.3584e-06, 
    1.366194e-06, 1.371159e-06, 1.368702e-06, 1.383901e-06, 1.377982e-06, 
    1.409309e-06, 1.395771e-06, 1.431203e-06, 1.422683e-06, 1.433248e-06, 
    1.427852e-06, 1.437104e-06, 1.428775e-06, 1.443218e-06, 1.446373e-06, 
    1.444216e-06, 1.452508e-06, 1.428313e-06, 1.437581e-06, 1.368634e-06, 
    1.369035e-06, 1.370901e-06, 1.362706e-06, 1.362205e-06, 1.354717e-06, 
    1.361378e-06, 1.36422e-06, 1.371447e-06, 1.375731e-06, 1.37981e-06, 
    1.3888e-06, 1.398875e-06, 1.413025e-06, 1.423234e-06, 1.430099e-06, 
    1.425887e-06, 1.429605e-06, 1.425449e-06, 1.423503e-06, 1.44519e-06, 
    1.432992e-06, 1.451313e-06, 1.450296e-06, 1.441993e-06, 1.45041e-06, 
    1.369316e-06, 1.367011e-06, 1.359027e-06, 1.365273e-06, 1.353902e-06, 
    1.360262e-06, 1.363925e-06, 1.378106e-06, 1.38123e-06, 1.384132e-06, 
    1.389872e-06, 1.397255e-06, 1.410257e-06, 1.421618e-06, 1.432029e-06, 
    1.431264e-06, 1.431533e-06, 1.433864e-06, 1.428094e-06, 1.434812e-06, 
    1.435942e-06, 1.43299e-06, 1.45016e-06, 1.445244e-06, 1.450274e-06, 
    1.447072e-06, 1.36776e-06, 1.371639e-06, 1.369542e-06, 1.373487e-06, 
    1.370707e-06, 1.38309e-06, 1.386813e-06, 1.404302e-06, 1.39711e-06, 
    1.408564e-06, 1.398271e-06, 1.400092e-06, 1.40894e-06, 1.398825e-06, 
    1.42099e-06, 1.405945e-06, 1.433955e-06, 1.418863e-06, 1.434903e-06, 
    1.431982e-06, 1.436818e-06, 1.441157e-06, 1.446624e-06, 1.45674e-06, 
    1.454394e-06, 1.462874e-06, 1.377433e-06, 1.382484e-06, 1.382038e-06, 
    1.387333e-06, 1.391256e-06, 1.399777e-06, 1.413499e-06, 1.40833e-06, 
    1.417825e-06, 1.419736e-06, 1.405312e-06, 1.41416e-06, 1.385868e-06, 
    1.39042e-06, 1.387708e-06, 1.377829e-06, 1.40952e-06, 1.393211e-06, 
    1.423401e-06, 1.41451e-06, 1.440538e-06, 1.427564e-06, 1.453103e-06, 
    1.464094e-06, 1.474471e-06, 1.486651e-06, 1.385244e-06, 1.381807e-06, 
    1.387963e-06, 1.396505e-06, 1.404451e-06, 1.415053e-06, 1.41614e-06, 
    1.418131e-06, 1.423295e-06, 1.427645e-06, 1.418761e-06, 1.428736e-06, 
    1.391478e-06, 1.41094e-06, 1.380508e-06, 1.389637e-06, 1.395998e-06, 
    1.393205e-06, 1.407738e-06, 1.411175e-06, 1.425184e-06, 1.417933e-06, 
    1.461378e-06, 1.442074e-06, 1.495955e-06, 1.480797e-06, 1.380607e-06, 
    1.385231e-06, 1.401388e-06, 1.393688e-06, 1.415762e-06, 1.421222e-06, 
    1.425668e-06, 1.431364e-06, 1.431978e-06, 1.435359e-06, 1.429821e-06, 
    1.435139e-06, 1.415074e-06, 1.424023e-06, 1.399533e-06, 1.405474e-06, 
    1.402739e-06, 1.399743e-06, 1.409001e-06, 1.4189e-06, 1.41911e-06, 
    1.422292e-06, 1.43128e-06, 1.415848e-06, 1.46388e-06, 1.434123e-06, 
    1.390283e-06, 1.39923e-06, 1.400508e-06, 1.397038e-06, 1.420674e-06, 
    1.412087e-06, 1.435276e-06, 1.428989e-06, 1.439296e-06, 1.43417e-06, 
    1.433416e-06, 1.426847e-06, 1.422765e-06, 1.412479e-06, 1.404137e-06, 
    1.397539e-06, 1.399071e-06, 1.406323e-06, 1.419505e-06, 1.432032e-06, 
    1.429284e-06, 1.43851e-06, 1.414152e-06, 1.424341e-06, 1.420398e-06, 
    1.430688e-06, 1.408193e-06, 1.427344e-06, 1.403319e-06, 1.405417e-06, 
    1.411916e-06, 1.425036e-06, 1.427945e-06, 1.431057e-06, 1.429136e-06, 
    1.419842e-06, 1.418321e-06, 1.411756e-06, 1.409947e-06, 1.404958e-06, 
    1.400835e-06, 1.404602e-06, 1.408564e-06, 1.419844e-06, 1.430049e-06, 
    1.441217e-06, 1.443957e-06, 1.457077e-06, 1.446393e-06, 1.464046e-06, 
    1.449034e-06, 1.47507e-06, 1.428456e-06, 1.448594e-06, 1.412212e-06, 
    1.416108e-06, 1.423171e-06, 1.439435e-06, 1.430642e-06, 1.440928e-06, 
    1.418261e-06, 1.406575e-06, 1.403557e-06, 1.39794e-06, 1.403686e-06, 
    1.403218e-06, 1.408727e-06, 1.406955e-06, 1.420219e-06, 1.413086e-06, 
    1.433396e-06, 1.440844e-06, 1.461983e-06, 1.475019e-06, 1.488348e-06, 
    1.494252e-06, 1.496051e-06, 1.496804e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  8.662834e-06, 8.70057e-06, 8.69321e-06, 8.72367e-06, 8.706756e-06, 
    8.726694e-06, 8.670432e-06, 8.702013e-06, 8.681835e-06, 8.666148e-06, 
    8.782779e-06, 8.724958e-06, 8.84286e-06, 8.805921e-06, 8.898702e-06, 
    8.837093e-06, 8.911122e-06, 8.896888e-06, 8.939666e-06, 8.927392e-06, 
    8.982162e-06, 8.945302e-06, 9.010546e-06, 8.973335e-06, 8.979147e-06, 
    8.944045e-06, 8.73664e-06, 8.775646e-06, 8.734315e-06, 8.739877e-06, 
    8.737368e-06, 8.707071e-06, 8.691822e-06, 8.659862e-06, 8.665646e-06, 
    8.689109e-06, 8.742311e-06, 8.72422e-06, 8.769762e-06, 8.768734e-06, 
    8.819486e-06, 8.79659e-06, 8.881984e-06, 8.857679e-06, 8.927894e-06, 
    8.910212e-06, 8.927047e-06, 8.921926e-06, 8.927088e-06, 8.901182e-06, 
    8.912261e-06, 8.889468e-06, 8.800986e-06, 8.827021e-06, 8.749374e-06, 
    8.702751e-06, 8.671782e-06, 8.649837e-06, 8.65292e-06, 8.658838e-06, 
    8.689228e-06, 8.717808e-06, 8.73961e-06, 8.75419e-06, 8.76856e-06, 
    8.812151e-06, 8.835201e-06, 8.886883e-06, 8.877536e-06, 8.893343e-06, 
    8.908445e-06, 8.933815e-06, 8.92963e-06, 8.940805e-06, 8.892871e-06, 
    8.924721e-06, 8.872138e-06, 8.886513e-06, 8.772599e-06, 8.729135e-06, 
    8.710707e-06, 8.694545e-06, 8.655299e-06, 8.682394e-06, 8.671701e-06, 
    8.697095e-06, 8.713248e-06, 8.705241e-06, 8.754579e-06, 8.735377e-06, 
    8.836554e-06, 8.792945e-06, 8.906694e-06, 8.879432e-06, 8.9132e-06, 
    8.89596e-06, 8.92549e-06, 8.898897e-06, 8.944949e-06, 8.954992e-06, 
    8.948111e-06, 8.974463e-06, 8.897368e-06, 8.926962e-06, 8.705071e-06, 
    8.706377e-06, 8.712435e-06, 8.685745e-06, 8.684108e-06, 8.659651e-06, 
    8.681385e-06, 8.690653e-06, 8.714158e-06, 8.728067e-06, 8.741292e-06, 
    8.77041e-06, 8.802941e-06, 8.848461e-06, 8.881188e-06, 8.90313e-06, 
    8.88966e-06, 8.901535e-06, 8.888242e-06, 8.881999e-06, 8.951206e-06, 
    8.912332e-06, 8.970645e-06, 8.967417e-06, 8.941002e-06, 8.967755e-06, 
    8.707274e-06, 8.699759e-06, 8.673733e-06, 8.694083e-06, 8.656972e-06, 
    8.677741e-06, 8.689677e-06, 8.735774e-06, 8.74589e-06, 8.755298e-06, 
    8.773858e-06, 8.797693e-06, 8.839557e-06, 8.875995e-06, 8.909285e-06, 
    8.906831e-06, 8.907687e-06, 8.915117e-06, 8.89668e-06, 8.918126e-06, 
    8.921719e-06, 8.9123e-06, 8.966958e-06, 8.951332e-06, 8.967312e-06, 
    8.957121e-06, 8.702186e-06, 8.714794e-06, 8.707962e-06, 8.720792e-06, 
    8.711738e-06, 8.751937e-06, 8.763984e-06, 8.820423e-06, 8.797226e-06, 
    8.834124e-06, 8.800952e-06, 8.806828e-06, 8.835314e-06, 8.802716e-06, 
    8.873964e-06, 8.825647e-06, 8.915396e-06, 8.867121e-06, 8.918405e-06, 
    8.909068e-06, 8.92449e-06, 8.938321e-06, 8.955698e-06, 8.987827e-06, 
    8.980364e-06, 9.007238e-06, 8.733603e-06, 8.749975e-06, 8.748521e-06, 
    8.765656e-06, 8.778333e-06, 8.805837e-06, 8.849977e-06, 8.833353e-06, 
    8.863831e-06, 8.869958e-06, 8.823615e-06, 8.852061e-06, 8.760848e-06, 
    8.775564e-06, 8.766784e-06, 8.734763e-06, 8.837115e-06, 8.784549e-06, 
    8.881623e-06, 8.853106e-06, 8.936324e-06, 8.894925e-06, 8.976263e-06, 
    9.011102e-06, 9.043863e-06, 9.08221e-06, 8.758902e-06, 8.747753e-06, 
    8.767676e-06, 8.795285e-06, 8.820874e-06, 8.854954e-06, 8.858427e-06, 
    8.864802e-06, 8.881335e-06, 8.895256e-06, 8.866808e-06, 8.898719e-06, 
    8.778986e-06, 8.841675e-06, 8.743433e-06, 8.773003e-06, 8.793529e-06, 
    8.78451e-06, 8.831337e-06, 8.842372e-06, 8.887285e-06, 8.864055e-06, 
    9.002481e-06, 8.941187e-06, 9.111393e-06, 9.063778e-06, 8.743854e-06, 
    8.758823e-06, 8.811003e-06, 8.786164e-06, 8.8572e-06, 8.874711e-06, 
    8.888923e-06, 8.907135e-06, 8.909076e-06, 8.91987e-06, 8.902168e-06, 
    8.919152e-06, 8.85493e-06, 8.883611e-06, 8.804927e-06, 8.824055e-06, 
    8.815242e-06, 8.805573e-06, 8.835367e-06, 8.867156e-06, 8.867812e-06, 
    8.877996e-06, 8.906763e-06, 8.857322e-06, 9.010385e-06, 8.915807e-06, 
    8.775157e-06, 8.804041e-06, 8.808143e-06, 8.796951e-06, 8.872929e-06, 
    8.845383e-06, 8.919606e-06, 8.899516e-06, 8.932399e-06, 8.916053e-06, 
    8.913629e-06, 8.89264e-06, 8.87956e-06, 8.846577e-06, 8.819732e-06, 
    8.798467e-06, 8.803391e-06, 8.826757e-06, 8.869071e-06, 8.909148e-06, 
    8.900357e-06, 8.929786e-06, 8.851861e-06, 8.884525e-06, 8.871882e-06, 
    8.904802e-06, 8.832877e-06, 8.894315e-06, 8.817181e-06, 8.823921e-06, 
    8.84481e-06, 8.886885e-06, 8.89616e-06, 8.90611e-06, 8.89995e-06, 
    8.870211e-06, 8.865324e-06, 8.84424e-06, 8.838418e-06, 8.82237e-06, 
    8.809071e-06, 8.821208e-06, 8.833937e-06, 8.870148e-06, 8.902795e-06, 
    8.938409e-06, 8.947123e-06, 8.988802e-06, 8.954871e-06, 9.01087e-06, 
    8.963264e-06, 9.045664e-06, 8.897833e-06, 8.962027e-06, 8.845759e-06, 
    8.858254e-06, 8.880896e-06, 8.932834e-06, 8.904756e-06, 8.937577e-06, 
    8.865126e-06, 8.827584e-06, 8.817852e-06, 8.79975e-06, 8.818249e-06, 
    8.816744e-06, 8.83446e-06, 8.828748e-06, 8.871325e-06, 8.848445e-06, 
    8.913452e-06, 8.937208e-06, 9.004321e-06, 9.045504e-06, 9.087448e-06, 
    9.105968e-06, 9.111606e-06, 9.113955e-06,
  4.951148e-06, 4.988322e-06, 4.981086e-06, 5.011128e-06, 4.994453e-06, 
    5.014138e-06, 4.958675e-06, 4.989801e-06, 4.969922e-06, 4.954488e-06, 
    5.069619e-06, 5.012469e-06, 5.129206e-06, 5.092583e-06, 5.18475e-06, 
    5.123503e-06, 5.197129e-06, 5.182975e-06, 5.225605e-06, 5.21338e-06, 
    5.268048e-06, 5.231251e-06, 5.296456e-06, 5.25925e-06, 5.265066e-06, 
    5.23004e-06, 5.023947e-06, 5.062493e-06, 5.021668e-06, 5.027157e-06, 
    5.024693e-06, 4.994799e-06, 4.979762e-06, 4.948308e-06, 4.954013e-06, 
    4.977115e-06, 5.029626e-06, 5.011776e-06, 5.056797e-06, 5.055779e-06, 
    5.106067e-06, 5.083372e-06, 5.168154e-06, 5.144007e-06, 5.21389e-06, 
    5.196285e-06, 5.213063e-06, 5.207973e-06, 5.213129e-06, 5.187318e-06, 
    5.198372e-06, 5.175677e-06, 5.087621e-06, 5.113446e-06, 5.036561e-06, 
    4.990536e-06, 4.960039e-06, 4.938443e-06, 4.941494e-06, 4.947313e-06, 
    4.97725e-06, 5.005453e-06, 5.026985e-06, 5.041408e-06, 5.055632e-06, 
    5.098786e-06, 5.121669e-06, 5.173044e-06, 5.163755e-06, 5.179491e-06, 
    5.194534e-06, 5.21983e-06, 5.215662e-06, 5.226818e-06, 5.179073e-06, 
    5.210789e-06, 5.158468e-06, 5.172761e-06, 5.059517e-06, 5.016588e-06, 
    4.998394e-06, 4.982477e-06, 4.94384e-06, 4.970511e-06, 4.959992e-06, 
    4.985029e-06, 5.000963e-06, 4.99308e-06, 5.041803e-06, 5.022841e-06, 
    5.123027e-06, 5.079787e-06, 5.192779e-06, 5.165661e-06, 5.199286e-06, 
    5.182118e-06, 5.211547e-06, 5.185058e-06, 5.230971e-06, 5.240989e-06, 
    5.234142e-06, 5.260453e-06, 5.183591e-06, 5.213065e-06, 4.992859e-06, 
    4.994145e-06, 5.000134e-06, 4.973827e-06, 4.972218e-06, 4.948153e-06, 
    4.969563e-06, 4.978692e-06, 5.001887e-06, 5.015627e-06, 5.0287e-06, 
    5.057488e-06, 5.089708e-06, 5.134881e-06, 5.167417e-06, 5.189268e-06, 
    5.175865e-06, 5.187698e-06, 5.174471e-06, 5.168275e-06, 5.237236e-06, 
    5.198476e-06, 5.256666e-06, 5.25344e-06, 5.227084e-06, 5.253803e-06, 
    4.995048e-06, 4.987651e-06, 4.962007e-06, 4.982072e-06, 4.945534e-06, 
    4.965976e-06, 4.977745e-06, 5.02324e-06, 5.033252e-06, 5.042547e-06, 
    5.060919e-06, 5.084533e-06, 5.126051e-06, 5.162271e-06, 5.195409e-06, 
    5.192979e-06, 5.193834e-06, 5.201248e-06, 5.182892e-06, 5.204264e-06, 
    5.207855e-06, 5.198469e-06, 5.253008e-06, 5.237406e-06, 5.253371e-06, 
    5.243211e-06, 4.990055e-06, 5.002504e-06, 4.995775e-06, 5.008431e-06, 
    4.999515e-06, 5.039208e-06, 5.05113e-06, 5.107046e-06, 5.084068e-06, 
    5.120651e-06, 5.087779e-06, 5.093599e-06, 5.121852e-06, 5.089552e-06, 
    5.160274e-06, 5.112295e-06, 5.201537e-06, 5.153497e-06, 5.204553e-06, 
    5.195266e-06, 5.210643e-06, 5.22443e-06, 5.241789e-06, 5.273877e-06, 
    5.26644e-06, 5.293311e-06, 5.021082e-06, 5.037268e-06, 5.03584e-06, 
    5.052795e-06, 5.065348e-06, 5.092591e-06, 5.136394e-06, 5.119906e-06, 
    5.150187e-06, 5.156275e-06, 5.110274e-06, 5.138503e-06, 5.048109e-06, 
    5.062679e-06, 5.054e-06, 5.022359e-06, 5.123708e-06, 5.071608e-06, 
    5.167956e-06, 5.139623e-06, 5.222464e-06, 5.181211e-06, 5.262348e-06, 
    5.297174e-06, 5.330007e-06, 5.368479e-06, 5.046107e-06, 5.0351e-06, 
    5.054812e-06, 5.082135e-06, 5.107524e-06, 5.14135e-06, 5.144814e-06, 
    5.151162e-06, 5.167615e-06, 5.181464e-06, 5.153173e-06, 5.184937e-06, 
    5.066065e-06, 5.128237e-06, 5.030944e-06, 5.060176e-06, 5.080521e-06, 
    5.07159e-06, 5.118022e-06, 5.128988e-06, 5.173636e-06, 5.150537e-06, 
    5.288573e-06, 5.227348e-06, 5.397825e-06, 5.35e-06, 5.031257e-06, 
    5.046068e-06, 5.097738e-06, 5.07313e-06, 5.14361e-06, 5.161012e-06, 
    5.175171e-06, 5.193295e-06, 5.195251e-06, 5.206001e-06, 5.18839e-06, 
    5.205304e-06, 5.141423e-06, 5.169935e-06, 5.091819e-06, 5.110795e-06, 
    5.102062e-06, 5.09249e-06, 5.122052e-06, 5.153619e-06, 5.154289e-06, 
    5.164427e-06, 5.193038e-06, 5.143896e-06, 5.296502e-06, 5.202082e-06, 
    5.062236e-06, 5.090846e-06, 5.094931e-06, 5.08384e-06, 5.159266e-06, 
    5.131892e-06, 5.205738e-06, 5.185743e-06, 5.218518e-06, 5.202223e-06, 
    5.199827e-06, 5.178927e-06, 5.165931e-06, 5.133147e-06, 5.106525e-06, 
    5.085447e-06, 5.090345e-06, 5.113508e-06, 5.15555e-06, 5.195431e-06, 
    5.186686e-06, 5.216024e-06, 5.138488e-06, 5.170954e-06, 5.158398e-06, 
    5.191157e-06, 5.119469e-06, 5.180507e-06, 5.103909e-06, 5.110608e-06, 
    5.131349e-06, 5.173161e-06, 5.182421e-06, 5.192323e-06, 5.186211e-06, 
    5.156618e-06, 5.151774e-06, 5.130844e-06, 5.125072e-06, 5.109149e-06, 
    5.095982e-06, 5.108013e-06, 5.12066e-06, 5.156629e-06, 5.189122e-06, 
    5.224627e-06, 5.233327e-06, 5.274951e-06, 5.241065e-06, 5.297031e-06, 
    5.249446e-06, 5.331905e-06, 5.184045e-06, 5.24804e-06, 5.132292e-06, 
    5.144718e-06, 5.167223e-06, 5.218961e-06, 5.191002e-06, 5.223702e-06, 
    5.151584e-06, 5.114311e-06, 5.104677e-06, 5.086729e-06, 5.105087e-06, 
    5.103593e-06, 5.12118e-06, 5.115526e-06, 5.157825e-06, 5.135088e-06, 
    5.199768e-06, 5.223443e-06, 5.290494e-06, 5.331745e-06, 5.373839e-06, 
    5.392461e-06, 5.398133e-06, 5.400505e-06,
  4.464231e-06, 4.503533e-06, 4.495881e-06, 4.527663e-06, 4.51002e-06, 
    4.530849e-06, 4.472186e-06, 4.505097e-06, 4.484075e-06, 4.467761e-06, 
    4.589611e-06, 4.529083e-06, 4.652822e-06, 4.613964e-06, 4.711826e-06, 
    4.646768e-06, 4.724988e-06, 4.709941e-06, 4.755282e-06, 4.742274e-06, 
    4.800466e-06, 4.76129e-06, 4.83074e-06, 4.791097e-06, 4.797291e-06, 
    4.76e-06, 4.541234e-06, 4.582058e-06, 4.538821e-06, 4.544632e-06, 
    4.542024e-06, 4.510385e-06, 4.494478e-06, 4.461231e-06, 4.467259e-06, 
    4.491681e-06, 4.547246e-06, 4.52835e-06, 4.576028e-06, 4.574949e-06, 
    4.628268e-06, 4.604196e-06, 4.69419e-06, 4.668538e-06, 4.742817e-06, 
    4.724092e-06, 4.741937e-06, 4.736522e-06, 4.742007e-06, 4.714557e-06, 
    4.726311e-06, 4.702184e-06, 4.608701e-06, 4.636096e-06, 4.55459e-06, 
    4.505873e-06, 4.473628e-06, 4.450807e-06, 4.454031e-06, 4.460178e-06, 
    4.491824e-06, 4.521659e-06, 4.544452e-06, 4.559725e-06, 4.574794e-06, 
    4.62054e-06, 4.644822e-06, 4.699385e-06, 4.689516e-06, 4.706237e-06, 
    4.722231e-06, 4.749135e-06, 4.744702e-06, 4.756571e-06, 4.705794e-06, 
    4.739517e-06, 4.683899e-06, 4.699085e-06, 4.578904e-06, 4.533444e-06, 
    4.514187e-06, 4.497351e-06, 4.456509e-06, 4.484698e-06, 4.473578e-06, 
    4.500051e-06, 4.516908e-06, 4.508567e-06, 4.560143e-06, 4.540063e-06, 
    4.646263e-06, 4.600395e-06, 4.720364e-06, 4.691541e-06, 4.727283e-06, 
    4.70903e-06, 4.740324e-06, 4.712156e-06, 4.760991e-06, 4.771653e-06, 
    4.764366e-06, 4.792379e-06, 4.710597e-06, 4.741938e-06, 4.508334e-06, 
    4.509694e-06, 4.516031e-06, 4.488204e-06, 4.486503e-06, 4.461066e-06, 
    4.483696e-06, 4.493348e-06, 4.517885e-06, 4.532426e-06, 4.546267e-06, 
    4.57676e-06, 4.610914e-06, 4.658847e-06, 4.693407e-06, 4.716632e-06, 
    4.702385e-06, 4.714962e-06, 4.700903e-06, 4.694319e-06, 4.767658e-06, 
    4.726421e-06, 4.788346e-06, 4.78491e-06, 4.756854e-06, 4.785297e-06, 
    4.510649e-06, 4.502825e-06, 4.475708e-06, 4.496924e-06, 4.4583e-06, 
    4.479904e-06, 4.492346e-06, 4.540484e-06, 4.551087e-06, 4.560931e-06, 
    4.580396e-06, 4.605427e-06, 4.649474e-06, 4.687938e-06, 4.723161e-06, 
    4.720577e-06, 4.721487e-06, 4.72937e-06, 4.709853e-06, 4.732577e-06, 
    4.736396e-06, 4.726415e-06, 4.784451e-06, 4.76784e-06, 4.784838e-06, 
    4.774019e-06, 4.505367e-06, 4.518538e-06, 4.511419e-06, 4.52481e-06, 
    4.515375e-06, 4.557393e-06, 4.570022e-06, 4.629305e-06, 4.604934e-06, 
    4.643742e-06, 4.608869e-06, 4.615041e-06, 4.645015e-06, 4.610751e-06, 
    4.685815e-06, 4.634873e-06, 4.729677e-06, 4.678614e-06, 4.732884e-06, 
    4.723009e-06, 4.739362e-06, 4.75403e-06, 4.772506e-06, 4.806678e-06, 
    4.798756e-06, 4.827387e-06, 4.538201e-06, 4.555339e-06, 4.553828e-06, 
    4.571788e-06, 4.58509e-06, 4.613973e-06, 4.660455e-06, 4.642952e-06, 
    4.675102e-06, 4.681568e-06, 4.632731e-06, 4.662693e-06, 4.566823e-06, 
    4.582258e-06, 4.573064e-06, 4.539553e-06, 4.646986e-06, 4.591723e-06, 
    4.693979e-06, 4.663883e-06, 4.751938e-06, 4.708065e-06, 4.794397e-06, 
    4.831502e-06, 4.86652e-06, 4.907582e-06, 4.564702e-06, 4.553044e-06, 
    4.573925e-06, 4.602883e-06, 4.629812e-06, 4.665717e-06, 4.669396e-06, 
    4.676138e-06, 4.693617e-06, 4.708335e-06, 4.678272e-06, 4.712027e-06, 
    4.585845e-06, 4.651795e-06, 4.548642e-06, 4.579606e-06, 4.601173e-06, 
    4.591705e-06, 4.640953e-06, 4.652592e-06, 4.700014e-06, 4.675474e-06, 
    4.822336e-06, 4.757133e-06, 4.938933e-06, 4.887854e-06, 4.548975e-06, 
    4.564661e-06, 4.619431e-06, 4.593338e-06, 4.668118e-06, 4.686601e-06, 
    4.701647e-06, 4.720912e-06, 4.722993e-06, 4.734424e-06, 4.715698e-06, 
    4.733683e-06, 4.665794e-06, 4.696083e-06, 4.613155e-06, 4.633284e-06, 
    4.624019e-06, 4.613866e-06, 4.645231e-06, 4.678746e-06, 4.67946e-06, 
    4.690228e-06, 4.720634e-06, 4.668421e-06, 4.830783e-06, 4.730251e-06, 
    4.581792e-06, 4.61212e-06, 4.616455e-06, 4.604693e-06, 4.684747e-06, 
    4.655675e-06, 4.734145e-06, 4.712884e-06, 4.74774e-06, 4.730407e-06, 
    4.727859e-06, 4.705639e-06, 4.691828e-06, 4.657007e-06, 4.628753e-06, 
    4.606397e-06, 4.611592e-06, 4.636163e-06, 4.680798e-06, 4.723183e-06, 
    4.713885e-06, 4.745087e-06, 4.662678e-06, 4.697164e-06, 4.683824e-06, 
    4.718639e-06, 4.642488e-06, 4.707313e-06, 4.625979e-06, 4.633086e-06, 
    4.655099e-06, 4.699509e-06, 4.709353e-06, 4.719878e-06, 4.713382e-06, 
    4.681933e-06, 4.676788e-06, 4.654562e-06, 4.648436e-06, 4.631538e-06, 
    4.617569e-06, 4.630332e-06, 4.643752e-06, 4.681945e-06, 4.716475e-06, 
    4.754239e-06, 4.763498e-06, 4.807819e-06, 4.771732e-06, 4.831346e-06, 
    4.78065e-06, 4.868541e-06, 4.711075e-06, 4.779156e-06, 4.6561e-06, 
    4.669294e-06, 4.693199e-06, 4.748209e-06, 4.718475e-06, 4.753254e-06, 
    4.676586e-06, 4.637013e-06, 4.626793e-06, 4.607756e-06, 4.627228e-06, 
    4.625643e-06, 4.644306e-06, 4.638305e-06, 4.683215e-06, 4.659069e-06, 
    4.727795e-06, 4.752978e-06, 4.824385e-06, 4.868373e-06, 4.91331e-06, 
    4.933202e-06, 4.939263e-06, 4.941798e-06,
  4.33327e-06, 4.374281e-06, 4.366293e-06, 4.399478e-06, 4.381054e-06, 
    4.402805e-06, 4.341568e-06, 4.375914e-06, 4.353973e-06, 4.336952e-06, 
    4.46422e-06, 4.40096e-06, 4.530367e-06, 4.489693e-06, 4.592192e-06, 
    4.524029e-06, 4.605994e-06, 4.590215e-06, 4.637773e-06, 4.624125e-06, 
    4.685212e-06, 4.644078e-06, 4.717022e-06, 4.675372e-06, 4.681877e-06, 
    4.642725e-06, 4.413654e-06, 4.456323e-06, 4.411133e-06, 4.417203e-06, 
    4.414478e-06, 4.381435e-06, 4.36483e-06, 4.330141e-06, 4.336428e-06, 
    4.36191e-06, 4.419934e-06, 4.400194e-06, 4.450017e-06, 4.448888e-06, 
    4.504662e-06, 4.479474e-06, 4.573704e-06, 4.546827e-06, 4.624694e-06, 
    4.605053e-06, 4.623771e-06, 4.618091e-06, 4.623845e-06, 4.595056e-06, 
    4.607381e-06, 4.582084e-06, 4.484187e-06, 4.512856e-06, 4.427608e-06, 
    4.376724e-06, 4.343072e-06, 4.31927e-06, 4.322631e-06, 4.329043e-06, 
    4.362059e-06, 4.393206e-06, 4.417015e-06, 4.432974e-06, 4.448726e-06, 
    4.496575e-06, 4.521991e-06, 4.57915e-06, 4.568806e-06, 4.586333e-06, 
    4.603101e-06, 4.631323e-06, 4.626672e-06, 4.639127e-06, 4.585868e-06, 
    4.621233e-06, 4.56292e-06, 4.578835e-06, 4.453025e-06, 4.405515e-06, 
    4.385405e-06, 4.367828e-06, 4.325217e-06, 4.354623e-06, 4.34302e-06, 
    4.370646e-06, 4.388245e-06, 4.379536e-06, 4.433412e-06, 4.412429e-06, 
    4.5235e-06, 4.475498e-06, 4.601144e-06, 4.570928e-06, 4.6084e-06, 
    4.58926e-06, 4.622079e-06, 4.592538e-06, 4.643765e-06, 4.654957e-06, 
    4.647307e-06, 4.676718e-06, 4.590903e-06, 4.623772e-06, 4.379293e-06, 
    4.380713e-06, 4.387329e-06, 4.358281e-06, 4.356506e-06, 4.329969e-06, 
    4.353577e-06, 4.36365e-06, 4.389266e-06, 4.404452e-06, 4.418911e-06, 
    4.450781e-06, 4.486503e-06, 4.536677e-06, 4.572884e-06, 4.597231e-06, 
    4.582294e-06, 4.59548e-06, 4.580741e-06, 4.57384e-06, 4.650763e-06, 
    4.607496e-06, 4.672483e-06, 4.668875e-06, 4.639423e-06, 4.669282e-06, 
    4.38171e-06, 4.373542e-06, 4.345242e-06, 4.367382e-06, 4.327083e-06, 
    4.34962e-06, 4.362604e-06, 4.41287e-06, 4.423948e-06, 4.434235e-06, 
    4.454583e-06, 4.480762e-06, 4.526862e-06, 4.567152e-06, 4.604077e-06, 
    4.601367e-06, 4.602321e-06, 4.610589e-06, 4.590124e-06, 4.613953e-06, 
    4.617959e-06, 4.60749e-06, 4.668392e-06, 4.650954e-06, 4.668798e-06, 
    4.65744e-06, 4.376196e-06, 4.389947e-06, 4.382514e-06, 4.396497e-06, 
    4.386644e-06, 4.430538e-06, 4.443738e-06, 4.505748e-06, 4.480246e-06, 
    4.52086e-06, 4.484363e-06, 4.490821e-06, 4.522193e-06, 4.486331e-06, 
    4.564929e-06, 4.511576e-06, 4.61091e-06, 4.557384e-06, 4.614275e-06, 
    4.603917e-06, 4.62107e-06, 4.636459e-06, 4.655852e-06, 4.691737e-06, 
    4.683415e-06, 4.713498e-06, 4.410485e-06, 4.428392e-06, 4.426811e-06, 
    4.445583e-06, 4.459491e-06, 4.489702e-06, 4.538361e-06, 4.520033e-06, 
    4.553704e-06, 4.560478e-06, 4.509334e-06, 4.540706e-06, 4.440393e-06, 
    4.456531e-06, 4.446918e-06, 4.411897e-06, 4.524257e-06, 4.466428e-06, 
    4.573484e-06, 4.541952e-06, 4.634264e-06, 4.588249e-06, 4.678838e-06, 
    4.717824e-06, 4.754643e-06, 4.797853e-06, 4.438177e-06, 4.425993e-06, 
    4.447817e-06, 4.4781e-06, 4.506279e-06, 4.543873e-06, 4.547726e-06, 
    4.554789e-06, 4.573104e-06, 4.588532e-06, 4.557025e-06, 4.592403e-06, 
    4.460282e-06, 4.529292e-06, 4.421393e-06, 4.453757e-06, 4.476312e-06, 
    4.466409e-06, 4.51794e-06, 4.530127e-06, 4.579809e-06, 4.554093e-06, 
    4.708189e-06, 4.639716e-06, 4.830869e-06, 4.777088e-06, 4.42174e-06, 
    4.438134e-06, 4.495414e-06, 4.468117e-06, 4.546387e-06, 4.565752e-06, 
    4.581521e-06, 4.601719e-06, 4.603901e-06, 4.615891e-06, 4.596251e-06, 
    4.615113e-06, 4.543953e-06, 4.575688e-06, 4.488847e-06, 4.509913e-06, 
    4.500215e-06, 4.489591e-06, 4.522419e-06, 4.557521e-06, 4.558269e-06, 
    4.569553e-06, 4.601428e-06, 4.546705e-06, 4.717069e-06, 4.611515e-06, 
    4.456042e-06, 4.487765e-06, 4.4923e-06, 4.479994e-06, 4.563808e-06, 
    4.533355e-06, 4.615598e-06, 4.593301e-06, 4.629859e-06, 4.611676e-06, 
    4.609004e-06, 4.585705e-06, 4.571229e-06, 4.53475e-06, 4.50517e-06, 
    4.481777e-06, 4.487211e-06, 4.512926e-06, 4.559672e-06, 4.6041e-06, 
    4.594351e-06, 4.627076e-06, 4.54069e-06, 4.576822e-06, 4.562842e-06, 
    4.599336e-06, 4.519547e-06, 4.587461e-06, 4.502266e-06, 4.509705e-06, 
    4.532752e-06, 4.57928e-06, 4.589599e-06, 4.600635e-06, 4.593823e-06, 
    4.560861e-06, 4.555469e-06, 4.53219e-06, 4.525774e-06, 4.508085e-06, 
    4.493465e-06, 4.506822e-06, 4.52087e-06, 4.560873e-06, 4.597066e-06, 
    4.636679e-06, 4.646396e-06, 4.692937e-06, 4.655039e-06, 4.71766e-06, 
    4.664404e-06, 4.756769e-06, 4.591406e-06, 4.662834e-06, 4.533801e-06, 
    4.547619e-06, 4.572667e-06, 4.630352e-06, 4.599163e-06, 4.635646e-06, 
    4.555258e-06, 4.513816e-06, 4.503118e-06, 4.483198e-06, 4.503574e-06, 
    4.501915e-06, 4.52145e-06, 4.515168e-06, 4.562204e-06, 4.53691e-06, 
    4.608938e-06, 4.635357e-06, 4.710342e-06, 4.756592e-06, 4.803882e-06, 
    4.824832e-06, 4.831216e-06, 4.833886e-06,
  4.365276e-06, 4.405923e-06, 4.398003e-06, 4.430912e-06, 4.412638e-06, 
    4.434213e-06, 4.373498e-06, 4.407543e-06, 4.385791e-06, 4.368924e-06, 
    4.495179e-06, 4.432383e-06, 4.560924e-06, 4.520485e-06, 4.622454e-06, 
    4.55462e-06, 4.6362e-06, 4.620485e-06, 4.667867e-06, 4.654264e-06, 
    4.715183e-06, 4.674153e-06, 4.746933e-06, 4.705363e-06, 4.711854e-06, 
    4.672804e-06, 4.444976e-06, 4.487335e-06, 4.442474e-06, 4.448499e-06, 
    4.445794e-06, 4.413017e-06, 4.396554e-06, 4.362175e-06, 4.368404e-06, 
    4.393658e-06, 4.451209e-06, 4.431623e-06, 4.48107e-06, 4.47995e-06, 
    4.535363e-06, 4.510331e-06, 4.604045e-06, 4.577297e-06, 4.654832e-06, 
    4.635263e-06, 4.653912e-06, 4.648252e-06, 4.653986e-06, 4.625305e-06, 
    4.637581e-06, 4.612388e-06, 4.515014e-06, 4.543509e-06, 4.458825e-06, 
    4.408347e-06, 4.374988e-06, 4.351407e-06, 4.354737e-06, 4.361088e-06, 
    4.393806e-06, 4.424691e-06, 4.44831e-06, 4.464151e-06, 4.479789e-06, 
    4.527327e-06, 4.552594e-06, 4.609467e-06, 4.599169e-06, 4.616619e-06, 
    4.633318e-06, 4.661439e-06, 4.656803e-06, 4.669217e-06, 4.616155e-06, 
    4.651383e-06, 4.59331e-06, 4.609153e-06, 4.484061e-06, 4.436901e-06, 
    4.416954e-06, 4.399526e-06, 4.357298e-06, 4.386436e-06, 4.374936e-06, 
    4.402319e-06, 4.41977e-06, 4.411133e-06, 4.464584e-06, 4.443761e-06, 
    4.554094e-06, 4.50638e-06, 4.631369e-06, 4.601281e-06, 4.638597e-06, 
    4.619533e-06, 4.652226e-06, 4.622797e-06, 4.673841e-06, 4.685e-06, 
    4.677373e-06, 4.706706e-06, 4.621169e-06, 4.653913e-06, 4.410892e-06, 
    4.4123e-06, 4.418861e-06, 4.390061e-06, 4.388302e-06, 4.362005e-06, 
    4.385399e-06, 4.395383e-06, 4.420782e-06, 4.435847e-06, 4.450193e-06, 
    4.48183e-06, 4.517315e-06, 4.5672e-06, 4.603229e-06, 4.627471e-06, 
    4.612596e-06, 4.625727e-06, 4.61105e-06, 4.60418e-06, 4.680818e-06, 
    4.637696e-06, 4.70248e-06, 4.698881e-06, 4.669513e-06, 4.699287e-06, 
    4.413288e-06, 4.405189e-06, 4.377139e-06, 4.399082e-06, 4.359147e-06, 
    4.381477e-06, 4.394347e-06, 4.444199e-06, 4.455191e-06, 4.465402e-06, 
    4.485605e-06, 4.51161e-06, 4.557437e-06, 4.597523e-06, 4.63429e-06, 
    4.63159e-06, 4.632541e-06, 4.640777e-06, 4.620393e-06, 4.644129e-06, 
    4.64812e-06, 4.637689e-06, 4.6984e-06, 4.681009e-06, 4.698805e-06, 
    4.687476e-06, 4.407821e-06, 4.421458e-06, 4.414086e-06, 4.427955e-06, 
    4.418183e-06, 4.461733e-06, 4.474837e-06, 4.536443e-06, 4.511098e-06, 
    4.551468e-06, 4.515188e-06, 4.521606e-06, 4.552795e-06, 4.517144e-06, 
    4.595311e-06, 4.542238e-06, 4.641098e-06, 4.587803e-06, 4.644449e-06, 
    4.634131e-06, 4.65122e-06, 4.666559e-06, 4.685893e-06, 4.721692e-06, 
    4.713388e-06, 4.743414e-06, 4.441831e-06, 4.459602e-06, 4.458033e-06, 
    4.476668e-06, 4.49048e-06, 4.520494e-06, 4.568874e-06, 4.550645e-06, 
    4.584138e-06, 4.590881e-06, 4.540007e-06, 4.571207e-06, 4.471516e-06, 
    4.487541e-06, 4.477994e-06, 4.443233e-06, 4.554846e-06, 4.497371e-06, 
    4.603826e-06, 4.572446e-06, 4.66437e-06, 4.618527e-06, 4.708821e-06, 
    4.747735e-06, 4.784514e-06, 4.827719e-06, 4.469315e-06, 4.457221e-06, 
    4.478887e-06, 4.508966e-06, 4.53697e-06, 4.574357e-06, 4.578191e-06, 
    4.585218e-06, 4.603448e-06, 4.618808e-06, 4.587445e-06, 4.622663e-06, 
    4.491267e-06, 4.559854e-06, 4.452656e-06, 4.484787e-06, 4.507189e-06, 
    4.497351e-06, 4.548564e-06, 4.560683e-06, 4.610123e-06, 4.584526e-06, 
    4.738116e-06, 4.669806e-06, 4.860757e-06, 4.806951e-06, 4.453e-06, 
    4.469272e-06, 4.526171e-06, 4.499047e-06, 4.576858e-06, 4.596129e-06, 
    4.611827e-06, 4.631942e-06, 4.634115e-06, 4.64606e-06, 4.626495e-06, 
    4.645285e-06, 4.574437e-06, 4.60602e-06, 4.519643e-06, 4.540583e-06, 
    4.530942e-06, 4.520383e-06, 4.553018e-06, 4.587938e-06, 4.588681e-06, 
    4.599913e-06, 4.631655e-06, 4.577174e-06, 4.746983e-06, 4.641703e-06, 
    4.487054e-06, 4.518569e-06, 4.523075e-06, 4.510846e-06, 4.594195e-06, 
    4.563894e-06, 4.645768e-06, 4.623557e-06, 4.659979e-06, 4.64186e-06, 
    4.639198e-06, 4.615993e-06, 4.601581e-06, 4.565282e-06, 4.535868e-06, 
    4.512618e-06, 4.518018e-06, 4.543579e-06, 4.590078e-06, 4.634314e-06, 
    4.624604e-06, 4.657205e-06, 4.57119e-06, 4.607149e-06, 4.593233e-06, 
    4.629567e-06, 4.550162e-06, 4.617745e-06, 4.532981e-06, 4.540376e-06, 
    4.563294e-06, 4.609597e-06, 4.61987e-06, 4.630862e-06, 4.624077e-06, 
    4.591261e-06, 4.585896e-06, 4.562735e-06, 4.556355e-06, 4.538765e-06, 
    4.524234e-06, 4.53751e-06, 4.551478e-06, 4.591273e-06, 4.627308e-06, 
    4.666778e-06, 4.676464e-06, 4.722892e-06, 4.685084e-06, 4.747574e-06, 
    4.694426e-06, 4.786642e-06, 4.621671e-06, 4.692859e-06, 4.564337e-06, 
    4.578084e-06, 4.603013e-06, 4.660472e-06, 4.629396e-06, 4.665748e-06, 
    4.585685e-06, 4.544464e-06, 4.533828e-06, 4.51403e-06, 4.534281e-06, 
    4.532632e-06, 4.552054e-06, 4.545807e-06, 4.592598e-06, 4.56743e-06, 
    4.639133e-06, 4.66546e-06, 4.740264e-06, 4.786463e-06, 4.833749e-06, 
    4.854713e-06, 4.861104e-06, 4.863777e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 SNOW_SOURCES =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 SOIL1C =
  5.777962, 5.777942, 5.777946, 5.777929, 5.777938, 5.777928, 5.777958, 
    5.777941, 5.777952, 5.77796, 5.777898, 5.777929, 5.777866, 5.777885, 
    5.777836, 5.777869, 5.77783, 5.777837, 5.777814, 5.777821, 5.777792, 
    5.777811, 5.777777, 5.777796, 5.777793, 5.777812, 5.777923, 5.777902, 
    5.777924, 5.777921, 5.777922, 5.777938, 5.777946, 5.777964, 5.77796, 
    5.777948, 5.777919, 5.777929, 5.777905, 5.777905, 5.777878, 5.777891, 
    5.777845, 5.777858, 5.777821, 5.77783, 5.777821, 5.777823, 5.777821, 
    5.777835, 5.777829, 5.777841, 5.777888, 5.777874, 5.777916, 5.777941, 
    5.777957, 5.777969, 5.777967, 5.777964, 5.777948, 5.777933, 5.777921, 
    5.777913, 5.777905, 5.777882, 5.77787, 5.777843, 5.777847, 5.777839, 
    5.777831, 5.777817, 5.77782, 5.777813, 5.777839, 5.777822, 5.77785, 
    5.777843, 5.777904, 5.777926, 5.777936, 5.777945, 5.777966, 5.777952, 
    5.777957, 5.777944, 5.777935, 5.777939, 5.777913, 5.777923, 5.777869, 
    5.777893, 5.777832, 5.777846, 5.777828, 5.777837, 5.777822, 5.777836, 
    5.777812, 5.777806, 5.77781, 5.777796, 5.777837, 5.777821, 5.777939, 
    5.777939, 5.777936, 5.77795, 5.777951, 5.777964, 5.777952, 5.777947, 
    5.777935, 5.777927, 5.77792, 5.777905, 5.777887, 5.777863, 5.777845, 
    5.777833, 5.777841, 5.777834, 5.777842, 5.777845, 5.777808, 5.777829, 
    5.777798, 5.7778, 5.777813, 5.777799, 5.777938, 5.777942, 5.777956, 
    5.777945, 5.777965, 5.777954, 5.777947, 5.777923, 5.777917, 5.777913, 
    5.777903, 5.77789, 5.777867, 5.777848, 5.777831, 5.777832, 5.777831, 
    5.777827, 5.777837, 5.777826, 5.777824, 5.777829, 5.7778, 5.777808, 
    5.7778, 5.777805, 5.777941, 5.777934, 5.777938, 5.777931, 5.777936, 
    5.777915, 5.777908, 5.777878, 5.77789, 5.777871, 5.777888, 5.777885, 
    5.77787, 5.777887, 5.777849, 5.777875, 5.777827, 5.777853, 5.777825, 
    5.777831, 5.777822, 5.777815, 5.777806, 5.777789, 5.777792, 5.777778, 
    5.777924, 5.777915, 5.777916, 5.777907, 5.7779, 5.777885, 5.777862, 
    5.777871, 5.777854, 5.777851, 5.777876, 5.777861, 5.777909, 5.777902, 
    5.777906, 5.777924, 5.777869, 5.777897, 5.777845, 5.77786, 5.777816, 
    5.777838, 5.777795, 5.777776, 5.777759, 5.777739, 5.777911, 5.777916, 
    5.777906, 5.777891, 5.777877, 5.777859, 5.777857, 5.777854, 5.777845, 
    5.777838, 5.777853, 5.777836, 5.7779, 5.777866, 5.777919, 5.777903, 
    5.777892, 5.777897, 5.777872, 5.777866, 5.777842, 5.777854, 5.777781, 
    5.777813, 5.777723, 5.777748, 5.777919, 5.777911, 5.777883, 5.777896, 
    5.777858, 5.777849, 5.777841, 5.777832, 5.777831, 5.777825, 5.777834, 
    5.777825, 5.777859, 5.777844, 5.777886, 5.777876, 5.77788, 5.777885, 
    5.77787, 5.777853, 5.777853, 5.777847, 5.777832, 5.777858, 5.777777, 
    5.777827, 5.777902, 5.777886, 5.777884, 5.77789, 5.77785, 5.777864, 
    5.777825, 5.777835, 5.777818, 5.777827, 5.777828, 5.777839, 5.777846, 
    5.777864, 5.777878, 5.777889, 5.777887, 5.777874, 5.777852, 5.777831, 
    5.777835, 5.777819, 5.777861, 5.777843, 5.77785, 5.777833, 5.777871, 
    5.777838, 5.777879, 5.777876, 5.777864, 5.777842, 5.777837, 5.777832, 
    5.777835, 5.777851, 5.777853, 5.777865, 5.777868, 5.777876, 5.777884, 
    5.777877, 5.777871, 5.777851, 5.777834, 5.777815, 5.77781, 5.777788, 
    5.777806, 5.777776, 5.777802, 5.777758, 5.777836, 5.777802, 5.777864, 
    5.777857, 5.777845, 5.777818, 5.777833, 5.777815, 5.777854, 5.777874, 
    5.777879, 5.777889, 5.777879, 5.77788, 5.77787, 5.777873, 5.777851, 
    5.777863, 5.777828, 5.777815, 5.77778, 5.777758, 5.777736, 5.777726, 
    5.777723, 5.777721 ;

 SOIL1C_TO_SOIL2C =
  3.181218e-08, 3.195197e-08, 3.192479e-08, 3.203753e-08, 3.197499e-08, 
    3.204882e-08, 3.184052e-08, 3.195752e-08, 3.188283e-08, 3.182477e-08, 
    3.225633e-08, 3.204256e-08, 3.247835e-08, 3.234203e-08, 3.268446e-08, 
    3.245713e-08, 3.273029e-08, 3.26779e-08, 3.283559e-08, 3.279041e-08, 
    3.299211e-08, 3.285644e-08, 3.309666e-08, 3.295971e-08, 3.298113e-08, 
    3.285196e-08, 3.208558e-08, 3.222972e-08, 3.207704e-08, 3.209759e-08, 
    3.208837e-08, 3.197628e-08, 3.19198e-08, 3.180149e-08, 3.182297e-08, 
    3.190986e-08, 3.210684e-08, 3.203997e-08, 3.220848e-08, 3.220467e-08, 
    3.239226e-08, 3.230768e-08, 3.262297e-08, 3.253336e-08, 3.27923e-08, 
    3.272718e-08, 3.278924e-08, 3.277042e-08, 3.278948e-08, 3.269398e-08, 
    3.27349e-08, 3.265086e-08, 3.232352e-08, 3.241973e-08, 3.21328e-08, 
    3.196026e-08, 3.184565e-08, 3.176433e-08, 3.177582e-08, 3.179774e-08, 
    3.191037e-08, 3.201626e-08, 3.209696e-08, 3.215094e-08, 3.220412e-08, 
    3.236512e-08, 3.245032e-08, 3.264109e-08, 3.260666e-08, 3.266499e-08, 
    3.27207e-08, 3.281425e-08, 3.279885e-08, 3.284006e-08, 3.266344e-08, 
    3.278083e-08, 3.258705e-08, 3.264005e-08, 3.22186e-08, 3.205801e-08, 
    3.198976e-08, 3.193001e-08, 3.178466e-08, 3.188504e-08, 3.184547e-08, 
    3.193961e-08, 3.199942e-08, 3.196984e-08, 3.215241e-08, 3.208143e-08, 
    3.245537e-08, 3.229431e-08, 3.27142e-08, 3.261373e-08, 3.273828e-08, 
    3.267472e-08, 3.278363e-08, 3.268562e-08, 3.28554e-08, 3.289237e-08, 
    3.286711e-08, 3.296415e-08, 3.268018e-08, 3.278924e-08, 3.196901e-08, 
    3.197383e-08, 3.199631e-08, 3.189751e-08, 3.189146e-08, 3.180091e-08, 
    3.188148e-08, 3.191579e-08, 3.200289e-08, 3.205441e-08, 3.210338e-08, 
    3.221105e-08, 3.23313e-08, 3.249945e-08, 3.262024e-08, 3.270121e-08, 
    3.265156e-08, 3.269539e-08, 3.264639e-08, 3.262342e-08, 3.287852e-08, 
    3.273528e-08, 3.295019e-08, 3.29383e-08, 3.284104e-08, 3.293964e-08, 
    3.197722e-08, 3.194945e-08, 3.185306e-08, 3.19285e-08, 3.179105e-08, 
    3.186799e-08, 3.191223e-08, 3.208292e-08, 3.212042e-08, 3.21552e-08, 
    3.222387e-08, 3.231201e-08, 3.246663e-08, 3.260114e-08, 3.272394e-08, 
    3.271494e-08, 3.271811e-08, 3.274554e-08, 3.267759e-08, 3.27567e-08, 
    3.276998e-08, 3.273526e-08, 3.293671e-08, 3.287916e-08, 3.293805e-08, 
    3.290058e-08, 3.195848e-08, 3.20052e-08, 3.197995e-08, 3.202743e-08, 
    3.199398e-08, 3.214269e-08, 3.218728e-08, 3.23959e-08, 3.231028e-08, 
    3.244654e-08, 3.232412e-08, 3.234581e-08, 3.245099e-08, 3.233073e-08, 
    3.259373e-08, 3.241543e-08, 3.274661e-08, 3.256857e-08, 3.275777e-08, 
    3.272341e-08, 3.278029e-08, 3.283124e-08, 3.289533e-08, 3.301359e-08, 
    3.29862e-08, 3.30851e-08, 3.207485e-08, 3.213544e-08, 3.213011e-08, 
    3.219352e-08, 3.224041e-08, 3.234206e-08, 3.250507e-08, 3.244377e-08, 
    3.255631e-08, 3.25789e-08, 3.240793e-08, 3.251291e-08, 3.2176e-08, 
    3.223044e-08, 3.219802e-08, 3.207963e-08, 3.24579e-08, 3.226378e-08, 
    3.262224e-08, 3.251708e-08, 3.282398e-08, 3.267136e-08, 3.297113e-08, 
    3.309929e-08, 3.321988e-08, 3.336083e-08, 3.216851e-08, 3.212734e-08, 
    3.220106e-08, 3.230306e-08, 3.239769e-08, 3.252349e-08, 3.253636e-08, 
    3.255993e-08, 3.262097e-08, 3.26723e-08, 3.256739e-08, 3.268517e-08, 
    3.224307e-08, 3.247475e-08, 3.211177e-08, 3.222108e-08, 3.229704e-08, 
    3.226372e-08, 3.243677e-08, 3.247755e-08, 3.264329e-08, 3.255761e-08, 
    3.306766e-08, 3.284201e-08, 3.346814e-08, 3.329317e-08, 3.211295e-08, 
    3.216837e-08, 3.236123e-08, 3.226947e-08, 3.253189e-08, 3.259648e-08, 
    3.264899e-08, 3.271611e-08, 3.272335e-08, 3.276312e-08, 3.269795e-08, 
    3.276055e-08, 3.252376e-08, 3.262958e-08, 3.233918e-08, 3.240987e-08, 
    3.237735e-08, 3.234168e-08, 3.245176e-08, 3.256904e-08, 3.257154e-08, 
    3.260914e-08, 3.271512e-08, 3.253295e-08, 3.309679e-08, 3.274859e-08, 
    3.22288e-08, 3.233554e-08, 3.235078e-08, 3.230943e-08, 3.259001e-08, 
    3.248834e-08, 3.276215e-08, 3.268815e-08, 3.28094e-08, 3.274915e-08, 
    3.274029e-08, 3.26629e-08, 3.261473e-08, 3.249301e-08, 3.239397e-08, 
    3.231543e-08, 3.233369e-08, 3.241997e-08, 3.257621e-08, 3.272401e-08, 
    3.269164e-08, 3.280018e-08, 3.251286e-08, 3.263334e-08, 3.258678e-08, 
    3.27082e-08, 3.244214e-08, 3.266872e-08, 3.238423e-08, 3.240917e-08, 
    3.248633e-08, 3.264152e-08, 3.267585e-08, 3.271251e-08, 3.268989e-08, 
    3.258018e-08, 3.25622e-08, 3.248445e-08, 3.246299e-08, 3.240374e-08, 
    3.235469e-08, 3.239951e-08, 3.244657e-08, 3.258022e-08, 3.270066e-08, 
    3.283197e-08, 3.28641e-08, 3.301752e-08, 3.289264e-08, 3.309873e-08, 
    3.292352e-08, 3.322681e-08, 3.268184e-08, 3.291836e-08, 3.248984e-08, 
    3.2536e-08, 3.261951e-08, 3.281102e-08, 3.270763e-08, 3.282854e-08, 
    3.256149e-08, 3.242294e-08, 3.238709e-08, 3.23202e-08, 3.238862e-08, 
    3.238305e-08, 3.244852e-08, 3.242748e-08, 3.258465e-08, 3.250023e-08, 
    3.274006e-08, 3.282759e-08, 3.307474e-08, 3.322625e-08, 3.338046e-08, 
    3.344855e-08, 3.346927e-08, 3.347793e-08 ;

 SOIL1C_TO_SOIL3C =
  3.773021e-10, 3.789605e-10, 3.786381e-10, 3.799758e-10, 3.792337e-10, 
    3.801096e-10, 3.776383e-10, 3.790264e-10, 3.781402e-10, 3.774513e-10, 
    3.825717e-10, 3.800354e-10, 3.85206e-10, 3.835885e-10, 3.876515e-10, 
    3.849543e-10, 3.881954e-10, 3.875737e-10, 3.894448e-10, 3.889087e-10, 
    3.91302e-10, 3.896921e-10, 3.925426e-10, 3.909175e-10, 3.911718e-10, 
    3.89639e-10, 3.805458e-10, 3.82256e-10, 3.804445e-10, 3.806884e-10, 
    3.805789e-10, 3.792491e-10, 3.785789e-10, 3.771753e-10, 3.774301e-10, 
    3.78461e-10, 3.80798e-10, 3.800047e-10, 3.82004e-10, 3.819588e-10, 
    3.841846e-10, 3.83181e-10, 3.869219e-10, 3.858587e-10, 3.889311e-10, 
    3.881584e-10, 3.888948e-10, 3.886715e-10, 3.888977e-10, 3.877645e-10, 
    3.8825e-10, 3.872529e-10, 3.83369e-10, 3.845105e-10, 3.81106e-10, 
    3.79059e-10, 3.776992e-10, 3.767343e-10, 3.768707e-10, 3.771307e-10, 
    3.784671e-10, 3.797234e-10, 3.806808e-10, 3.813213e-10, 3.819523e-10, 
    3.838625e-10, 3.848734e-10, 3.87137e-10, 3.867284e-10, 3.874205e-10, 
    3.880816e-10, 3.891915e-10, 3.890088e-10, 3.894979e-10, 3.874022e-10, 
    3.88795e-10, 3.864957e-10, 3.871246e-10, 3.821241e-10, 3.802187e-10, 
    3.79409e-10, 3.787001e-10, 3.769756e-10, 3.781665e-10, 3.77697e-10, 
    3.788139e-10, 3.795236e-10, 3.791726e-10, 3.813388e-10, 3.804967e-10, 
    3.849333e-10, 3.830223e-10, 3.880045e-10, 3.868123e-10, 3.882902e-10, 
    3.87536e-10, 3.888283e-10, 3.876653e-10, 3.896798e-10, 3.901185e-10, 
    3.898187e-10, 3.909702e-10, 3.876008e-10, 3.888948e-10, 3.791628e-10, 
    3.7922e-10, 3.794867e-10, 3.783144e-10, 3.782427e-10, 3.771683e-10, 
    3.781243e-10, 3.785313e-10, 3.795647e-10, 3.801759e-10, 3.80757e-10, 
    3.820345e-10, 3.834613e-10, 3.854563e-10, 3.868895e-10, 3.878503e-10, 
    3.872612e-10, 3.877813e-10, 3.871999e-10, 3.869274e-10, 3.899542e-10, 
    3.882546e-10, 3.908046e-10, 3.906635e-10, 3.895095e-10, 3.906794e-10, 
    3.792602e-10, 3.789307e-10, 3.77787e-10, 3.786821e-10, 3.770513e-10, 
    3.779642e-10, 3.784891e-10, 3.805143e-10, 3.809592e-10, 3.813718e-10, 
    3.821867e-10, 3.832324e-10, 3.850669e-10, 3.86663e-10, 3.8812e-10, 
    3.880133e-10, 3.880508e-10, 3.883764e-10, 3.875701e-10, 3.885087e-10, 
    3.886663e-10, 3.882543e-10, 3.906446e-10, 3.899617e-10, 3.906605e-10, 
    3.902159e-10, 3.790378e-10, 3.795921e-10, 3.792926e-10, 3.798559e-10, 
    3.794591e-10, 3.812235e-10, 3.817525e-10, 3.842277e-10, 3.832119e-10, 
    3.848286e-10, 3.833761e-10, 3.836334e-10, 3.848814e-10, 3.834545e-10, 
    3.86575e-10, 3.844595e-10, 3.88389e-10, 3.862765e-10, 3.885214e-10, 
    3.881137e-10, 3.887887e-10, 3.893932e-10, 3.901536e-10, 3.915569e-10, 
    3.912319e-10, 3.924054e-10, 3.804185e-10, 3.811375e-10, 3.810741e-10, 
    3.818265e-10, 3.823829e-10, 3.835889e-10, 3.855231e-10, 3.847958e-10, 
    3.86131e-10, 3.863991e-10, 3.843705e-10, 3.856161e-10, 3.816186e-10, 
    3.822645e-10, 3.818799e-10, 3.804752e-10, 3.849634e-10, 3.826601e-10, 
    3.869133e-10, 3.856655e-10, 3.89307e-10, 3.874961e-10, 3.910531e-10, 
    3.925737e-10, 3.940047e-10, 3.956772e-10, 3.815298e-10, 3.810413e-10, 
    3.819159e-10, 3.831262e-10, 3.842489e-10, 3.857416e-10, 3.858943e-10, 
    3.86174e-10, 3.868983e-10, 3.875073e-10, 3.862624e-10, 3.8766e-10, 
    3.824144e-10, 3.851633e-10, 3.808566e-10, 3.821535e-10, 3.830548e-10, 
    3.826594e-10, 3.847126e-10, 3.851965e-10, 3.87163e-10, 3.861465e-10, 
    3.921984e-10, 3.895209e-10, 3.969504e-10, 3.948743e-10, 3.808706e-10, 
    3.815281e-10, 3.838164e-10, 3.827277e-10, 3.858412e-10, 3.866076e-10, 
    3.872307e-10, 3.880271e-10, 3.88113e-10, 3.885849e-10, 3.878117e-10, 
    3.885544e-10, 3.857448e-10, 3.870003e-10, 3.835548e-10, 3.843935e-10, 
    3.840077e-10, 3.835845e-10, 3.848905e-10, 3.86282e-10, 3.863117e-10, 
    3.867579e-10, 3.880153e-10, 3.858539e-10, 3.925441e-10, 3.884125e-10, 
    3.822451e-10, 3.835116e-10, 3.836924e-10, 3.832018e-10, 3.865308e-10, 
    3.853246e-10, 3.885734e-10, 3.876954e-10, 3.89134e-10, 3.884191e-10, 
    3.88314e-10, 3.873958e-10, 3.868242e-10, 3.853799e-10, 3.842048e-10, 
    3.832729e-10, 3.834896e-10, 3.845133e-10, 3.863671e-10, 3.881209e-10, 
    3.877367e-10, 3.890247e-10, 3.856155e-10, 3.870451e-10, 3.864925e-10, 
    3.879332e-10, 3.847765e-10, 3.874648e-10, 3.840893e-10, 3.843852e-10, 
    3.853007e-10, 3.871421e-10, 3.875494e-10, 3.879844e-10, 3.877159e-10, 
    3.864142e-10, 3.862009e-10, 3.852784e-10, 3.850237e-10, 3.843208e-10, 
    3.837389e-10, 3.842706e-10, 3.84829e-10, 3.864147e-10, 3.878438e-10, 
    3.894018e-10, 3.89783e-10, 3.916036e-10, 3.901217e-10, 3.925671e-10, 
    3.904881e-10, 3.940869e-10, 3.876205e-10, 3.904269e-10, 3.853423e-10, 
    3.858901e-10, 3.868809e-10, 3.891533e-10, 3.879264e-10, 3.893612e-10, 
    3.861926e-10, 3.845486e-10, 3.841232e-10, 3.833296e-10, 3.841413e-10, 
    3.840753e-10, 3.848521e-10, 3.846025e-10, 3.864674e-10, 3.854656e-10, 
    3.883114e-10, 3.893498e-10, 3.922824e-10, 3.940802e-10, 3.959101e-10, 
    3.96718e-10, 3.969639e-10, 3.970667e-10 ;

 SOIL1C_vr =
  19.97937, 19.97932, 19.97933, 19.97929, 19.97931, 19.97928, 19.97936, 
    19.97932, 19.97935, 19.97937, 19.9792, 19.97929, 19.97912, 19.97917, 
    19.97904, 19.97913, 19.97902, 19.97904, 19.97898, 19.979, 19.97892, 
    19.97897, 19.97888, 19.97894, 19.97893, 19.97898, 19.97927, 19.97921, 
    19.97927, 19.97927, 19.97927, 19.97931, 19.97933, 19.97938, 19.97937, 
    19.97934, 19.97926, 19.97929, 19.97922, 19.97922, 19.97915, 19.97918, 
    19.97906, 19.9791, 19.979, 19.97902, 19.979, 19.97901, 19.979, 19.97904, 
    19.97902, 19.97905, 19.97918, 19.97914, 19.97925, 19.97932, 19.97936, 
    19.97939, 19.97939, 19.97938, 19.97934, 19.9793, 19.97927, 19.97924, 
    19.97922, 19.97916, 19.97913, 19.97906, 19.97907, 19.97905, 19.97902, 
    19.97899, 19.979, 19.97898, 19.97905, 19.979, 19.97908, 19.97906, 
    19.97922, 19.97928, 19.97931, 19.97933, 19.97939, 19.97935, 19.97936, 
    19.97932, 19.9793, 19.97931, 19.97924, 19.97927, 19.97913, 19.97919, 
    19.97903, 19.97907, 19.97902, 19.97904, 19.979, 19.97904, 19.97897, 
    19.97896, 19.97897, 19.97893, 19.97904, 19.979, 19.97931, 19.97931, 
    19.9793, 19.97934, 19.97934, 19.97938, 19.97935, 19.97933, 19.9793, 
    19.97928, 19.97926, 19.97922, 19.97917, 19.97911, 19.97906, 19.97903, 
    19.97905, 19.97903, 19.97905, 19.97906, 19.97897, 19.97902, 19.97894, 
    19.97894, 19.97898, 19.97894, 19.97931, 19.97932, 19.97936, 19.97933, 
    19.97938, 19.97935, 19.97934, 19.97927, 19.97926, 19.97924, 19.97922, 
    19.97918, 19.97912, 19.97907, 19.97902, 19.97903, 19.97903, 19.97902, 
    19.97904, 19.97901, 19.97901, 19.97902, 19.97894, 19.97897, 19.97894, 
    19.97896, 19.97932, 19.9793, 19.97931, 19.97929, 19.9793, 19.97925, 
    19.97923, 19.97915, 19.97918, 19.97913, 19.97918, 19.97917, 19.97913, 
    19.97918, 19.97907, 19.97914, 19.97902, 19.97908, 19.97901, 19.97902, 
    19.979, 19.97898, 19.97896, 19.97891, 19.97892, 19.97889, 19.97927, 
    19.97925, 19.97925, 19.97923, 19.97921, 19.97917, 19.97911, 19.97913, 
    19.97909, 19.97908, 19.97915, 19.9791, 19.97923, 19.97921, 19.97923, 
    19.97927, 19.97913, 19.9792, 19.97906, 19.9791, 19.97899, 19.97904, 
    19.97893, 19.97888, 19.97884, 19.97878, 19.97924, 19.97925, 19.97923, 
    19.97919, 19.97915, 19.9791, 19.9791, 19.97909, 19.97906, 19.97904, 
    19.97908, 19.97904, 19.97921, 19.97912, 19.97926, 19.97922, 19.97919, 
    19.9792, 19.97913, 19.97912, 19.97906, 19.97909, 19.97889, 19.97898, 
    19.97874, 19.97881, 19.97926, 19.97924, 19.97916, 19.9792, 19.9791, 
    19.97907, 19.97905, 19.97903, 19.97902, 19.97901, 19.97903, 19.97901, 
    19.9791, 19.97906, 19.97917, 19.97915, 19.97916, 19.97917, 19.97913, 
    19.97908, 19.97908, 19.97907, 19.97903, 19.9791, 19.97888, 19.97902, 
    19.97921, 19.97917, 19.97917, 19.97918, 19.97908, 19.97911, 19.97901, 
    19.97904, 19.97899, 19.97902, 19.97902, 19.97905, 19.97907, 19.97911, 
    19.97915, 19.97918, 19.97917, 19.97914, 19.97908, 19.97902, 19.97904, 
    19.97899, 19.9791, 19.97906, 19.97908, 19.97903, 19.97913, 19.97905, 
    19.97915, 19.97915, 19.97911, 19.97906, 19.97904, 19.97903, 19.97904, 
    19.97908, 19.97909, 19.97912, 19.97912, 19.97915, 19.97917, 19.97915, 
    19.97913, 19.97908, 19.97903, 19.97898, 19.97897, 19.97891, 19.97896, 
    19.97888, 19.97895, 19.97883, 19.97904, 19.97895, 19.97911, 19.9791, 
    19.97906, 19.97899, 19.97903, 19.97898, 19.97909, 19.97914, 19.97915, 
    19.97918, 19.97915, 19.97915, 19.97913, 19.97914, 19.97908, 19.97911, 
    19.97902, 19.97898, 19.97889, 19.97883, 19.97878, 19.97875, 19.97874, 
    19.97874,
  19.981, 19.98093, 19.98094, 19.98088, 19.98091, 19.98088, 19.98098, 
    19.98092, 19.98096, 19.98099, 19.98077, 19.98088, 19.98066, 19.98073, 
    19.98055, 19.98067, 19.98053, 19.98056, 19.98048, 19.9805, 19.9804, 
    19.98047, 19.98035, 19.98042, 19.9804, 19.98047, 19.98086, 19.98079, 
    19.98086, 19.98085, 19.98086, 19.98091, 19.98094, 19.981, 19.98099, 
    19.98095, 19.98085, 19.98088, 19.98079, 19.9808, 19.9807, 19.98075, 
    19.98059, 19.98063, 19.9805, 19.98053, 19.9805, 19.98051, 19.9805, 
    19.98055, 19.98053, 19.98057, 19.98074, 19.98069, 19.98083, 19.98092, 
    19.98098, 19.98102, 19.98101, 19.981, 19.98095, 19.98089, 19.98085, 
    19.98083, 19.9808, 19.98072, 19.98067, 19.98058, 19.98059, 19.98056, 
    19.98054, 19.98049, 19.9805, 19.98048, 19.98056, 19.9805, 19.9806, 
    19.98058, 19.98079, 19.98087, 19.98091, 19.98094, 19.98101, 19.98096, 
    19.98098, 19.98093, 19.9809, 19.98092, 19.98082, 19.98086, 19.98067, 
    19.98075, 19.98054, 19.98059, 19.98053, 19.98056, 19.9805, 19.98055, 
    19.98047, 19.98045, 19.98046, 19.98041, 19.98056, 19.9805, 19.98092, 
    19.98092, 19.9809, 19.98095, 19.98096, 19.981, 19.98096, 19.98094, 
    19.9809, 19.98087, 19.98085, 19.98079, 19.98073, 19.98065, 19.98059, 
    19.98055, 19.98057, 19.98055, 19.98057, 19.98059, 19.98046, 19.98053, 
    19.98042, 19.98043, 19.98047, 19.98042, 19.98091, 19.98093, 19.98098, 
    19.98094, 19.98101, 19.98097, 19.98095, 19.98086, 19.98084, 19.98082, 
    19.98079, 19.98074, 19.98067, 19.9806, 19.98053, 19.98054, 19.98054, 
    19.98052, 19.98056, 19.98052, 19.98051, 19.98053, 19.98043, 19.98046, 
    19.98043, 19.98045, 19.98092, 19.9809, 19.98091, 19.98089, 19.9809, 
    19.98083, 19.98081, 19.9807, 19.98074, 19.98067, 19.98074, 19.98073, 
    19.98067, 19.98073, 19.9806, 19.98069, 19.98052, 19.98061, 19.98052, 
    19.98054, 19.98051, 19.98048, 19.98045, 19.98039, 19.9804, 19.98035, 
    19.98086, 19.98083, 19.98083, 19.9808, 19.98078, 19.98073, 19.98064, 
    19.98068, 19.98062, 19.98061, 19.98069, 19.98064, 19.98081, 19.98078, 
    19.9808, 19.98086, 19.98067, 19.98077, 19.98059, 19.98064, 19.98048, 
    19.98056, 19.98041, 19.98034, 19.98028, 19.98021, 19.98082, 19.98084, 
    19.9808, 19.98075, 19.9807, 19.98064, 19.98063, 19.98062, 19.98059, 
    19.98056, 19.98061, 19.98055, 19.98078, 19.98066, 19.98084, 19.98079, 
    19.98075, 19.98077, 19.98068, 19.98066, 19.98058, 19.98062, 19.98036, 
    19.98047, 19.98016, 19.98025, 19.98084, 19.98082, 19.98072, 19.98076, 
    19.98063, 19.9806, 19.98057, 19.98054, 19.98054, 19.98051, 19.98055, 
    19.98052, 19.98064, 19.98058, 19.98073, 19.98069, 19.98071, 19.98073, 
    19.98067, 19.98061, 19.98061, 19.98059, 19.98054, 19.98063, 19.98035, 
    19.98052, 19.98079, 19.98073, 19.98072, 19.98074, 19.9806, 19.98065, 
    19.98051, 19.98055, 19.98049, 19.98052, 19.98053, 19.98057, 19.98059, 
    19.98065, 19.9807, 19.98074, 19.98073, 19.98069, 19.98061, 19.98053, 
    19.98055, 19.9805, 19.98064, 19.98058, 19.9806, 19.98054, 19.98068, 
    19.98056, 19.98071, 19.98069, 19.98065, 19.98058, 19.98056, 19.98054, 
    19.98055, 19.98061, 19.98062, 19.98066, 19.98067, 19.9807, 19.98072, 
    19.9807, 19.98067, 19.98061, 19.98055, 19.98048, 19.98046, 19.98039, 
    19.98045, 19.98034, 19.98043, 19.98028, 19.98056, 19.98044, 19.98065, 
    19.98063, 19.98059, 19.98049, 19.98054, 19.98048, 19.98062, 19.98069, 
    19.98071, 19.98074, 19.9807, 19.98071, 19.98067, 19.98068, 19.9806, 
    19.98065, 19.98053, 19.98048, 19.98036, 19.98028, 19.9802, 19.98017, 
    19.98016, 19.98015,
  19.98272, 19.98265, 19.98266, 19.9826, 19.98263, 19.98259, 19.98271, 
    19.98264, 19.98268, 19.98272, 19.98248, 19.9826, 19.98236, 19.98244, 
    19.98225, 19.98237, 19.98223, 19.98225, 19.98217, 19.98219, 19.98208, 
    19.98216, 19.98203, 19.9821, 19.98209, 19.98216, 19.98257, 19.9825, 
    19.98258, 19.98257, 19.98257, 19.98263, 19.98266, 19.98273, 19.98272, 
    19.98267, 19.98256, 19.9826, 19.98251, 19.98251, 19.98241, 19.98245, 
    19.98228, 19.98233, 19.98219, 19.98223, 19.98219, 19.9822, 19.98219, 
    19.98224, 19.98222, 19.98227, 19.98244, 19.98239, 19.98255, 19.98264, 
    19.9827, 19.98275, 19.98274, 19.98273, 19.98267, 19.98261, 19.98257, 
    19.98254, 19.98251, 19.98242, 19.98238, 19.98227, 19.98229, 19.98226, 
    19.98223, 19.98218, 19.98219, 19.98217, 19.98226, 19.9822, 19.9823, 
    19.98227, 19.9825, 19.98259, 19.98263, 19.98266, 19.98274, 19.98268, 
    19.9827, 19.98265, 19.98262, 19.98264, 19.98254, 19.98258, 19.98237, 
    19.98246, 19.98223, 19.98229, 19.98222, 19.98226, 19.9822, 19.98225, 
    19.98216, 19.98214, 19.98215, 19.9821, 19.98225, 19.98219, 19.98264, 
    19.98263, 19.98262, 19.98268, 19.98268, 19.98273, 19.98269, 19.98267, 
    19.98262, 19.98259, 19.98256, 19.98251, 19.98244, 19.98235, 19.98228, 
    19.98224, 19.98227, 19.98224, 19.98227, 19.98228, 19.98215, 19.98222, 
    19.98211, 19.98211, 19.98217, 19.98211, 19.98263, 19.98265, 19.9827, 
    19.98266, 19.98273, 19.98269, 19.98267, 19.98257, 19.98256, 19.98254, 
    19.9825, 19.98245, 19.98237, 19.9823, 19.98223, 19.98223, 19.98223, 
    19.98222, 19.98225, 19.98221, 19.9822, 19.98222, 19.98211, 19.98215, 
    19.98211, 19.98213, 19.98264, 19.98262, 19.98263, 19.9826, 19.98262, 
    19.98254, 19.98252, 19.98241, 19.98245, 19.98238, 19.98244, 19.98243, 
    19.98238, 19.98244, 19.9823, 19.9824, 19.98222, 19.98231, 19.98221, 
    19.98223, 19.9822, 19.98217, 19.98214, 19.98207, 19.98209, 19.98203, 
    19.98258, 19.98255, 19.98255, 19.98252, 19.98249, 19.98244, 19.98235, 
    19.98238, 19.98232, 19.98231, 19.9824, 19.98234, 19.98252, 19.9825, 
    19.98251, 19.98258, 19.98237, 19.98248, 19.98228, 19.98234, 19.98217, 
    19.98226, 19.9821, 19.98203, 19.98196, 19.98189, 19.98253, 19.98255, 
    19.98251, 19.98246, 19.9824, 19.98234, 19.98233, 19.98232, 19.98228, 
    19.98226, 19.98231, 19.98225, 19.98249, 19.98236, 19.98256, 19.9825, 
    19.98246, 19.98248, 19.98238, 19.98236, 19.98227, 19.98232, 19.98204, 
    19.98216, 19.98183, 19.98192, 19.98256, 19.98253, 19.98243, 19.98248, 
    19.98233, 19.9823, 19.98227, 19.98223, 19.98223, 19.98221, 19.98224, 
    19.98221, 19.98234, 19.98228, 19.98244, 19.9824, 19.98242, 19.98244, 
    19.98238, 19.98231, 19.98231, 19.98229, 19.98223, 19.98233, 19.98203, 
    19.98222, 19.9825, 19.98244, 19.98243, 19.98245, 19.9823, 19.98236, 
    19.98221, 19.98225, 19.98218, 19.98222, 19.98222, 19.98226, 19.98229, 
    19.98235, 19.98241, 19.98245, 19.98244, 19.98239, 19.98231, 19.98223, 
    19.98225, 19.98219, 19.98234, 19.98228, 19.9823, 19.98224, 19.98238, 
    19.98226, 19.98241, 19.9824, 19.98236, 19.98227, 19.98225, 19.98223, 
    19.98225, 19.98231, 19.98232, 19.98236, 19.98237, 19.9824, 19.98243, 
    19.9824, 19.98238, 19.98231, 19.98224, 19.98217, 19.98215, 19.98207, 
    19.98214, 19.98203, 19.98212, 19.98196, 19.98225, 19.98212, 19.98236, 
    19.98233, 19.98228, 19.98218, 19.98224, 19.98217, 19.98232, 19.98239, 
    19.98241, 19.98245, 19.98241, 19.98241, 19.98238, 19.98239, 19.9823, 
    19.98235, 19.98222, 19.98217, 19.98204, 19.98196, 19.98187, 19.98184, 
    19.98183, 19.98182,
  19.9841, 19.98402, 19.98404, 19.98398, 19.98401, 19.98397, 19.98408, 
    19.98402, 19.98406, 19.98409, 19.98386, 19.98397, 19.98374, 19.98381, 
    19.98363, 19.98375, 19.98361, 19.98363, 19.98355, 19.98357, 19.98347, 
    19.98354, 19.98341, 19.98348, 19.98347, 19.98354, 19.98395, 19.98388, 
    19.98396, 19.98395, 19.98395, 19.98401, 19.98404, 19.9841, 19.98409, 
    19.98405, 19.98394, 19.98398, 19.98389, 19.98389, 19.98379, 19.98383, 
    19.98366, 19.98371, 19.98357, 19.98361, 19.98357, 19.98359, 19.98357, 
    19.98363, 19.9836, 19.98365, 19.98382, 19.98377, 19.98393, 19.98402, 
    19.98408, 19.98413, 19.98412, 19.98411, 19.98405, 19.98399, 19.98395, 
    19.98392, 19.98389, 19.9838, 19.98376, 19.98365, 19.98367, 19.98364, 
    19.98361, 19.98356, 19.98357, 19.98355, 19.98364, 19.98358, 19.98368, 
    19.98365, 19.98388, 19.98397, 19.984, 19.98404, 19.98411, 19.98406, 
    19.98408, 19.98403, 19.984, 19.98401, 19.98392, 19.98396, 19.98375, 
    19.98384, 19.98362, 19.98367, 19.9836, 19.98364, 19.98358, 19.98363, 
    19.98354, 19.98352, 19.98353, 19.98348, 19.98363, 19.98357, 19.98401, 
    19.98401, 19.984, 19.98405, 19.98406, 19.9841, 19.98406, 19.98404, 
    19.984, 19.98397, 19.98394, 19.98388, 19.98382, 19.98373, 19.98367, 
    19.98362, 19.98365, 19.98363, 19.98365, 19.98366, 19.98353, 19.9836, 
    19.98349, 19.9835, 19.98355, 19.98349, 19.98401, 19.98403, 19.98408, 
    19.98404, 19.98411, 19.98407, 19.98405, 19.98395, 19.98393, 19.98392, 
    19.98388, 19.98383, 19.98375, 19.98368, 19.98361, 19.98361, 19.98361, 
    19.9836, 19.98363, 19.98359, 19.98359, 19.9836, 19.9835, 19.98353, 
    19.9835, 19.98351, 19.98402, 19.984, 19.98401, 19.98398, 19.984, 
    19.98392, 19.9839, 19.98379, 19.98383, 19.98376, 19.98382, 19.98381, 
    19.98376, 19.98382, 19.98368, 19.98378, 19.9836, 19.98369, 19.98359, 
    19.98361, 19.98358, 19.98355, 19.98352, 19.98345, 19.98347, 19.98342, 
    19.98396, 19.98392, 19.98393, 19.98389, 19.98387, 19.98381, 19.98373, 
    19.98376, 19.9837, 19.98369, 19.98378, 19.98372, 19.9839, 19.98388, 
    19.98389, 19.98396, 19.98375, 19.98386, 19.98366, 19.98372, 19.98356, 
    19.98364, 19.98348, 19.98341, 19.98334, 19.98327, 19.98391, 19.98393, 
    19.98389, 19.98384, 19.98379, 19.98372, 19.98371, 19.9837, 19.98367, 
    19.98364, 19.98369, 19.98363, 19.98387, 19.98374, 19.98394, 19.98388, 
    19.98384, 19.98386, 19.98376, 19.98374, 19.98365, 19.9837, 19.98343, 
    19.98355, 19.98321, 19.9833, 19.98394, 19.98391, 19.9838, 19.98385, 
    19.98371, 19.98368, 19.98365, 19.98361, 19.98361, 19.98359, 19.98362, 
    19.98359, 19.98372, 19.98366, 19.98382, 19.98378, 19.9838, 19.98381, 
    19.98376, 19.98369, 19.98369, 19.98367, 19.98361, 19.98371, 19.98341, 
    19.9836, 19.98388, 19.98382, 19.98381, 19.98383, 19.98368, 19.98374, 
    19.98359, 19.98363, 19.98356, 19.9836, 19.9836, 19.98364, 19.98367, 
    19.98373, 19.98379, 19.98383, 19.98382, 19.98377, 19.98369, 19.98361, 
    19.98363, 19.98357, 19.98372, 19.98366, 19.98368, 19.98362, 19.98376, 
    19.98364, 19.98379, 19.98378, 19.98374, 19.98365, 19.98363, 19.98362, 
    19.98363, 19.98369, 19.9837, 19.98374, 19.98375, 19.98378, 19.98381, 
    19.98378, 19.98376, 19.98369, 19.98362, 19.98355, 19.98353, 19.98345, 
    19.98352, 19.98341, 19.9835, 19.98334, 19.98363, 19.98351, 19.98374, 
    19.98371, 19.98367, 19.98356, 19.98362, 19.98355, 19.9837, 19.98377, 
    19.98379, 19.98383, 19.98379, 19.98379, 19.98376, 19.98377, 19.98368, 
    19.98373, 19.9836, 19.98355, 19.98342, 19.98334, 19.98326, 19.98322, 
    19.98321, 19.98321,
  19.9857, 19.98564, 19.98565, 19.9856, 19.98563, 19.98559, 19.98569, 
    19.98564, 19.98567, 19.9857, 19.98549, 19.9856, 19.98539, 19.98545, 
    19.98529, 19.9854, 19.98527, 19.98529, 19.98522, 19.98524, 19.98514, 
    19.98521, 19.98509, 19.98516, 19.98515, 19.98521, 19.98557, 19.98551, 
    19.98558, 19.98557, 19.98557, 19.98563, 19.98565, 19.98571, 19.9857, 
    19.98566, 19.98557, 19.9856, 19.98552, 19.98552, 19.98543, 19.98547, 
    19.98532, 19.98536, 19.98524, 19.98527, 19.98524, 19.98525, 19.98524, 
    19.98528, 19.98527, 19.98531, 19.98546, 19.98542, 19.98555, 19.98563, 
    19.98569, 19.98573, 19.98572, 19.98571, 19.98566, 19.98561, 19.98557, 
    19.98554, 19.98552, 19.98544, 19.9854, 19.98531, 19.98533, 19.9853, 
    19.98527, 19.98523, 19.98524, 19.98521, 19.9853, 19.98524, 19.98534, 
    19.98531, 19.98551, 19.98559, 19.98562, 19.98565, 19.98572, 19.98567, 
    19.98569, 19.98564, 19.98561, 19.98563, 19.98554, 19.98558, 19.9854, 
    19.98548, 19.98528, 19.98532, 19.98526, 19.98529, 19.98524, 19.98529, 
    19.98521, 19.98519, 19.9852, 19.98516, 19.98529, 19.98524, 19.98563, 
    19.98563, 19.98562, 19.98566, 19.98567, 19.98571, 19.98567, 19.98565, 
    19.98561, 19.98559, 19.98557, 19.98552, 19.98546, 19.98538, 19.98532, 
    19.98528, 19.98531, 19.98528, 19.98531, 19.98532, 19.9852, 19.98527, 
    19.98516, 19.98517, 19.98521, 19.98517, 19.98563, 19.98564, 19.98569, 
    19.98565, 19.98571, 19.98568, 19.98566, 19.98558, 19.98556, 19.98554, 
    19.98551, 19.98547, 19.98539, 19.98533, 19.98527, 19.98528, 19.98527, 
    19.98526, 19.98529, 19.98525, 19.98525, 19.98527, 19.98517, 19.9852, 
    19.98517, 19.98519, 19.98564, 19.98561, 19.98562, 19.9856, 19.98562, 
    19.98555, 19.98553, 19.98543, 19.98547, 19.9854, 19.98546, 19.98545, 
    19.9854, 19.98546, 19.98533, 19.98542, 19.98526, 19.98534, 19.98525, 
    19.98527, 19.98524, 19.98522, 19.98519, 19.98513, 19.98515, 19.9851, 
    19.98558, 19.98555, 19.98555, 19.98552, 19.9855, 19.98545, 19.98537, 
    19.9854, 19.98535, 19.98534, 19.98542, 19.98537, 19.98553, 19.98551, 
    19.98552, 19.98558, 19.9854, 19.98549, 19.98532, 19.98537, 19.98522, 
    19.9853, 19.98515, 19.98509, 19.98503, 19.98497, 19.98553, 19.98556, 
    19.98552, 19.98547, 19.98543, 19.98537, 19.98536, 19.98535, 19.98532, 
    19.98529, 19.98535, 19.98529, 19.9855, 19.98539, 19.98556, 19.98551, 
    19.98547, 19.98549, 19.98541, 19.98539, 19.98531, 19.98535, 19.98511, 
    19.98521, 19.98491, 19.985, 19.98556, 19.98553, 19.98544, 19.98549, 
    19.98536, 19.98533, 19.98531, 19.98527, 19.98527, 19.98525, 19.98528, 
    19.98525, 19.98537, 19.98532, 19.98545, 19.98542, 19.98544, 19.98545, 
    19.9854, 19.98534, 19.98534, 19.98532, 19.98528, 19.98536, 19.98509, 
    19.98526, 19.98551, 19.98546, 19.98545, 19.98547, 19.98533, 19.98538, 
    19.98525, 19.98529, 19.98523, 19.98526, 19.98526, 19.9853, 19.98532, 
    19.98538, 19.98543, 19.98547, 19.98546, 19.98541, 19.98534, 19.98527, 
    19.98529, 19.98523, 19.98537, 19.98531, 19.98534, 19.98528, 19.9854, 
    19.9853, 19.98543, 19.98542, 19.98538, 19.98531, 19.98529, 19.98528, 
    19.98529, 19.98534, 19.98535, 19.98538, 19.9854, 19.98542, 19.98545, 
    19.98543, 19.9854, 19.98534, 19.98528, 19.98522, 19.9852, 19.98513, 
    19.98519, 19.98509, 19.98517, 19.98503, 19.98529, 19.98518, 19.98538, 
    19.98536, 19.98532, 19.98523, 19.98528, 19.98522, 19.98535, 19.98541, 
    19.98543, 19.98546, 19.98543, 19.98543, 19.9854, 19.98541, 19.98534, 
    19.98538, 19.98526, 19.98522, 19.9851, 19.98503, 19.98496, 19.98492, 
    19.98491, 19.98491,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222453, 0.7222427, 0.7222432, 0.7222412, 0.7222423, 0.722241, 0.7222447, 
    0.7222427, 0.722244, 0.722245, 0.7222372, 0.7222411, 0.7222332, 
    0.7222357, 0.7222295, 0.7222336, 0.7222287, 0.7222296, 0.7222268, 
    0.7222276, 0.7222239, 0.7222264, 0.7222221, 0.7222245, 0.7222242, 
    0.7222265, 0.7222403, 0.7222377, 0.7222404, 0.7222401, 0.7222403, 
    0.7222423, 0.7222433, 0.7222455, 0.722245, 0.7222435, 0.7222399, 
    0.7222412, 0.7222381, 0.7222382, 0.7222348, 0.7222363, 0.7222306, 
    0.7222322, 0.7222276, 0.7222288, 0.7222276, 0.7222279, 0.7222276, 
    0.7222294, 0.7222286, 0.7222301, 0.722236, 0.7222343, 0.7222395, 
    0.7222426, 0.7222446, 0.7222461, 0.7222459, 0.7222455, 0.7222435, 
    0.7222416, 0.7222401, 0.7222391, 0.7222382, 0.7222353, 0.7222337, 
    0.7222303, 0.7222309, 0.7222298, 0.7222289, 0.7222272, 0.7222275, 
    0.7222267, 0.7222299, 0.7222278, 0.7222313, 0.7222303, 0.7222379, 
    0.7222408, 0.7222421, 0.7222431, 0.7222458, 0.722244, 0.7222447, 
    0.722243, 0.7222419, 0.7222424, 0.7222391, 0.7222404, 0.7222337, 
    0.7222366, 0.7222289, 0.7222308, 0.7222285, 0.7222297, 0.7222277, 
    0.7222295, 0.7222264, 0.7222258, 0.7222262, 0.7222245, 0.7222296, 
    0.7222276, 0.7222424, 0.7222424, 0.7222419, 0.7222437, 0.7222438, 
    0.7222455, 0.722244, 0.7222434, 0.7222418, 0.7222409, 0.72224, 0.7222381, 
    0.7222359, 0.7222328, 0.7222307, 0.7222292, 0.7222301, 0.7222293, 
    0.7222302, 0.7222306, 0.722226, 0.7222286, 0.7222247, 0.722225, 
    0.7222267, 0.7222249, 0.7222423, 0.7222428, 0.7222445, 0.7222431, 
    0.7222456, 0.7222443, 0.7222434, 0.7222404, 0.7222397, 0.7222391, 
    0.7222378, 0.7222362, 0.7222334, 0.722231, 0.7222288, 0.7222289, 
    0.7222289, 0.7222284, 0.7222297, 0.7222282, 0.722228, 0.7222286, 
    0.722225, 0.722226, 0.722225, 0.7222256, 0.7222426, 0.7222418, 0.7222422, 
    0.7222413, 0.722242, 0.7222393, 0.7222385, 0.7222347, 0.7222363, 
    0.7222338, 0.722236, 0.7222356, 0.7222337, 0.7222359, 0.7222311, 
    0.7222344, 0.7222284, 0.7222316, 0.7222282, 0.7222288, 0.7222278, 
    0.7222269, 0.7222257, 0.7222236, 0.7222241, 0.7222223, 0.7222405, 
    0.7222394, 0.7222395, 0.7222384, 0.7222375, 0.7222357, 0.7222328, 
    0.7222338, 0.7222318, 0.7222314, 0.7222345, 0.7222326, 0.7222387, 
    0.7222377, 0.7222383, 0.7222404, 0.7222336, 0.7222371, 0.7222306, 
    0.7222325, 0.722227, 0.7222297, 0.7222244, 0.722222, 0.7222198, 
    0.7222173, 0.7222388, 0.7222396, 0.7222382, 0.7222364, 0.7222347, 
    0.7222324, 0.7222322, 0.7222317, 0.7222307, 0.7222297, 0.7222316, 
    0.7222295, 0.7222375, 0.7222333, 0.7222399, 0.7222379, 0.7222365, 
    0.7222371, 0.722234, 0.7222332, 0.7222303, 0.7222318, 0.7222226, 
    0.7222267, 0.7222154, 0.7222185, 0.7222399, 0.7222388, 0.7222353, 
    0.722237, 0.7222323, 0.7222311, 0.7222301, 0.7222289, 0.7222288, 
    0.7222281, 0.7222292, 0.7222281, 0.7222324, 0.7222305, 0.7222357, 
    0.7222345, 0.722235, 0.7222357, 0.7222337, 0.7222316, 0.7222316, 
    0.7222309, 0.7222289, 0.7222322, 0.7222221, 0.7222283, 0.7222377, 
    0.7222358, 0.7222356, 0.7222363, 0.7222312, 0.7222331, 0.7222281, 
    0.7222294, 0.7222273, 0.7222283, 0.7222285, 0.7222299, 0.7222308, 
    0.7222329, 0.7222347, 0.7222362, 0.7222359, 0.7222343, 0.7222314, 
    0.7222288, 0.7222294, 0.7222274, 0.7222326, 0.7222304, 0.7222313, 
    0.7222291, 0.7222339, 0.7222298, 0.7222349, 0.7222345, 0.7222331, 
    0.7222303, 0.7222297, 0.722229, 0.7222294, 0.7222314, 0.7222317, 
    0.7222331, 0.7222335, 0.7222345, 0.7222354, 0.7222347, 0.7222338, 
    0.7222314, 0.7222292, 0.7222269, 0.7222263, 0.7222235, 0.7222257, 
    0.722222, 0.7222252, 0.7222197, 0.7222295, 0.7222253, 0.722233, 
    0.7222322, 0.7222307, 0.7222272, 0.7222291, 0.7222269, 0.7222317, 
    0.7222342, 0.7222349, 0.7222361, 0.7222348, 0.722235, 0.7222338, 
    0.7222341, 0.7222313, 0.7222328, 0.7222285, 0.7222269, 0.7222224, 
    0.7222197, 0.722217, 0.7222157, 0.7222154, 0.7222152 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  -5.139921e-21, -4.111937e-20, 1.541976e-20, -2.055969e-20, -5.139921e-20, 
    2.055969e-20, 1.541976e-20, 1.541976e-20, 1.027984e-20, -2.569961e-20, 
    3.597945e-20, -2.055969e-20, 2.569961e-20, 1.541976e-20, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -2.569961e-20, 0, -2.055969e-20, 
    3.083953e-20, -1.541976e-20, -2.055969e-20, -5.139921e-21, 1.027984e-20, 
    3.083953e-20, 1.541976e-20, 1.027984e-20, -4.111937e-20, 5.139921e-21, 
    5.139921e-21, 2.055969e-20, 0, -5.139921e-21, -1.541976e-20, 0, 
    1.541976e-20, 2.055969e-20, -5.139921e-21, 2.569961e-20, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, -3.597945e-20, 2.055969e-20, -2.006177e-36, 
    -1.027984e-20, -1.027984e-20, 2.569961e-20, 5.139921e-21, -2.055969e-20, 
    1.541976e-20, 1.541976e-20, -5.139921e-21, 2.569961e-20, 2.569961e-20, 
    2.055969e-20, 2.569961e-20, 1.541976e-20, 2.569961e-20, 1.027984e-20, 0, 
    -1.541976e-20, -1.541976e-20, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 0, -5.139921e-21, 2.055969e-20, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, -4.111937e-20, -2.055969e-20, 
    -1.027984e-20, 1.541976e-20, 2.569961e-20, 1.027984e-20, -5.139921e-21, 
    -4.625929e-20, -3.083953e-20, 2.006177e-36, 5.139921e-21, -2.055969e-20, 
    3.597945e-20, 3.597945e-20, 1.027984e-20, 1.541976e-20, 5.139921e-21, 
    -1.027984e-20, 1.541976e-20, 2.055969e-20, 5.139921e-21, -2.569961e-20, 
    1.027984e-20, 1.027984e-20, 2.569961e-20, 3.597945e-20, 3.083953e-20, 
    -5.139921e-21, 1.541976e-20, -1.027984e-20, 3.597945e-20, 4.111937e-20, 
    2.569961e-20, 1.027984e-20, -2.055969e-20, -1.541976e-20, 5.653913e-20, 
    0, 4.111937e-20, -1.541976e-20, 3.083953e-20, 5.139921e-21, 0, 
    -2.569961e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -2.569961e-20, 1.541976e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    1.541976e-20, 1.541976e-20, -1.027984e-20, -5.139921e-21, -1.541976e-20, 
    -1.541976e-20, 2.055969e-20, -1.027984e-20, -2.055969e-20, -1.027984e-20, 
    2.569961e-20, -1.541976e-20, -2.055969e-20, -2.569961e-20, 2.055969e-20, 
    -4.625929e-20, -2.055969e-20, -1.541976e-20, -2.006177e-36, 
    -5.139921e-21, -1.541976e-20, -3.083953e-20, -2.055969e-20, 5.139921e-21, 
    2.569961e-20, -2.569961e-20, -2.569961e-20, -5.139921e-21, -1.027984e-20, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, 2.055969e-20, 
    -1.541976e-20, 2.006177e-36, 2.569961e-20, 1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, 3.597945e-20, 2.055969e-20, 
    2.055969e-20, -2.055969e-20, -2.569961e-20, -1.027984e-20, -5.139921e-21, 
    0, -2.055969e-20, -1.027984e-20, 1.541976e-20, 1.027984e-20, 
    2.006177e-36, 5.139921e-21, 2.006177e-36, -2.055969e-20, -5.139921e-21, 
    -5.139921e-21, 2.055969e-20, -1.027984e-20, 5.139921e-21, -2.006177e-36, 
    1.027984e-20, -3.083953e-20, -1.027984e-20, 4.111937e-20, -1.027984e-20, 
    -1.541976e-20, 1.027984e-20, 2.569961e-20, 2.055969e-20, -2.569961e-20, 
    -1.027984e-20, -2.569961e-20, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    1.541976e-20, 1.027984e-20, 3.597945e-20, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 1.027984e-20, 1.541976e-20, -2.569961e-20, 
    1.541976e-20, 5.139921e-21, -2.055969e-20, -3.597945e-20, -5.139921e-21, 
    2.055969e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 2.569961e-20, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, -1.541976e-20, 1.541976e-20, 
    -5.139921e-21, 2.055969e-20, 1.541976e-20, -3.083953e-20, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, -2.569961e-20, -1.027984e-20, 
    1.541976e-20, 2.569961e-20, 5.139921e-21, 2.006177e-36, -5.139921e-21, 
    2.569961e-20, 1.541976e-20, 2.569961e-20, 2.055969e-20, -5.139921e-21, 
    -1.541976e-20, 3.083953e-20, 2.006177e-36, 1.027984e-20, 1.541976e-20, 
    -2.055969e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 3.597945e-20, 
    2.055969e-20, 1.027984e-20, -2.569961e-20, -2.055969e-20, 5.139921e-21, 
    2.569961e-20, 2.006177e-36, 5.139921e-21, 4.625929e-20, 1.027984e-20, 
    -2.006177e-36, -1.027984e-20, 0, 1.027984e-20, 5.139921e-21, 
    1.541976e-20, 1.027984e-20, -5.139921e-20, 0, 2.006177e-36, 5.139921e-21, 
    -2.055969e-20, 0, 1.027984e-20, 2.569961e-20, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 5.139921e-21, 1.027984e-20, -2.569961e-20, 
    2.006177e-36, 1.541976e-20, -1.027984e-20, 2.006177e-36, 5.139921e-21, 0, 
    1.541976e-20, -3.083953e-20, 1.541976e-20, 1.027984e-20, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, -2.569961e-20, 1.027984e-20, 
    -2.006177e-36, 0, 1.027984e-20, 1.027984e-20, 2.055969e-20, 
    -3.083953e-20, 5.139921e-21, -2.055969e-20, -5.139921e-21, -2.569961e-20, 
    -5.139921e-21, -2.055969e-20, -1.541976e-20, 1.541976e-20, 0, 
    -1.027984e-20, 0, -1.027984e-20, 2.569961e-20, -2.569961e-20, 
    1.027984e-20, -4.625929e-20, -5.139921e-21, -2.569961e-20, 0,
  5.139921e-21, -1.027984e-20, 1.027984e-20, 1.541976e-20, -1.541976e-20, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -3.597945e-20, -1.027984e-20, -1.541976e-20, 
    -1.541976e-20, -1.027984e-20, 3.083953e-20, 1.541976e-20, -1.541976e-20, 
    -2.006177e-36, 5.139921e-21, -2.055969e-20, 5.139921e-21, -1.027984e-20, 
    2.006177e-36, -1.027984e-20, 5.139921e-21, 5.139921e-21, 1.541976e-20, 
    3.597945e-20, 2.055969e-20, 0, 1.541976e-20, -5.139921e-21, 1.541976e-20, 
    2.006177e-36, 5.139921e-21, -2.006177e-36, 2.006177e-36, -5.139921e-21, 
    2.569961e-20, -2.006177e-36, -1.027984e-20, 2.006177e-36, 1.541976e-20, 
    -1.541976e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 2.006177e-36, 
    -2.055969e-20, -5.139921e-21, 2.055969e-20, 2.569961e-20, -3.083953e-20, 
    1.541976e-20, 2.006177e-36, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -1.541976e-20, -1.027984e-20, 2.055969e-20, 1.027984e-20, 1.027984e-20, 
    -5.139921e-21, 2.055969e-20, 2.006177e-36, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 2.055969e-20, -1.027984e-20, -5.139921e-21, -1.541976e-20, 
    3.597945e-20, 0, 1.027984e-20, 0, 1.027984e-20, 1.541976e-20, 
    -2.569961e-20, -5.139921e-21, -5.139921e-21, 0, 1.027984e-20, 
    -5.139921e-21, 0, 1.541976e-20, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 1.541976e-20, -2.006177e-36, 2.055969e-20, -2.055969e-20, 
    1.027984e-20, 0, 1.541976e-20, -3.083953e-20, 0, -5.139921e-21, 
    -5.139921e-21, -2.006177e-36, -2.055969e-20, 1.027984e-20, 1.541976e-20, 
    5.139921e-21, 1.027984e-20, -2.569961e-20, -5.139921e-21, 0, 
    1.027984e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 2.055969e-20, -1.027984e-20, 2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, 1.541976e-20, -2.569961e-20, 
    2.006177e-36, -1.027984e-20, 1.027984e-20, 1.541976e-20, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -2.055969e-20, -1.027984e-20, 0, 
    1.027984e-20, -2.569961e-20, 0, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, 0, -2.055969e-20, 3.597945e-20, -1.027984e-20, 
    -1.027984e-20, 0, -2.055969e-20, 2.055969e-20, -1.541976e-20, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, -1.541976e-20, -2.006177e-36, 
    1.027984e-20, 2.055969e-20, 5.139921e-21, -2.006177e-36, -1.027984e-20, 
    2.006177e-36, 2.569961e-20, 0, 1.541976e-20, -2.055969e-20, 2.055969e-20, 
    2.006177e-36, -5.139921e-21, 1.541976e-20, 2.569961e-20, -1.541976e-20, 
    2.006177e-36, -1.541976e-20, 1.541976e-20, 2.569961e-20, 1.027984e-20, 
    -2.006177e-36, 5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 1.541976e-20, 1.541976e-20, 5.139921e-21, 2.055969e-20, 
    -2.006177e-36, 5.139921e-21, 1.541976e-20, -1.027984e-20, 2.055969e-20, 
    -1.541976e-20, -1.027984e-20, -1.541976e-20, 2.055969e-20, 2.055969e-20, 
    -1.541976e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, -2.006177e-36, 
    3.597945e-20, -1.541976e-20, 5.139921e-21, -2.055969e-20, -1.027984e-20, 
    -5.139921e-21, -2.569961e-20, 5.139921e-21, 5.139921e-21, 3.083953e-20, 
    1.027984e-20, 2.006177e-36, 1.027984e-20, 0, -1.541976e-20, 0, 
    1.541976e-20, 0, 3.083953e-20, -2.006177e-36, 2.006177e-36, 2.055969e-20, 
    2.055969e-20, 0, -3.083953e-20, -5.139921e-21, 1.541976e-20, 
    -1.541976e-20, -2.006177e-36, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -3.597945e-20, -4.111937e-20, -2.006177e-36, 1.027984e-20, 1.027984e-20, 
    1.027984e-20, -3.083953e-20, -1.541976e-20, 1.027984e-20, -2.055969e-20, 
    -1.541976e-20, 3.083953e-20, 1.027984e-20, 2.006177e-36, -5.139921e-21, 
    -2.055969e-20, -1.027984e-20, -2.006177e-36, -1.541976e-20, 0, 
    -2.569961e-20, 1.027984e-20, -1.541976e-20, 1.541976e-20, -2.055969e-20, 
    2.055969e-20, 0, 1.027984e-20, -5.139921e-20, 1.541976e-20, 2.569961e-20, 
    5.139921e-21, 5.139921e-21, -2.006177e-36, -1.027984e-20, -2.055969e-20, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, 1.541976e-20, 1.027984e-20, 
    -2.055969e-20, -1.027984e-20, 1.027984e-20, 0, 1.027984e-20, 
    -5.139921e-21, -2.055969e-20, 2.006177e-36, 1.027984e-20, 5.139921e-21, 
    -3.083953e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, -1.027984e-20, 
    1.541976e-20, -2.055969e-20, -5.139921e-21, 0, -1.027984e-20, 
    1.027984e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    4.111937e-20, 0, 1.027984e-20, -1.027984e-20, -2.055969e-20, 
    1.541976e-20, -5.139921e-21, 1.541976e-20, 5.139921e-21, 1.027984e-20, 
    -2.055969e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 0, 
    -1.027984e-20, -1.027984e-20, -1.027984e-20, 1.541976e-20, 2.055969e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -2.006177e-36, 1.541976e-20, 1.027984e-20, -1.541976e-20, 1.027984e-20, 
    0, -1.541976e-20, -2.055969e-20, -2.055969e-20, -2.006177e-36,
  2.006177e-36, -1.027984e-20, -2.006177e-36, 1.541976e-20, -2.055969e-20, 
    -1.027984e-20, 1.541976e-20, -5.139921e-21, 1.541976e-20, 4.111937e-20, 
    -3.597945e-20, -1.027984e-20, -3.083953e-20, -2.006177e-36, 1.541976e-20, 
    0, -1.027984e-20, 2.055969e-20, 2.055969e-20, 2.055969e-20, 
    -1.027984e-20, 1.027984e-20, 5.139921e-21, 2.006177e-36, 0, 
    -2.006177e-36, 5.139921e-21, -5.139921e-21, 5.139921e-21, 2.055969e-20, 
    2.569961e-20, 1.541976e-20, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    3.083953e-20, 1.027984e-20, 5.139921e-21, -2.569961e-20, -2.006177e-36, 
    2.055969e-20, 2.569961e-20, 2.569961e-20, 1.541976e-20, 5.139921e-21, 
    -3.083953e-20, -1.541976e-20, 1.027984e-20, 0, 1.027984e-20, 
    3.083953e-20, 5.139921e-21, -1.027984e-20, -3.083953e-20, 0, 
    1.541976e-20, 2.055969e-20, 1.027984e-20, 3.597945e-20, -2.055969e-20, 
    1.027984e-20, -5.139921e-21, -2.055969e-20, 0, 1.541976e-20, 
    -3.597945e-20, -5.139921e-21, -2.569961e-20, 0, -1.541976e-20, 
    1.027984e-20, 2.569961e-20, -1.541976e-20, -5.139921e-21, -5.139921e-21, 
    -2.055969e-20, -1.541976e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    4.111937e-20, -5.139921e-21, -1.541976e-20, 5.139921e-21, 1.027984e-20, 
    1.541976e-20, -2.055969e-20, 2.006177e-36, -1.541976e-20, 0, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 2.055969e-20, 
    1.027984e-20, -1.027984e-20, 1.027984e-20, 2.569961e-20, -1.027984e-20, 
    -3.083953e-20, 5.139921e-21, -5.139921e-21, 2.055969e-20, 4.111937e-20, 
    -3.597945e-20, -1.541976e-20, 1.541976e-20, 3.083953e-20, -5.139921e-21, 
    -1.027984e-20, 2.569961e-20, -1.027984e-20, 1.027984e-20, 0, 
    -1.027984e-20, 1.027984e-20, 5.139921e-21, 1.541976e-20, -2.569961e-20, 
    -1.027984e-20, 2.055969e-20, -2.006177e-36, 1.027984e-20, -1.541976e-20, 
    -5.139921e-21, 1.541976e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, 
    -2.569961e-20, -2.569961e-20, 5.139921e-21, -1.541976e-20, -3.597945e-20, 
    1.027984e-20, -2.055969e-20, 1.541976e-20, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, -4.111937e-20, 5.139921e-21, -1.027984e-20, -5.139921e-20, 
    -2.006177e-36, -5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -1.541976e-20, 2.055969e-20, -2.055969e-20, -3.083953e-20, -1.027984e-20, 
    -5.139921e-21, 2.569961e-20, -3.083953e-20, -5.139921e-21, 3.597945e-20, 
    -2.055969e-20, -1.027984e-20, -2.055969e-20, 1.027984e-20, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, 0, 
    1.541976e-20, 2.569961e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, 
    2.055969e-20, 2.055969e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, 1.027984e-20, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, -2.055969e-20, -2.006177e-36, -2.055969e-20, 1.541976e-20, 
    -5.139921e-21, 3.597945e-20, 1.027984e-20, 5.139921e-21, 2.569961e-20, 
    2.569961e-20, -2.055969e-20, -1.541976e-20, -5.139921e-21, 1.027984e-20, 
    -2.006177e-36, -1.541976e-20, 2.055969e-20, -1.027984e-20, 1.541976e-20, 
    1.541976e-20, 2.055969e-20, 5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -1.541976e-20, 5.139921e-21, -2.055969e-20, -2.055969e-20, -5.139921e-21, 
    0, -2.569961e-20, -5.139921e-21, 1.541976e-20, 2.569961e-20, 
    -2.055969e-20, 3.083953e-20, -2.055969e-20, 2.055969e-20, -1.541976e-20, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, -2.569961e-20, 3.083953e-20, 
    -2.569961e-20, -5.139921e-21, 0, -1.541976e-20, -1.027984e-20, 
    5.139921e-21, 2.569961e-20, 2.055969e-20, -5.139921e-21, -2.055969e-20, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, 1.541976e-20, -2.569961e-20, 
    1.541976e-20, -2.569961e-20, -5.139921e-21, 5.139921e-21, 0, 
    2.006177e-36, -5.139921e-21, 5.139921e-21, 2.569961e-20, -5.139921e-21, 
    3.083953e-20, 3.083953e-20, 1.541976e-20, 2.055969e-20, 1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 1.541976e-20, -2.006177e-36, 2.006177e-36, 
    0, -1.027984e-20, 1.027984e-20, 0, 1.541976e-20, 5.139921e-21, 
    -2.055969e-20, 0, 1.541976e-20, 5.139921e-21, 1.541976e-20, 
    -1.541976e-20, -1.541976e-20, 2.055969e-20, -1.541976e-20, -5.139921e-21, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, 2.055969e-20, -1.541976e-20, 
    1.027984e-20, -2.055969e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    1.541976e-20, -1.027984e-20, 1.541976e-20, 1.027984e-20, 1.027984e-20, 
    2.569961e-20, -3.083953e-20, -2.569961e-20, 0, 2.569961e-20, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, -1.541976e-20, -2.006177e-36, 
    2.055969e-20, 0, -5.139921e-21, 4.625929e-20, -5.139921e-21, 
    1.541976e-20, 1.027984e-20, 5.139921e-21, -2.569961e-20, 1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -1.027984e-20, 2.055969e-20, -1.541976e-20, 1.027984e-20, 
    5.139921e-21, -2.055969e-20,
  -5.139921e-21, -1.541976e-20, -1.027984e-20, 3.083953e-20, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, 0, 1.541976e-20, 
    -2.569961e-20, -1.541976e-20, -1.027984e-20, 1.027984e-20, -4.111937e-20, 
    -1.541976e-20, -5.139921e-21, -2.569961e-20, 5.139921e-21, -1.541976e-20, 
    -1.541976e-20, 1.027984e-20, 2.569961e-20, 4.111937e-20, 5.139921e-21, 
    2.006177e-36, 4.625929e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -2.055969e-20, -3.083953e-20, 1.541976e-20, -2.055969e-20, 
    2.569961e-20, 1.541976e-20, -5.139921e-21, 2.569961e-20, -1.541976e-20, 
    -1.541976e-20, 3.083953e-20, -1.027984e-20, -1.027984e-20, -4.625929e-20, 
    -5.139921e-21, 1.027984e-20, 2.055969e-20, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, -2.569961e-20, 1.541976e-20, 1.541976e-20, -1.541976e-20, 
    2.055969e-20, -2.055969e-20, 0, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 2.569961e-20, 5.139921e-21, -4.111937e-20, 5.139921e-21, 
    2.055969e-20, 5.139921e-20, -1.541976e-20, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -2.569961e-20, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -2.569961e-20, 5.139921e-21, -1.541976e-20, 
    -3.083953e-20, -1.541976e-20, 0, -5.139921e-21, 1.027984e-20, 
    -2.006177e-36, -2.569961e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, 3.083953e-20, 3.083953e-20, -5.139921e-21, 
    -2.006177e-36, -3.083953e-20, 2.055969e-20, 2.006177e-36, 1.027984e-20, 
    1.027984e-20, -1.027984e-20, 2.569961e-20, 0, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, -1.027984e-20, 3.083953e-20, -2.006177e-36, 
    0, 0, -1.027984e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, 
    -1.027984e-20, 1.541976e-20, -2.006177e-36, -3.083953e-20, 5.139921e-21, 
    -4.625929e-20, -1.541976e-20, -2.055969e-20, -1.027984e-20, 
    -5.139921e-20, -3.597945e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    2.569961e-20, 1.027984e-20, -6.681898e-20, -1.541976e-20, 0, 
    2.569961e-20, -1.027984e-20, 3.083953e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 0, 5.139921e-21, -4.625929e-20, 
    -5.139921e-20, 1.027984e-20, 0, 4.625929e-20, 1.541976e-20, 
    -5.139921e-21, -2.569961e-20, 3.083953e-20, -1.027984e-20, 2.055969e-20, 
    5.139921e-21, -2.055969e-20, -2.569961e-20, -1.541976e-20, 5.139921e-21, 
    2.569961e-20, 5.139921e-21, 1.027984e-20, 1.541976e-20, -1.027984e-20, 
    5.139921e-21, 2.006177e-36, -1.027984e-20, -3.597945e-20, -5.139921e-21, 
    -1.541976e-20, 0, -1.027984e-20, 5.139921e-21, -1.541976e-20, 
    -2.055969e-20, -3.083953e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, -1.541976e-20, 0, -5.139921e-21, 1.541976e-20, 
    -2.055969e-20, -2.055969e-20, -1.541976e-20, 3.083953e-20, 2.569961e-20, 
    3.083953e-20, -2.006177e-36, 1.027984e-20, -1.541976e-20, -2.055969e-20, 
    1.027984e-20, 2.055969e-20, -1.027984e-20, 1.027984e-20, -1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 3.083953e-20, -2.569961e-20, -1.541976e-20, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -5.139921e-21, 3.597945e-20, -3.083953e-20, 
    -2.006177e-36, 3.083953e-20, 5.139921e-21, 1.027984e-20, -2.569961e-20, 
    -2.006177e-36, -3.083953e-20, 1.541976e-20, 5.139921e-21, -2.006177e-36, 
    -2.055969e-20, 2.569961e-20, 2.055969e-20, -2.055969e-20, 1.541976e-20, 
    2.006177e-36, -1.541976e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    1.541976e-20, -2.569961e-20, 5.139921e-21, -1.541976e-20, 3.597945e-20, 
    5.139921e-21, 2.055969e-20, 0, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    -5.139921e-21, -2.055969e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, 2.055969e-20, 1.027984e-20, -2.055969e-20, -1.027984e-20, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, 
    -2.569961e-20, 2.006177e-36, -2.569961e-20, -3.083953e-20, -1.027984e-20, 
    1.541976e-20, -1.541976e-20, 1.541976e-20, -5.139921e-21, -3.597945e-20, 
    2.055969e-20, -4.625929e-20, -1.027984e-20, -5.139921e-21, 1.541976e-20, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, 2.006177e-36, 
    2.055969e-20, 5.139921e-21, -2.055969e-20, 2.006177e-36, -2.055969e-20, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, -2.569961e-20, -2.569961e-20, 
    1.541976e-20, -5.139921e-21, -1.027984e-20, 1.541976e-20, -4.625929e-20, 
    -3.083953e-20, 5.139921e-21, -2.569961e-20, 1.027984e-20, -2.569961e-20, 
    -5.139921e-21, 0, 0, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    5.139921e-21, -3.083953e-20, -5.139921e-21, 0, -1.027984e-20, 
    1.027984e-20, 1.027984e-20, 2.569961e-20, -5.139921e-21, 1.541976e-20, 
    5.139921e-21, 3.083953e-20, -2.569961e-20, 2.006177e-36, -1.027984e-20, 
    -5.139921e-21, 0, 3.597945e-20, -2.569961e-20, -1.541976e-20, 
    -2.569961e-20, 1.027984e-20, 3.597945e-20, -2.569961e-20, -1.541976e-20, 
    2.569961e-20, 1.541976e-20,
  -2.055969e-20, 4.111937e-20, 0, 1.027984e-20, -2.055969e-20, 0, 0, 
    2.055969e-20, 0, -5.139921e-21, 1.027984e-20, -3.083953e-20, 
    -1.541976e-20, 5.139921e-21, 1.027984e-20, 1.541976e-20, 1.541976e-20, 0, 
    -1.541976e-20, 5.139921e-21, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    1.541976e-20, 5.139921e-21, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    -1.541976e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 1.541976e-20, 
    3.083953e-20, -2.055969e-20, 1.027984e-20, 1.541976e-20, -2.055969e-20, 
    0, -5.139921e-21, -2.055969e-20, 0, 0, 5.139921e-21, -4.111937e-20, 
    5.139921e-21, 2.006177e-36, 5.139921e-21, -1.541976e-20, -1.541976e-20, 
    3.083953e-20, -2.569961e-20, 3.083953e-20, 5.139921e-21, 5.139921e-21, 
    5.653913e-20, 2.569961e-20, -5.139921e-21, -1.541976e-20, 2.569961e-20, 
    -3.083953e-20, -1.541976e-20, -2.055969e-20, -5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 1.027984e-20, 1.541976e-20, 1.027984e-20, 
    0, -1.027984e-20, -1.541976e-20, 5.139921e-21, 0, 5.139921e-21, 
    1.027984e-20, 0, 1.027984e-20, 1.541976e-20, 1.541976e-20, 1.027984e-20, 
    1.541976e-20, -1.027984e-20, -3.083953e-20, 0, 5.139921e-21, 0, 
    2.006177e-36, 2.569961e-20, -2.569961e-20, 2.006177e-36, 1.541976e-20, 0, 
    2.569961e-20, -2.055969e-20, -3.597945e-20, 5.139921e-21, 2.006177e-36, 
    0, -1.027984e-20, 5.139921e-21, -1.027984e-20, 1.541976e-20, 
    -3.597945e-20, 5.139921e-21, 2.569961e-20, 5.139921e-21, 1.541976e-20, 
    2.055969e-20, 2.055969e-20, 0, -5.139921e-21, 2.006177e-36, 
    -5.139921e-21, -5.139921e-21, 0, -5.139921e-21, -1.541976e-20, 
    2.569961e-20, 1.541976e-20, -2.055969e-20, 0, -2.055969e-20, 
    -1.541976e-20, 2.055969e-20, 2.006177e-36, -1.027984e-20, -1.541976e-20, 
    -2.006177e-36, -3.083953e-20, 1.027984e-20, -1.541976e-20, 2.055969e-20, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, 0, -2.055969e-20, 
    5.139921e-21, -2.055969e-20, -1.027984e-20, -5.139921e-21, -2.569961e-20, 
    -1.541976e-20, -1.027984e-20, 1.027984e-20, -2.055969e-20, -2.055969e-20, 
    1.541976e-20, 5.139921e-21, 1.541976e-20, -2.055969e-20, -2.055969e-20, 
    1.027984e-20, -1.541976e-20, 2.006177e-36, -5.139921e-21, 2.569961e-20, 
    5.139921e-21, 0, -2.055969e-20, -3.597945e-20, 0, 4.111937e-20, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    2.006177e-36, -5.139921e-21, -3.083953e-20, 4.625929e-20, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, -2.569961e-20, -4.625929e-20, 
    -2.569961e-20, -3.083953e-20, 1.027984e-20, 1.541976e-20, 2.006177e-36, 
    0, 5.139921e-21, 2.006177e-36, 3.083953e-20, -1.027984e-20, 
    -4.111937e-20, 1.027984e-20, 1.541976e-20, -1.541976e-20, 5.139921e-21, 
    5.139921e-21, 0, 1.541976e-20, 0, 5.139921e-21, 1.027984e-20, 
    -1.541976e-20, -2.569961e-20, 2.006177e-36, -1.541976e-20, 1.027984e-20, 
    -3.597945e-20, 0, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 2.055969e-20, 
    2.055969e-20, -5.139921e-21, 5.139921e-21, 2.569961e-20, 5.139921e-21, 
    -1.541976e-20, -1.027984e-20, -1.541976e-20, 3.083953e-20, 2.569961e-20, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -1.541976e-20, 1.027984e-20, 1.541976e-20, 5.139921e-21, 2.569961e-20, 
    5.139921e-21, -1.541976e-20, -1.541976e-20, 2.569961e-20, -2.006177e-36, 
    -2.569961e-20, -1.027984e-20, 2.569961e-20, 1.027984e-20, -1.027984e-20, 
    1.027984e-20, 4.111937e-20, 1.027984e-20, 5.139921e-21, -2.569961e-20, 0, 
    2.569961e-20, 0, 0, 2.055969e-20, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, -2.055969e-20, -1.541976e-20, -1.541976e-20, 5.139921e-21, 
    1.541976e-20, -2.006177e-36, 1.027984e-20, 1.027984e-20, -2.055969e-20, 
    -1.027984e-20, 4.625929e-20, 1.027984e-20, -1.027984e-20, 1.541976e-20, 
    -2.006177e-36, -2.006177e-36, 0, 1.027984e-20, -1.541976e-20, 
    1.541976e-20, 5.139921e-21, 2.055969e-20, 0, 1.027984e-20, -2.055969e-20, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, -2.055969e-20, 0, 
    -2.569961e-20, 1.027984e-20, -1.027984e-20, -5.139921e-20, 2.006177e-36, 
    -1.541976e-20, 0, -1.541976e-20, -5.139921e-21, 2.006177e-36, 
    -3.597945e-20, -2.006177e-36, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -2.055969e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-20, 3.597945e-20, 3.083953e-20, 2.055969e-20, 2.569961e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -3.083953e-20, 5.139921e-21, 1.541976e-20, -2.055969e-20, 5.139921e-21, 
    2.055969e-20, 1.541976e-20, -5.139921e-21, 3.083953e-20, -4.111937e-20, 
    4.111937e-20, 1.027984e-20, -2.055969e-20, -2.569961e-20, -2.055969e-20, 
    -5.139921e-21, 2.055969e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21,
  8.598663e-29, 8.598634e-29, 8.59864e-29, 8.598617e-29, 8.59863e-29, 
    8.598615e-29, 8.598657e-29, 8.598634e-29, 8.598649e-29, 8.598661e-29, 
    8.598572e-29, 8.598616e-29, 8.598527e-29, 8.598555e-29, 8.598485e-29, 
    8.598531e-29, 8.598475e-29, 8.598486e-29, 8.598453e-29, 8.598463e-29, 
    8.598421e-29, 8.598449e-29, 8.5984e-29, 8.598428e-29, 8.598424e-29, 
    8.59845e-29, 8.598607e-29, 8.598578e-29, 8.598609e-29, 8.598605e-29, 
    8.598607e-29, 8.59863e-29, 8.598641e-29, 8.598666e-29, 8.598661e-29, 
    8.598643e-29, 8.598603e-29, 8.598616e-29, 8.598582e-29, 8.598583e-29, 
    8.598545e-29, 8.598562e-29, 8.598497e-29, 8.598516e-29, 8.598462e-29, 
    8.598476e-29, 8.598463e-29, 8.598467e-29, 8.598463e-29, 8.598483e-29, 
    8.598474e-29, 8.598491e-29, 8.598559e-29, 8.598539e-29, 8.598598e-29, 
    8.598633e-29, 8.598657e-29, 8.598673e-29, 8.598671e-29, 8.598666e-29, 
    8.598643e-29, 8.598622e-29, 8.598605e-29, 8.598594e-29, 8.598583e-29, 
    8.59855e-29, 8.598533e-29, 8.598494e-29, 8.598501e-29, 8.598489e-29, 
    8.598477e-29, 8.598458e-29, 8.598461e-29, 8.598453e-29, 8.598489e-29, 
    8.598465e-29, 8.598504e-29, 8.598494e-29, 8.59858e-29, 8.598613e-29, 
    8.598627e-29, 8.598639e-29, 8.598669e-29, 8.598648e-29, 8.598657e-29, 
    8.598637e-29, 8.598625e-29, 8.598631e-29, 8.598593e-29, 8.598608e-29, 
    8.598532e-29, 8.598565e-29, 8.598479e-29, 8.598499e-29, 8.598474e-29, 
    8.598486e-29, 8.598464e-29, 8.598485e-29, 8.59845e-29, 8.598442e-29, 
    8.598447e-29, 8.598427e-29, 8.598485e-29, 8.598463e-29, 8.598631e-29, 
    8.59863e-29, 8.598625e-29, 8.598646e-29, 8.598647e-29, 8.598666e-29, 
    8.598649e-29, 8.598642e-29, 8.598624e-29, 8.598614e-29, 8.598604e-29, 
    8.598581e-29, 8.598557e-29, 8.598522e-29, 8.598498e-29, 8.598481e-29, 
    8.598491e-29, 8.598482e-29, 8.598492e-29, 8.598497e-29, 8.598445e-29, 
    8.598474e-29, 8.59843e-29, 8.598432e-29, 8.598453e-29, 8.598432e-29, 
    8.59863e-29, 8.598635e-29, 8.598655e-29, 8.598639e-29, 8.598668e-29, 
    8.598652e-29, 8.598643e-29, 8.598608e-29, 8.5986e-29, 8.598593e-29, 
    8.598579e-29, 8.598561e-29, 8.598529e-29, 8.598501e-29, 8.598477e-29, 
    8.598479e-29, 8.598478e-29, 8.598472e-29, 8.598486e-29, 8.59847e-29, 
    8.598467e-29, 8.598474e-29, 8.598433e-29, 8.598445e-29, 8.598432e-29, 
    8.59844e-29, 8.598633e-29, 8.598624e-29, 8.598629e-29, 8.598619e-29, 
    8.598626e-29, 8.598596e-29, 8.598586e-29, 8.598544e-29, 8.598562e-29, 
    8.598533e-29, 8.598559e-29, 8.598554e-29, 8.598533e-29, 8.598557e-29, 
    8.598503e-29, 8.59854e-29, 8.598472e-29, 8.598508e-29, 8.59847e-29, 
    8.598477e-29, 8.598465e-29, 8.598454e-29, 8.598441e-29, 8.598417e-29, 
    8.598423e-29, 8.598402e-29, 8.59861e-29, 8.598597e-29, 8.598598e-29, 
    8.598585e-29, 8.598575e-29, 8.598555e-29, 8.598521e-29, 8.598534e-29, 
    8.598511e-29, 8.598506e-29, 8.598541e-29, 8.598519e-29, 8.598589e-29, 
    8.598578e-29, 8.598584e-29, 8.598609e-29, 8.598531e-29, 8.598571e-29, 
    8.598497e-29, 8.598519e-29, 8.598456e-29, 8.598487e-29, 8.598426e-29, 
    8.598399e-29, 8.598374e-29, 8.598346e-29, 8.59859e-29, 8.598599e-29, 
    8.598584e-29, 8.598563e-29, 8.598544e-29, 8.598518e-29, 8.598515e-29, 
    8.59851e-29, 8.598498e-29, 8.598487e-29, 8.598509e-29, 8.598485e-29, 
    8.598575e-29, 8.598527e-29, 8.598602e-29, 8.59858e-29, 8.598564e-29, 
    8.598571e-29, 8.598535e-29, 8.598527e-29, 8.598493e-29, 8.59851e-29, 
    8.598406e-29, 8.598452e-29, 8.598323e-29, 8.598359e-29, 8.598602e-29, 
    8.59859e-29, 8.598551e-29, 8.598569e-29, 8.598516e-29, 8.598503e-29, 
    8.598492e-29, 8.598478e-29, 8.598477e-29, 8.598468e-29, 8.598482e-29, 
    8.598469e-29, 8.598518e-29, 8.598496e-29, 8.598556e-29, 8.598541e-29, 
    8.598548e-29, 8.598555e-29, 8.598532e-29, 8.598508e-29, 8.598507e-29, 
    8.5985e-29, 8.598479e-29, 8.598516e-29, 8.5984e-29, 8.598471e-29, 
    8.598578e-29, 8.598556e-29, 8.598553e-29, 8.598562e-29, 8.598504e-29, 
    8.598525e-29, 8.598468e-29, 8.598484e-29, 8.598459e-29, 8.598471e-29, 
    8.598473e-29, 8.598489e-29, 8.598499e-29, 8.598524e-29, 8.598544e-29, 
    8.59856e-29, 8.598557e-29, 8.598539e-29, 8.598507e-29, 8.598476e-29, 
    8.598483e-29, 8.59846e-29, 8.598519e-29, 8.598495e-29, 8.598504e-29, 
    8.59848e-29, 8.598535e-29, 8.598488e-29, 8.598546e-29, 8.598541e-29, 
    8.598525e-29, 8.598494e-29, 8.598486e-29, 8.598479e-29, 8.598483e-29, 
    8.598506e-29, 8.59851e-29, 8.598525e-29, 8.59853e-29, 8.598542e-29, 
    8.598552e-29, 8.598543e-29, 8.598533e-29, 8.598506e-29, 8.598481e-29, 
    8.598454e-29, 8.598448e-29, 8.598416e-29, 8.598442e-29, 8.5984e-29, 
    8.598435e-29, 8.598373e-29, 8.598485e-29, 8.598436e-29, 8.598524e-29, 
    8.598515e-29, 8.598498e-29, 8.598459e-29, 8.59848e-29, 8.598455e-29, 
    8.59851e-29, 8.598538e-29, 8.598545e-29, 8.598559e-29, 8.598545e-29, 
    8.598547e-29, 8.598533e-29, 8.598538e-29, 8.598505e-29, 8.598522e-29, 
    8.598473e-29, 8.598455e-29, 8.598405e-29, 8.598373e-29, 8.598341e-29, 
    8.598327e-29, 8.598323e-29, 8.598321e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.165244e-08, 1.170366e-08, 1.16937e-08, 1.173501e-08, 1.171209e-08, 
    1.173914e-08, 1.166282e-08, 1.170569e-08, 1.167832e-08, 1.165705e-08, 
    1.181518e-08, 1.173685e-08, 1.189654e-08, 1.184658e-08, 1.197206e-08, 
    1.188876e-08, 1.198886e-08, 1.196966e-08, 1.202744e-08, 1.201089e-08, 
    1.20848e-08, 1.203508e-08, 1.212312e-08, 1.207293e-08, 1.208078e-08, 
    1.203345e-08, 1.175262e-08, 1.180543e-08, 1.174949e-08, 1.175702e-08, 
    1.175364e-08, 1.171257e-08, 1.169187e-08, 1.164852e-08, 1.165639e-08, 
    1.168823e-08, 1.17604e-08, 1.17359e-08, 1.179765e-08, 1.179625e-08, 
    1.186499e-08, 1.1834e-08, 1.194953e-08, 1.19167e-08, 1.201158e-08, 
    1.198772e-08, 1.201046e-08, 1.200356e-08, 1.201055e-08, 1.197555e-08, 
    1.199055e-08, 1.195975e-08, 1.183981e-08, 1.187506e-08, 1.176992e-08, 
    1.17067e-08, 1.16647e-08, 1.16349e-08, 1.163911e-08, 1.164715e-08, 
    1.168842e-08, 1.172722e-08, 1.175679e-08, 1.177657e-08, 1.179605e-08, 
    1.185505e-08, 1.188627e-08, 1.195617e-08, 1.194356e-08, 1.196493e-08, 
    1.198535e-08, 1.201962e-08, 1.201398e-08, 1.202908e-08, 1.196436e-08, 
    1.200738e-08, 1.193637e-08, 1.195579e-08, 1.180136e-08, 1.174251e-08, 
    1.171751e-08, 1.169561e-08, 1.164235e-08, 1.167913e-08, 1.166464e-08, 
    1.169913e-08, 1.172105e-08, 1.171021e-08, 1.177711e-08, 1.17511e-08, 
    1.188812e-08, 1.18291e-08, 1.198296e-08, 1.194615e-08, 1.199179e-08, 
    1.19685e-08, 1.200841e-08, 1.197249e-08, 1.20347e-08, 1.204825e-08, 
    1.203899e-08, 1.207456e-08, 1.19705e-08, 1.201046e-08, 1.17099e-08, 
    1.171167e-08, 1.171991e-08, 1.16837e-08, 1.168149e-08, 1.164831e-08, 
    1.167783e-08, 1.16904e-08, 1.172232e-08, 1.174119e-08, 1.175914e-08, 
    1.179859e-08, 1.184266e-08, 1.190427e-08, 1.194853e-08, 1.19782e-08, 
    1.196001e-08, 1.197607e-08, 1.195812e-08, 1.19497e-08, 1.204318e-08, 
    1.199069e-08, 1.206944e-08, 1.206508e-08, 1.202944e-08, 1.206558e-08, 
    1.171291e-08, 1.170274e-08, 1.166741e-08, 1.169506e-08, 1.164469e-08, 
    1.167289e-08, 1.16891e-08, 1.175164e-08, 1.176538e-08, 1.177813e-08, 
    1.180329e-08, 1.183559e-08, 1.189224e-08, 1.194153e-08, 1.198653e-08, 
    1.198324e-08, 1.19844e-08, 1.199445e-08, 1.196955e-08, 1.199854e-08, 
    1.20034e-08, 1.199068e-08, 1.20645e-08, 1.204341e-08, 1.206499e-08, 
    1.205126e-08, 1.170604e-08, 1.172316e-08, 1.171391e-08, 1.173131e-08, 
    1.171905e-08, 1.177354e-08, 1.178988e-08, 1.186632e-08, 1.183495e-08, 
    1.188488e-08, 1.184002e-08, 1.184797e-08, 1.188651e-08, 1.184245e-08, 
    1.193882e-08, 1.187348e-08, 1.199484e-08, 1.19296e-08, 1.199893e-08, 
    1.198634e-08, 1.200718e-08, 1.202585e-08, 1.204934e-08, 1.209267e-08, 
    1.208264e-08, 1.211888e-08, 1.174868e-08, 1.177089e-08, 1.176893e-08, 
    1.179217e-08, 1.180935e-08, 1.18466e-08, 1.190633e-08, 1.188387e-08, 
    1.192511e-08, 1.193338e-08, 1.187073e-08, 1.19092e-08, 1.178575e-08, 
    1.180569e-08, 1.179382e-08, 1.175044e-08, 1.188905e-08, 1.181791e-08, 
    1.194926e-08, 1.191073e-08, 1.202319e-08, 1.196726e-08, 1.207711e-08, 
    1.212408e-08, 1.216827e-08, 1.221992e-08, 1.1783e-08, 1.176792e-08, 
    1.179493e-08, 1.183231e-08, 1.186698e-08, 1.191308e-08, 1.19178e-08, 
    1.192643e-08, 1.19488e-08, 1.196761e-08, 1.192916e-08, 1.197233e-08, 
    1.181032e-08, 1.189522e-08, 1.176221e-08, 1.180227e-08, 1.18301e-08, 
    1.181789e-08, 1.18813e-08, 1.189625e-08, 1.195698e-08, 1.192558e-08, 
    1.211249e-08, 1.20298e-08, 1.225925e-08, 1.219513e-08, 1.176265e-08, 
    1.178295e-08, 1.185362e-08, 1.182e-08, 1.191616e-08, 1.193983e-08, 
    1.195907e-08, 1.198366e-08, 1.198632e-08, 1.200089e-08, 1.197701e-08, 
    1.199995e-08, 1.191318e-08, 1.195195e-08, 1.184554e-08, 1.187144e-08, 
    1.185953e-08, 1.184646e-08, 1.18868e-08, 1.192977e-08, 1.193069e-08, 
    1.194447e-08, 1.19833e-08, 1.191655e-08, 1.212316e-08, 1.199557e-08, 
    1.180509e-08, 1.184421e-08, 1.184979e-08, 1.183464e-08, 1.193745e-08, 
    1.19002e-08, 1.200054e-08, 1.197342e-08, 1.201785e-08, 1.199577e-08, 
    1.199252e-08, 1.196417e-08, 1.194651e-08, 1.190191e-08, 1.186562e-08, 
    1.183684e-08, 1.184353e-08, 1.187514e-08, 1.19324e-08, 1.198656e-08, 
    1.19747e-08, 1.201447e-08, 1.190918e-08, 1.195333e-08, 1.193627e-08, 
    1.198076e-08, 1.188327e-08, 1.19663e-08, 1.186205e-08, 1.187119e-08, 
    1.189946e-08, 1.195633e-08, 1.196891e-08, 1.198234e-08, 1.197405e-08, 
    1.193385e-08, 1.192726e-08, 1.189877e-08, 1.189091e-08, 1.18692e-08, 
    1.185123e-08, 1.186765e-08, 1.188489e-08, 1.193387e-08, 1.1978e-08, 
    1.202612e-08, 1.203789e-08, 1.209412e-08, 1.204835e-08, 1.212387e-08, 
    1.205967e-08, 1.217081e-08, 1.19711e-08, 1.205778e-08, 1.190075e-08, 
    1.191767e-08, 1.194826e-08, 1.201844e-08, 1.198055e-08, 1.202486e-08, 
    1.192701e-08, 1.187624e-08, 1.18631e-08, 1.183859e-08, 1.186366e-08, 
    1.186162e-08, 1.188561e-08, 1.18779e-08, 1.193549e-08, 1.190456e-08, 
    1.199244e-08, 1.202451e-08, 1.211508e-08, 1.21706e-08, 1.222712e-08, 
    1.225207e-08, 1.225966e-08, 1.226284e-08 ;

 SOIL1N_TO_SOIL3N =
  1.382522e-10, 1.388602e-10, 1.38742e-10, 1.392323e-10, 1.389603e-10, 
    1.392814e-10, 1.383755e-10, 1.388843e-10, 1.385595e-10, 1.38307e-10, 
    1.401839e-10, 1.392542e-10, 1.411496e-10, 1.405566e-10, 1.42046e-10, 
    1.410573e-10, 1.422454e-10, 1.420175e-10, 1.427034e-10, 1.425069e-10, 
    1.433842e-10, 1.427941e-10, 1.43839e-10, 1.432433e-10, 1.433365e-10, 
    1.427746e-10, 1.394413e-10, 1.400682e-10, 1.394041e-10, 1.394935e-10, 
    1.394534e-10, 1.389659e-10, 1.387203e-10, 1.382058e-10, 1.382992e-10, 
    1.386771e-10, 1.395337e-10, 1.392429e-10, 1.399758e-10, 1.399592e-10, 
    1.407751e-10, 1.404073e-10, 1.417786e-10, 1.413888e-10, 1.425151e-10, 
    1.422319e-10, 1.425018e-10, 1.424199e-10, 1.425029e-10, 1.420875e-10, 
    1.422654e-10, 1.418999e-10, 1.404762e-10, 1.408946e-10, 1.396466e-10, 
    1.388963e-10, 1.383978e-10, 1.380441e-10, 1.380941e-10, 1.381894e-10, 
    1.386793e-10, 1.391398e-10, 1.394908e-10, 1.397255e-10, 1.399569e-10, 
    1.406571e-10, 1.410276e-10, 1.418574e-10, 1.417076e-10, 1.419613e-10, 
    1.422037e-10, 1.426106e-10, 1.425436e-10, 1.427229e-10, 1.419546e-10, 
    1.424652e-10, 1.416223e-10, 1.418529e-10, 1.400198e-10, 1.393214e-10, 
    1.390246e-10, 1.387647e-10, 1.381326e-10, 1.385691e-10, 1.38397e-10, 
    1.388064e-10, 1.390666e-10, 1.389379e-10, 1.39732e-10, 1.394233e-10, 
    1.410496e-10, 1.403491e-10, 1.421754e-10, 1.417384e-10, 1.422802e-10, 
    1.420037e-10, 1.424774e-10, 1.420511e-10, 1.427896e-10, 1.429504e-10, 
    1.428405e-10, 1.432626e-10, 1.420274e-10, 1.425018e-10, 1.389343e-10, 
    1.389553e-10, 1.39053e-10, 1.386233e-10, 1.38597e-10, 1.382032e-10, 
    1.385536e-10, 1.387028e-10, 1.390816e-10, 1.393057e-10, 1.395187e-10, 
    1.39987e-10, 1.4051e-10, 1.412413e-10, 1.417667e-10, 1.421189e-10, 
    1.419029e-10, 1.420936e-10, 1.418805e-10, 1.417806e-10, 1.428901e-10, 
    1.422671e-10, 1.432019e-10, 1.431502e-10, 1.427271e-10, 1.43156e-10, 
    1.3897e-10, 1.388493e-10, 1.3843e-10, 1.387581e-10, 1.381603e-10, 
    1.384949e-10, 1.386874e-10, 1.394297e-10, 1.395928e-10, 1.39744e-10, 
    1.400427e-10, 1.404261e-10, 1.410986e-10, 1.416837e-10, 1.422178e-10, 
    1.421786e-10, 1.421924e-10, 1.423117e-10, 1.420162e-10, 1.423603e-10, 
    1.42418e-10, 1.42267e-10, 1.431432e-10, 1.428929e-10, 1.431491e-10, 
    1.429861e-10, 1.388885e-10, 1.390917e-10, 1.389819e-10, 1.391884e-10, 
    1.390429e-10, 1.396897e-10, 1.398836e-10, 1.407909e-10, 1.404186e-10, 
    1.410112e-10, 1.404787e-10, 1.405731e-10, 1.410305e-10, 1.405075e-10, 
    1.416514e-10, 1.408759e-10, 1.423164e-10, 1.41542e-10, 1.423649e-10, 
    1.422155e-10, 1.424629e-10, 1.426845e-10, 1.429633e-10, 1.434777e-10, 
    1.433585e-10, 1.437887e-10, 1.393946e-10, 1.396581e-10, 1.396349e-10, 
    1.399107e-10, 1.401147e-10, 1.405568e-10, 1.412658e-10, 1.409992e-10, 
    1.414887e-10, 1.415869e-10, 1.408433e-10, 1.412999e-10, 1.398345e-10, 
    1.400713e-10, 1.399303e-10, 1.394154e-10, 1.410606e-10, 1.402163e-10, 
    1.417754e-10, 1.41318e-10, 1.426529e-10, 1.41989e-10, 1.43293e-10, 
    1.438504e-10, 1.44375e-10, 1.449882e-10, 1.39802e-10, 1.396229e-10, 
    1.399435e-10, 1.403871e-10, 1.407987e-10, 1.413459e-10, 1.414019e-10, 
    1.415044e-10, 1.417699e-10, 1.419932e-10, 1.415368e-10, 1.420491e-10, 
    1.401262e-10, 1.411339e-10, 1.395552e-10, 1.400306e-10, 1.40361e-10, 
    1.40216e-10, 1.409687e-10, 1.411461e-10, 1.418669e-10, 1.414943e-10, 
    1.437129e-10, 1.427313e-10, 1.45455e-10, 1.446938e-10, 1.395603e-10, 
    1.398013e-10, 1.406402e-10, 1.402411e-10, 1.413824e-10, 1.416634e-10, 
    1.418917e-10, 1.421837e-10, 1.422152e-10, 1.423882e-10, 1.421047e-10, 
    1.42377e-10, 1.413471e-10, 1.418073e-10, 1.405443e-10, 1.408517e-10, 
    1.407103e-10, 1.405551e-10, 1.410339e-10, 1.41544e-10, 1.415549e-10, 
    1.417184e-10, 1.421794e-10, 1.41387e-10, 1.438396e-10, 1.42325e-10, 
    1.400642e-10, 1.405284e-10, 1.405947e-10, 1.404149e-10, 1.416352e-10, 
    1.41193e-10, 1.42384e-10, 1.420621e-10, 1.425895e-10, 1.423274e-10, 
    1.422889e-10, 1.419523e-10, 1.417427e-10, 1.412133e-10, 1.407825e-10, 
    1.40441e-10, 1.405204e-10, 1.408956e-10, 1.415752e-10, 1.422181e-10, 
    1.420773e-10, 1.425494e-10, 1.412997e-10, 1.418237e-10, 1.416212e-10, 
    1.421493e-10, 1.409921e-10, 1.419776e-10, 1.407402e-10, 1.408487e-10, 
    1.411843e-10, 1.418593e-10, 1.420086e-10, 1.42168e-10, 1.420696e-10, 
    1.415924e-10, 1.415143e-10, 1.411761e-10, 1.410827e-10, 1.408251e-10, 
    1.406117e-10, 1.408066e-10, 1.410113e-10, 1.415926e-10, 1.421165e-10, 
    1.426876e-10, 1.428274e-10, 1.434948e-10, 1.429515e-10, 1.43848e-10, 
    1.430859e-10, 1.444052e-10, 1.420346e-10, 1.430634e-10, 1.411995e-10, 
    1.414003e-10, 1.417635e-10, 1.425965e-10, 1.421468e-10, 1.426727e-10, 
    1.415112e-10, 1.409086e-10, 1.407526e-10, 1.404617e-10, 1.407593e-10, 
    1.407351e-10, 1.410198e-10, 1.409283e-10, 1.416119e-10, 1.412447e-10, 
    1.422879e-10, 1.426686e-10, 1.437437e-10, 1.444027e-10, 1.450736e-10, 
    1.453697e-10, 1.454599e-10, 1.454976e-10 ;

 SOIL1N_vr =
  2.497422, 2.497415, 2.497416, 2.497411, 2.497414, 2.49741, 2.49742, 
    2.497415, 2.497418, 2.497421, 2.497401, 2.497411, 2.49739, 2.497396, 
    2.49738, 2.497391, 2.497378, 2.49738, 2.497373, 2.497375, 2.497365, 
    2.497372, 2.49736, 2.497367, 2.497366, 2.497372, 2.497409, 2.497402, 
    2.497409, 2.497408, 2.497408, 2.497414, 2.497416, 2.497422, 2.497421, 
    2.497417, 2.497408, 2.497411, 2.497403, 2.497403, 2.497394, 2.497398, 
    2.497383, 2.497387, 2.497375, 2.497378, 2.497375, 2.497376, 2.497375, 
    2.49738, 2.497377, 2.497381, 2.497397, 2.497393, 2.497406, 2.497415, 
    2.49742, 2.497424, 2.497423, 2.497422, 2.497417, 2.497412, 2.497408, 
    2.497406, 2.497403, 2.497395, 2.497391, 2.497382, 2.497384, 2.497381, 
    2.497378, 2.497374, 2.497375, 2.497372, 2.497381, 2.497375, 2.497385, 
    2.497382, 2.497402, 2.49741, 2.497413, 2.497416, 2.497423, 2.497418, 
    2.49742, 2.497416, 2.497413, 2.497414, 2.497406, 2.497409, 2.497391, 
    2.497399, 2.497379, 2.497383, 2.497377, 2.49738, 2.497375, 2.49738, 
    2.497372, 2.49737, 2.497371, 2.497367, 2.49738, 2.497375, 2.497414, 
    2.497414, 2.497413, 2.497418, 2.497418, 2.497422, 2.497418, 2.497417, 
    2.497413, 2.49741, 2.497408, 2.497403, 2.497397, 2.497389, 2.497383, 
    2.497379, 2.497381, 2.497379, 2.497382, 2.497383, 2.497371, 2.497377, 
    2.497367, 2.497368, 2.497372, 2.497368, 2.497414, 2.497415, 2.49742, 
    2.497416, 2.497423, 2.497419, 2.497417, 2.497409, 2.497407, 2.497405, 
    2.497402, 2.497398, 2.49739, 2.497384, 2.497378, 2.497378, 2.497378, 
    2.497377, 2.49738, 2.497376, 2.497376, 2.497377, 2.497368, 2.497371, 
    2.497368, 2.49737, 2.497415, 2.497412, 2.497414, 2.497411, 2.497413, 
    2.497406, 2.497404, 2.497394, 2.497398, 2.497391, 2.497397, 2.497396, 
    2.497391, 2.497397, 2.497384, 2.497393, 2.497377, 2.497386, 2.497376, 
    2.497378, 2.497375, 2.497373, 2.49737, 2.497364, 2.497365, 2.497361, 
    2.497409, 2.497406, 2.497406, 2.497403, 2.497401, 2.497396, 2.497389, 
    2.497391, 2.497386, 2.497385, 2.497393, 2.497388, 2.497404, 2.497402, 
    2.497403, 2.497409, 2.497391, 2.4974, 2.497383, 2.497388, 2.497373, 
    2.49738, 2.497366, 2.49736, 2.497355, 2.497348, 2.497405, 2.497407, 
    2.497403, 2.497398, 2.497394, 2.497388, 2.497387, 2.497386, 2.497383, 
    2.49738, 2.497386, 2.49738, 2.497401, 2.49739, 2.497407, 2.497402, 
    2.497398, 2.4974, 2.497392, 2.49739, 2.497382, 2.497386, 2.497362, 
    2.497372, 2.497343, 2.497351, 2.497407, 2.497405, 2.497395, 2.4974, 
    2.497387, 2.497384, 2.497382, 2.497378, 2.497378, 2.497376, 2.497379, 
    2.497376, 2.497388, 2.497383, 2.497396, 2.497393, 2.497395, 2.497396, 
    2.497391, 2.497386, 2.497385, 2.497384, 2.497378, 2.497387, 2.49736, 
    2.497377, 2.497402, 2.497397, 2.497396, 2.497398, 2.497385, 2.497389, 
    2.497376, 2.49738, 2.497374, 2.497377, 2.497377, 2.497381, 2.497383, 
    2.497389, 2.497394, 2.497398, 2.497397, 2.497393, 2.497385, 2.497378, 
    2.49738, 2.497374, 2.497388, 2.497382, 2.497385, 2.497379, 2.497391, 
    2.497381, 2.497394, 2.497393, 2.497389, 2.497382, 2.49738, 2.497379, 
    2.49738, 2.497385, 2.497386, 2.49739, 2.497391, 2.497393, 2.497396, 
    2.497394, 2.497391, 2.497385, 2.497379, 2.497373, 2.497371, 2.497364, 
    2.49737, 2.49736, 2.497369, 2.497354, 2.49738, 2.497369, 2.497389, 
    2.497387, 2.497383, 2.497374, 2.497379, 2.497373, 2.497386, 2.497392, 
    2.497394, 2.497397, 2.497394, 2.497394, 2.497391, 2.497392, 2.497385, 
    2.497389, 2.497377, 2.497373, 2.497361, 2.497354, 2.497347, 2.497344, 
    2.497343, 2.497342,
  2.497625, 2.497616, 2.497617, 2.49761, 2.497614, 2.49761, 2.497623, 
    2.497615, 2.49762, 2.497624, 2.497597, 2.49761, 2.497582, 2.497591, 
    2.497569, 2.497584, 2.497566, 2.49757, 2.49756, 2.497563, 2.49755, 
    2.497558, 2.497543, 2.497552, 2.49755, 2.497559, 2.497607, 2.497598, 
    2.497608, 2.497607, 2.497607, 2.497614, 2.497618, 2.497625, 2.497624, 
    2.497618, 2.497606, 2.49761, 2.497599, 2.4976, 2.497588, 2.497593, 
    2.497573, 2.497579, 2.497562, 2.497567, 2.497563, 2.497564, 2.497563, 
    2.497569, 2.497566, 2.497571, 2.497592, 2.497586, 2.497604, 2.497615, 
    2.497622, 2.497628, 2.497627, 2.497626, 2.497618, 2.497612, 2.497607, 
    2.497603, 2.4976, 2.49759, 2.497584, 2.497572, 2.497574, 2.497571, 
    2.497567, 2.497561, 2.497562, 2.49756, 2.497571, 2.497563, 2.497576, 
    2.497572, 2.497599, 2.497609, 2.497613, 2.497617, 2.497626, 2.49762, 
    2.497622, 2.497617, 2.497613, 2.497615, 2.497603, 2.497607, 2.497584, 
    2.497594, 2.497567, 2.497574, 2.497566, 2.49757, 2.497563, 2.497569, 
    2.497559, 2.497556, 2.497558, 2.497552, 2.49757, 2.497563, 2.497615, 
    2.497614, 2.497613, 2.497619, 2.49762, 2.497625, 2.49762, 2.497618, 
    2.497612, 2.497609, 2.497606, 2.497599, 2.497592, 2.497581, 2.497573, 
    2.497568, 2.497571, 2.497569, 2.497572, 2.497573, 2.497557, 2.497566, 
    2.497553, 2.497553, 2.497559, 2.497553, 2.497614, 2.497616, 2.497622, 
    2.497617, 2.497626, 2.497621, 2.497618, 2.497607, 2.497605, 2.497603, 
    2.497598, 2.497593, 2.497583, 2.497575, 2.497567, 2.497567, 2.497567, 
    2.497566, 2.49757, 2.497565, 2.497564, 2.497566, 2.497553, 2.497557, 
    2.497553, 2.497556, 2.497615, 2.497612, 2.497614, 2.497611, 2.497613, 
    2.497604, 2.497601, 2.497587, 2.497593, 2.497584, 2.497592, 2.497591, 
    2.497584, 2.497592, 2.497575, 2.497586, 2.497565, 2.497577, 2.497565, 
    2.497567, 2.497563, 2.49756, 2.497556, 2.497549, 2.49755, 2.497544, 
    2.497608, 2.497604, 2.497604, 2.4976, 2.497597, 2.497591, 2.497581, 
    2.497585, 2.497577, 2.497576, 2.497587, 2.49758, 2.497602, 2.497598, 
    2.4976, 2.497608, 2.497584, 2.497596, 2.497573, 2.49758, 2.497561, 
    2.49757, 2.497551, 2.497543, 2.497535, 2.497527, 2.497602, 2.497605, 
    2.4976, 2.497593, 2.497587, 2.49758, 2.497579, 2.497577, 2.497573, 
    2.49757, 2.497577, 2.497569, 2.497597, 2.497583, 2.497606, 2.497599, 
    2.497594, 2.497596, 2.497585, 2.497582, 2.497572, 2.497577, 2.497545, 
    2.497559, 2.49752, 2.497531, 2.497606, 2.497602, 2.49759, 2.497596, 
    2.497579, 2.497575, 2.497571, 2.497567, 2.497567, 2.497564, 2.497568, 
    2.497565, 2.49758, 2.497573, 2.497591, 2.497587, 2.497589, 2.497591, 
    2.497584, 2.497577, 2.497576, 2.497574, 2.497567, 2.497579, 2.497543, 
    2.497565, 2.497598, 2.497591, 2.49759, 2.497593, 2.497575, 2.497582, 
    2.497564, 2.497569, 2.497561, 2.497565, 2.497566, 2.497571, 2.497574, 
    2.497581, 2.497588, 2.497593, 2.497591, 2.497586, 2.497576, 2.497567, 
    2.497569, 2.497562, 2.49758, 2.497572, 2.497576, 2.497568, 2.497585, 
    2.49757, 2.497588, 2.497587, 2.497582, 2.497572, 2.49757, 2.497567, 
    2.497569, 2.497576, 2.497577, 2.497582, 2.497583, 2.497587, 2.49759, 
    2.497587, 2.497584, 2.497576, 2.497568, 2.49756, 2.497558, 2.497548, 
    2.497556, 2.497543, 2.497554, 2.497535, 2.49757, 2.497555, 2.497582, 
    2.497579, 2.497573, 2.497561, 2.497568, 2.49756, 2.497577, 2.497586, 
    2.497588, 2.497592, 2.497588, 2.497588, 2.497584, 2.497586, 2.497576, 
    2.497581, 2.497566, 2.49756, 2.497545, 2.497535, 2.497525, 2.497521, 
    2.49752, 2.497519,
  2.49784, 2.497831, 2.497833, 2.497825, 2.497829, 2.497824, 2.497838, 
    2.49783, 2.497835, 2.497839, 2.49781, 2.497825, 2.497795, 2.497804, 
    2.497781, 2.497797, 2.497778, 2.497782, 2.497771, 2.497774, 2.497761, 
    2.49777, 2.497753, 2.497763, 2.497761, 2.49777, 2.497822, 2.497812, 
    2.497822, 2.497821, 2.497822, 2.497829, 2.497833, 2.497841, 2.497839, 
    2.497834, 2.49782, 2.497825, 2.497813, 2.497814, 2.497801, 2.497807, 
    2.497785, 2.497792, 2.497774, 2.497778, 2.497774, 2.497776, 2.497774, 
    2.497781, 2.497778, 2.497783, 2.497806, 2.497799, 2.497818, 2.49783, 
    2.497838, 2.497844, 2.497843, 2.497841, 2.497834, 2.497826, 2.497821, 
    2.497817, 2.497814, 2.497803, 2.497797, 2.497784, 2.497787, 2.497782, 
    2.497779, 2.497772, 2.497774, 2.497771, 2.497783, 2.497775, 2.497788, 
    2.497784, 2.497813, 2.497824, 2.497828, 2.497832, 2.497842, 2.497835, 
    2.497838, 2.497832, 2.497828, 2.49783, 2.497817, 2.497822, 2.497797, 
    2.497808, 2.497779, 2.497786, 2.497778, 2.497782, 2.497775, 2.497781, 
    2.49777, 2.497767, 2.497769, 2.497762, 2.497782, 2.497774, 2.49783, 
    2.497829, 2.497828, 2.497834, 2.497835, 2.497841, 2.497836, 2.497833, 
    2.497827, 2.497824, 2.497821, 2.497813, 2.497805, 2.497794, 2.497786, 
    2.49778, 2.497783, 2.497781, 2.497784, 2.497785, 2.497768, 2.497778, 
    2.497763, 2.497764, 2.497771, 2.497764, 2.497829, 2.497831, 2.497838, 
    2.497832, 2.497842, 2.497837, 2.497833, 2.497822, 2.497819, 2.497817, 
    2.497812, 2.497806, 2.497796, 2.497787, 2.497779, 2.497779, 2.497779, 
    2.497777, 2.497782, 2.497776, 2.497776, 2.497778, 2.497764, 2.497768, 
    2.497764, 2.497767, 2.49783, 2.497827, 2.497829, 2.497826, 2.497828, 
    2.497818, 2.497815, 2.497801, 2.497807, 2.497797, 2.497806, 2.497804, 
    2.497797, 2.497805, 2.497787, 2.497799, 2.497777, 2.497789, 2.497776, 
    2.497779, 2.497775, 2.497771, 2.497767, 2.497759, 2.497761, 2.497754, 
    2.497823, 2.497818, 2.497819, 2.497814, 2.497811, 2.497804, 2.497793, 
    2.497797, 2.49779, 2.497788, 2.4978, 2.497793, 2.497816, 2.497812, 
    2.497814, 2.497822, 2.497797, 2.49781, 2.497786, 2.497792, 2.497772, 
    2.497782, 2.497762, 2.497753, 2.497745, 2.497736, 2.497816, 2.497819, 
    2.497814, 2.497807, 2.497801, 2.497792, 2.497791, 2.49779, 2.497786, 
    2.497782, 2.497789, 2.497781, 2.497811, 2.497795, 2.49782, 2.497813, 
    2.497808, 2.49781, 2.497798, 2.497795, 2.497784, 2.49779, 2.497756, 
    2.497771, 2.497729, 2.49774, 2.49782, 2.497816, 2.497803, 2.497809, 
    2.497792, 2.497787, 2.497784, 2.497779, 2.497779, 2.497776, 2.49778, 
    2.497776, 2.497792, 2.497785, 2.497805, 2.4978, 2.497802, 2.497804, 
    2.497797, 2.497789, 2.497789, 2.497786, 2.497779, 2.497792, 2.497753, 
    2.497777, 2.497812, 2.497805, 2.497804, 2.497807, 2.497788, 2.497794, 
    2.497776, 2.497781, 2.497773, 2.497777, 2.497777, 2.497783, 2.497786, 
    2.497794, 2.497801, 2.497806, 2.497805, 2.497799, 2.497789, 2.497779, 
    2.497781, 2.497773, 2.497793, 2.497785, 2.497788, 2.49778, 2.497798, 
    2.497782, 2.497802, 2.4978, 2.497795, 2.497784, 2.497782, 2.497779, 
    2.497781, 2.497788, 2.49779, 2.497795, 2.497796, 2.4978, 2.497803, 
    2.497801, 2.497797, 2.497788, 2.49778, 2.497771, 2.497769, 2.497759, 
    2.497767, 2.497753, 2.497765, 2.497745, 2.497782, 2.497766, 2.497794, 
    2.497791, 2.497786, 2.497773, 2.49778, 2.497772, 2.49779, 2.497799, 
    2.497801, 2.497806, 2.497801, 2.497802, 2.497797, 2.497799, 2.497788, 
    2.497794, 2.497777, 2.497772, 2.497755, 2.497745, 2.497734, 2.49773, 
    2.497728, 2.497728,
  2.498012, 2.498003, 2.498005, 2.497997, 2.498001, 2.497997, 2.49801, 
    2.498003, 2.498008, 2.498012, 2.497983, 2.497997, 2.497968, 2.497977, 
    2.497954, 2.497969, 2.497951, 2.497954, 2.497944, 2.497947, 2.497933, 
    2.497942, 2.497926, 2.497936, 2.497934, 2.497943, 2.497994, 2.497984, 
    2.497995, 2.497993, 2.497994, 2.498001, 2.498005, 2.498013, 2.498012, 
    2.498006, 2.497993, 2.497997, 2.497986, 2.497986, 2.497973, 2.497979, 
    2.497958, 2.497964, 2.497947, 2.497951, 2.497947, 2.497948, 2.497947, 
    2.497953, 2.497951, 2.497956, 2.497978, 2.497972, 2.497991, 2.498003, 
    2.49801, 2.498016, 2.498015, 2.498013, 2.498006, 2.497999, 2.497993, 
    2.49799, 2.497986, 2.497975, 2.49797, 2.497957, 2.497959, 2.497955, 
    2.497952, 2.497945, 2.497946, 2.497943, 2.497955, 2.497947, 2.49796, 
    2.497957, 2.497985, 2.497996, 2.498, 2.498004, 2.498014, 2.498008, 
    2.49801, 2.498004, 2.498, 2.498002, 2.49799, 2.497994, 2.497969, 2.49798, 
    2.497952, 2.497959, 2.49795, 2.497955, 2.497947, 2.497954, 2.497942, 
    2.49794, 2.497942, 2.497935, 2.497954, 2.497947, 2.498002, 2.498002, 
    2.498, 2.498007, 2.498007, 2.498013, 2.498008, 2.498005, 2.498, 2.497996, 
    2.497993, 2.497986, 2.497977, 2.497966, 2.497958, 2.497953, 2.497956, 
    2.497953, 2.497957, 2.497958, 2.497941, 2.497951, 2.497936, 2.497937, 
    2.497943, 2.497937, 2.498001, 2.498003, 2.49801, 2.498005, 2.498014, 
    2.498009, 2.498006, 2.497994, 2.497992, 2.497989, 2.497985, 2.497979, 
    2.497968, 2.497959, 2.497951, 2.497952, 2.497952, 2.49795, 2.497954, 
    2.497949, 2.497948, 2.497951, 2.497937, 2.497941, 2.497937, 2.497939, 
    2.498003, 2.497999, 2.498001, 2.497998, 2.498, 2.49799, 2.497987, 
    2.497973, 2.497979, 2.49797, 2.497978, 2.497977, 2.49797, 2.497977, 
    2.49796, 2.497972, 2.49795, 2.497962, 2.497949, 2.497951, 2.497947, 
    2.497944, 2.49794, 2.497932, 2.497934, 2.497927, 2.497995, 2.497991, 
    2.497991, 2.497987, 2.497984, 2.497977, 2.497966, 2.49797, 2.497962, 
    2.497961, 2.497972, 2.497965, 2.497988, 2.497984, 2.497987, 2.497994, 
    2.497969, 2.497982, 2.497958, 2.497965, 2.497945, 2.497955, 2.497935, 
    2.497926, 2.497918, 2.497909, 2.497988, 2.497991, 2.497986, 2.497979, 
    2.497973, 2.497965, 2.497964, 2.497962, 2.497958, 2.497955, 2.497962, 
    2.497954, 2.497983, 2.497968, 2.497992, 2.497985, 2.49798, 2.497982, 
    2.497971, 2.497968, 2.497957, 2.497962, 2.497928, 2.497943, 2.497901, 
    2.497913, 2.497992, 2.497988, 2.497976, 2.497982, 2.497964, 2.49796, 
    2.497956, 2.497952, 2.497951, 2.497949, 2.497953, 2.497949, 2.497965, 
    2.497957, 2.497977, 2.497972, 2.497974, 2.497977, 2.497969, 2.497962, 
    2.497962, 2.497959, 2.497952, 2.497964, 2.497926, 2.49795, 2.497984, 
    2.497977, 2.497976, 2.497979, 2.49796, 2.497967, 2.497949, 2.497954, 
    2.497946, 2.49795, 2.49795, 2.497955, 2.497959, 2.497967, 2.497973, 
    2.497979, 2.497977, 2.497972, 2.497961, 2.497951, 2.497953, 2.497946, 
    2.497965, 2.497957, 2.49796, 2.497952, 2.49797, 2.497955, 2.497974, 
    2.497972, 2.497967, 2.497957, 2.497954, 2.497952, 2.497953, 2.497961, 
    2.497962, 2.497967, 2.497969, 2.497973, 2.497976, 2.497973, 2.49797, 
    2.497961, 2.497953, 2.497944, 2.497942, 2.497931, 2.49794, 2.497926, 
    2.497938, 2.497918, 2.497954, 2.497938, 2.497967, 2.497964, 2.497958, 
    2.497945, 2.497952, 2.497944, 2.497962, 2.497971, 2.497974, 2.497978, 
    2.497974, 2.497974, 2.49797, 2.497971, 2.497961, 2.497966, 2.49795, 
    2.497944, 2.497928, 2.497918, 2.497907, 2.497903, 2.497901, 2.497901,
  2.498213, 2.498205, 2.498206, 2.4982, 2.498204, 2.498199, 2.498211, 
    2.498204, 2.498209, 2.498212, 2.498187, 2.498199, 2.498173, 2.498182, 
    2.498161, 2.498175, 2.498158, 2.498162, 2.498152, 2.498155, 2.498143, 
    2.498151, 2.498137, 2.498145, 2.498143, 2.498151, 2.498197, 2.498188, 
    2.498197, 2.498196, 2.498197, 2.498203, 2.498207, 2.498214, 2.498212, 
    2.498207, 2.498196, 2.498199, 2.498189, 2.49819, 2.498178, 2.498184, 
    2.498165, 2.49817, 2.498155, 2.498159, 2.498155, 2.498156, 2.498155, 
    2.498161, 2.498158, 2.498163, 2.498183, 2.498177, 2.498194, 2.498204, 
    2.498211, 2.498216, 2.498215, 2.498214, 2.498207, 2.498201, 2.498196, 
    2.498193, 2.49819, 2.49818, 2.498175, 2.498164, 2.498166, 2.498162, 
    2.498159, 2.498153, 2.498154, 2.498152, 2.498163, 2.498155, 2.498167, 
    2.498164, 2.498189, 2.498199, 2.498203, 2.498206, 2.498215, 2.498209, 
    2.498211, 2.498205, 2.498202, 2.498204, 2.498193, 2.498197, 2.498175, 
    2.498184, 2.498159, 2.498165, 2.498158, 2.498162, 2.498155, 2.498161, 
    2.498151, 2.498149, 2.49815, 2.498144, 2.498161, 2.498155, 2.498204, 
    2.498204, 2.498202, 2.498208, 2.498208, 2.498214, 2.498209, 2.498207, 
    2.498202, 2.498199, 2.498196, 2.498189, 2.498182, 2.498172, 2.498165, 
    2.49816, 2.498163, 2.498161, 2.498163, 2.498165, 2.49815, 2.498158, 
    2.498145, 2.498146, 2.498152, 2.498146, 2.498203, 2.498205, 2.498211, 
    2.498206, 2.498214, 2.49821, 2.498207, 2.498197, 2.498195, 2.498193, 
    2.498188, 2.498183, 2.498174, 2.498166, 2.498159, 2.498159, 2.498159, 
    2.498158, 2.498162, 2.498157, 2.498156, 2.498158, 2.498146, 2.49815, 
    2.498146, 2.498148, 2.498204, 2.498202, 2.498203, 2.4982, 2.498202, 
    2.498194, 2.498191, 2.498178, 2.498183, 2.498175, 2.498183, 2.498181, 
    2.498175, 2.498182, 2.498167, 2.498177, 2.498158, 2.498168, 2.498157, 
    2.498159, 2.498155, 2.498152, 2.498149, 2.498142, 2.498143, 2.498137, 
    2.498198, 2.498194, 2.498194, 2.49819, 2.498188, 2.498182, 2.498172, 
    2.498176, 2.498169, 2.498168, 2.498178, 2.498171, 2.498191, 2.498188, 
    2.49819, 2.498197, 2.498175, 2.498186, 2.498165, 2.498171, 2.498153, 
    2.498162, 2.498144, 2.498136, 2.498129, 2.498121, 2.498192, 2.498194, 
    2.49819, 2.498184, 2.498178, 2.498171, 2.49817, 2.498168, 2.498165, 
    2.498162, 2.498168, 2.498161, 2.498188, 2.498174, 2.498195, 2.498189, 
    2.498184, 2.498186, 2.498176, 2.498173, 2.498164, 2.498169, 2.498138, 
    2.498152, 2.498114, 2.498125, 2.498195, 2.498192, 2.49818, 2.498186, 
    2.49817, 2.498166, 2.498163, 2.498159, 2.498159, 2.498157, 2.49816, 
    2.498157, 2.498171, 2.498164, 2.498182, 2.498178, 2.498179, 2.498182, 
    2.498175, 2.498168, 2.498168, 2.498166, 2.498159, 2.49817, 2.498137, 
    2.498157, 2.498188, 2.498182, 2.498181, 2.498183, 2.498167, 2.498173, 
    2.498157, 2.498161, 2.498154, 2.498157, 2.498158, 2.498163, 2.498165, 
    2.498173, 2.498178, 2.498183, 2.498182, 2.498177, 2.498168, 2.498159, 
    2.498161, 2.498154, 2.498171, 2.498164, 2.498167, 2.49816, 2.498176, 
    2.498162, 2.498179, 2.498178, 2.498173, 2.498164, 2.498162, 2.498159, 
    2.498161, 2.498167, 2.498168, 2.498173, 2.498174, 2.498178, 2.498181, 
    2.498178, 2.498175, 2.498167, 2.49816, 2.498152, 2.49815, 2.498141, 
    2.498149, 2.498137, 2.498147, 2.498129, 2.498161, 2.498147, 2.498173, 
    2.49817, 2.498165, 2.498154, 2.49816, 2.498152, 2.498168, 2.498177, 
    2.498179, 2.498183, 2.498179, 2.498179, 2.498175, 2.498177, 2.498167, 
    2.498172, 2.498158, 2.498153, 2.498138, 2.498129, 2.49812, 2.498116, 
    2.498114, 2.498114,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  6.140732e-08, 6.167728e-08, 6.16248e-08, 6.184255e-08, 6.172176e-08, 
    6.186434e-08, 6.146205e-08, 6.168801e-08, 6.154376e-08, 6.143162e-08, 
    6.226513e-08, 6.185226e-08, 6.269395e-08, 6.243065e-08, 6.309206e-08, 
    6.265298e-08, 6.318059e-08, 6.307938e-08, 6.338397e-08, 6.329671e-08, 
    6.368631e-08, 6.342425e-08, 6.388827e-08, 6.362372e-08, 6.366511e-08, 
    6.34156e-08, 6.193535e-08, 6.221374e-08, 6.191885e-08, 6.195855e-08, 
    6.194074e-08, 6.172426e-08, 6.161517e-08, 6.138668e-08, 6.142816e-08, 
    6.159598e-08, 6.19764e-08, 6.184726e-08, 6.217271e-08, 6.216536e-08, 
    6.252768e-08, 6.236432e-08, 6.297329e-08, 6.280021e-08, 6.330036e-08, 
    6.317457e-08, 6.329445e-08, 6.32581e-08, 6.329492e-08, 6.311045e-08, 
    6.318949e-08, 6.302716e-08, 6.239492e-08, 6.258073e-08, 6.202654e-08, 
    6.169331e-08, 6.147196e-08, 6.131489e-08, 6.13371e-08, 6.137943e-08, 
    6.159696e-08, 6.180147e-08, 6.195733e-08, 6.206158e-08, 6.21643e-08, 
    6.247526e-08, 6.263982e-08, 6.300829e-08, 6.294179e-08, 6.305444e-08, 
    6.316206e-08, 6.334275e-08, 6.331301e-08, 6.339262e-08, 6.305147e-08, 
    6.32782e-08, 6.290391e-08, 6.300628e-08, 6.219226e-08, 6.18821e-08, 
    6.175029e-08, 6.163489e-08, 6.135417e-08, 6.154804e-08, 6.147161e-08, 
    6.165342e-08, 6.176894e-08, 6.17118e-08, 6.206443e-08, 6.192735e-08, 
    6.264957e-08, 6.233849e-08, 6.314951e-08, 6.295544e-08, 6.319603e-08, 
    6.307326e-08, 6.328361e-08, 6.30943e-08, 6.342224e-08, 6.349365e-08, 
    6.344485e-08, 6.363231e-08, 6.30838e-08, 6.329445e-08, 6.17102e-08, 
    6.171953e-08, 6.176293e-08, 6.157211e-08, 6.156043e-08, 6.138554e-08, 
    6.154116e-08, 6.160742e-08, 6.177564e-08, 6.187514e-08, 6.196972e-08, 
    6.217768e-08, 6.240995e-08, 6.273471e-08, 6.296802e-08, 6.312441e-08, 
    6.302851e-08, 6.311318e-08, 6.301853e-08, 6.297417e-08, 6.34669e-08, 
    6.319023e-08, 6.360534e-08, 6.358237e-08, 6.339451e-08, 6.358496e-08, 
    6.172607e-08, 6.167244e-08, 6.148626e-08, 6.163197e-08, 6.13665e-08, 
    6.15151e-08, 6.160054e-08, 6.193022e-08, 6.200263e-08, 6.20698e-08, 
    6.220245e-08, 6.237268e-08, 6.267131e-08, 6.293114e-08, 6.316832e-08, 
    6.315094e-08, 6.315706e-08, 6.321005e-08, 6.30788e-08, 6.32316e-08, 
    6.325725e-08, 6.319019e-08, 6.357929e-08, 6.346813e-08, 6.358189e-08, 
    6.35095e-08, 6.168987e-08, 6.178011e-08, 6.173135e-08, 6.182303e-08, 
    6.175844e-08, 6.204566e-08, 6.213178e-08, 6.25347e-08, 6.236933e-08, 
    6.263252e-08, 6.239606e-08, 6.243796e-08, 6.264111e-08, 6.240884e-08, 
    6.291682e-08, 6.257244e-08, 6.321211e-08, 6.286822e-08, 6.323366e-08, 
    6.316729e-08, 6.327717e-08, 6.337557e-08, 6.349937e-08, 6.37278e-08, 
    6.36749e-08, 6.386593e-08, 6.191462e-08, 6.203165e-08, 6.202134e-08, 
    6.214382e-08, 6.22344e-08, 6.243071e-08, 6.274558e-08, 6.262717e-08, 
    6.284454e-08, 6.288818e-08, 6.255794e-08, 6.276071e-08, 6.210998e-08, 
    6.221512e-08, 6.215252e-08, 6.192385e-08, 6.265446e-08, 6.227952e-08, 
    6.297187e-08, 6.276876e-08, 6.336155e-08, 6.306675e-08, 6.364579e-08, 
    6.389333e-08, 6.412628e-08, 6.439855e-08, 6.209552e-08, 6.2016e-08, 
    6.215839e-08, 6.235538e-08, 6.253816e-08, 6.278115e-08, 6.280601e-08, 
    6.285153e-08, 6.296944e-08, 6.306858e-08, 6.286593e-08, 6.309343e-08, 
    6.223951e-08, 6.268701e-08, 6.198594e-08, 6.219706e-08, 6.234377e-08, 
    6.22794e-08, 6.261364e-08, 6.269241e-08, 6.301254e-08, 6.284705e-08, 
    6.383225e-08, 6.339637e-08, 6.460584e-08, 6.426785e-08, 6.198822e-08, 
    6.209525e-08, 6.246775e-08, 6.229051e-08, 6.279737e-08, 6.292213e-08, 
    6.302354e-08, 6.315319e-08, 6.316719e-08, 6.3244e-08, 6.311813e-08, 
    6.323903e-08, 6.278167e-08, 6.298605e-08, 6.242517e-08, 6.256169e-08, 
    6.249888e-08, 6.242999e-08, 6.264261e-08, 6.286912e-08, 6.287395e-08, 
    6.294658e-08, 6.315128e-08, 6.279942e-08, 6.388851e-08, 6.321594e-08, 
    6.221196e-08, 6.241812e-08, 6.244756e-08, 6.23677e-08, 6.290962e-08, 
    6.271326e-08, 6.324213e-08, 6.309919e-08, 6.333339e-08, 6.321702e-08, 
    6.319989e-08, 6.305042e-08, 6.295737e-08, 6.272227e-08, 6.253098e-08, 
    6.237928e-08, 6.241455e-08, 6.258119e-08, 6.288298e-08, 6.316846e-08, 
    6.310592e-08, 6.331559e-08, 6.276061e-08, 6.299333e-08, 6.290339e-08, 
    6.313791e-08, 6.262403e-08, 6.306166e-08, 6.251217e-08, 6.256035e-08, 
    6.270937e-08, 6.300913e-08, 6.307543e-08, 6.314624e-08, 6.310254e-08, 
    6.289063e-08, 6.285591e-08, 6.270574e-08, 6.266428e-08, 6.254986e-08, 
    6.245513e-08, 6.254168e-08, 6.263258e-08, 6.289072e-08, 6.312335e-08, 
    6.337698e-08, 6.343905e-08, 6.37354e-08, 6.349416e-08, 6.389227e-08, 
    6.355383e-08, 6.413967e-08, 6.3087e-08, 6.354385e-08, 6.271615e-08, 
    6.280531e-08, 6.296661e-08, 6.333652e-08, 6.313681e-08, 6.337036e-08, 
    6.285455e-08, 6.258694e-08, 6.251769e-08, 6.23885e-08, 6.252064e-08, 
    6.25099e-08, 6.263634e-08, 6.25957e-08, 6.289929e-08, 6.273622e-08, 
    6.319947e-08, 6.336852e-08, 6.384592e-08, 6.413858e-08, 6.443647e-08, 
    6.456799e-08, 6.460802e-08, 6.462475e-08 ;

 SOIL1_HR_S3 =
  7.287159e-10, 7.319208e-10, 7.312977e-10, 7.338827e-10, 7.324487e-10, 
    7.341414e-10, 7.293656e-10, 7.320481e-10, 7.303356e-10, 7.290044e-10, 
    7.388995e-10, 7.33998e-10, 7.439904e-10, 7.408645e-10, 7.487168e-10, 
    7.43504e-10, 7.497678e-10, 7.485663e-10, 7.521824e-10, 7.511464e-10, 
    7.557719e-10, 7.526605e-10, 7.581696e-10, 7.550289e-10, 7.555202e-10, 
    7.525579e-10, 7.349844e-10, 7.382893e-10, 7.347886e-10, 7.352599e-10, 
    7.350484e-10, 7.324784e-10, 7.311834e-10, 7.284708e-10, 7.289633e-10, 
    7.309555e-10, 7.354717e-10, 7.339386e-10, 7.378023e-10, 7.37715e-10, 
    7.420164e-10, 7.400771e-10, 7.473067e-10, 7.452519e-10, 7.511897e-10, 
    7.496964e-10, 7.511196e-10, 7.50688e-10, 7.511252e-10, 7.489351e-10, 
    7.498734e-10, 7.479463e-10, 7.404403e-10, 7.426463e-10, 7.36067e-10, 
    7.32111e-10, 7.294833e-10, 7.276186e-10, 7.278823e-10, 7.283848e-10, 
    7.309672e-10, 7.333951e-10, 7.352453e-10, 7.36483e-10, 7.377025e-10, 
    7.413941e-10, 7.433477e-10, 7.477223e-10, 7.469327e-10, 7.482702e-10, 
    7.495478e-10, 7.51693e-10, 7.513399e-10, 7.52285e-10, 7.482348e-10, 
    7.509267e-10, 7.464829e-10, 7.476983e-10, 7.380344e-10, 7.343522e-10, 
    7.327874e-10, 7.314175e-10, 7.280849e-10, 7.303864e-10, 7.294791e-10, 
    7.316374e-10, 7.330089e-10, 7.323305e-10, 7.365168e-10, 7.348893e-10, 
    7.434635e-10, 7.397703e-10, 7.493988e-10, 7.470947e-10, 7.49951e-10, 
    7.484935e-10, 7.509909e-10, 7.487433e-10, 7.526367e-10, 7.534846e-10, 
    7.529052e-10, 7.551307e-10, 7.486187e-10, 7.511196e-10, 7.323115e-10, 
    7.324222e-10, 7.329375e-10, 7.306721e-10, 7.305335e-10, 7.284573e-10, 
    7.303047e-10, 7.310914e-10, 7.330884e-10, 7.342696e-10, 7.353925e-10, 
    7.378613e-10, 7.406187e-10, 7.444742e-10, 7.472441e-10, 7.491008e-10, 
    7.479623e-10, 7.489674e-10, 7.478438e-10, 7.473171e-10, 7.531669e-10, 
    7.498822e-10, 7.548106e-10, 7.545379e-10, 7.523075e-10, 7.545686e-10, 
    7.324999e-10, 7.318632e-10, 7.296531e-10, 7.313827e-10, 7.282313e-10, 
    7.299953e-10, 7.310097e-10, 7.349234e-10, 7.357832e-10, 7.365806e-10, 
    7.381553e-10, 7.401763e-10, 7.437216e-10, 7.468062e-10, 7.496221e-10, 
    7.494158e-10, 7.494885e-10, 7.501175e-10, 7.485593e-10, 7.503734e-10, 
    7.506779e-10, 7.498818e-10, 7.545014e-10, 7.531816e-10, 7.545321e-10, 
    7.536727e-10, 7.320702e-10, 7.331414e-10, 7.325626e-10, 7.33651e-10, 
    7.328842e-10, 7.36294e-10, 7.373163e-10, 7.420998e-10, 7.401366e-10, 
    7.43261e-10, 7.404539e-10, 7.409513e-10, 7.43363e-10, 7.406056e-10, 
    7.466363e-10, 7.425477e-10, 7.50142e-10, 7.460594e-10, 7.503979e-10, 
    7.4961e-10, 7.509144e-10, 7.520827e-10, 7.535525e-10, 7.562645e-10, 
    7.556365e-10, 7.579045e-10, 7.347383e-10, 7.361277e-10, 7.360053e-10, 
    7.374593e-10, 7.385346e-10, 7.408652e-10, 7.446033e-10, 7.431976e-10, 
    7.457782e-10, 7.462962e-10, 7.423757e-10, 7.447829e-10, 7.370575e-10, 
    7.383057e-10, 7.375625e-10, 7.348479e-10, 7.435216e-10, 7.390703e-10, 
    7.472899e-10, 7.448785e-10, 7.519161e-10, 7.484162e-10, 7.552908e-10, 
    7.582298e-10, 7.609955e-10, 7.642281e-10, 7.368859e-10, 7.359418e-10, 
    7.376322e-10, 7.39971e-10, 7.421408e-10, 7.450256e-10, 7.453207e-10, 
    7.458612e-10, 7.47261e-10, 7.48438e-10, 7.460321e-10, 7.48733e-10, 
    7.385954e-10, 7.43908e-10, 7.35585e-10, 7.380913e-10, 7.398331e-10, 
    7.390689e-10, 7.430369e-10, 7.439722e-10, 7.477726e-10, 7.45808e-10, 
    7.575045e-10, 7.523296e-10, 7.666892e-10, 7.626763e-10, 7.35612e-10, 
    7.368826e-10, 7.41305e-10, 7.392008e-10, 7.452181e-10, 7.466993e-10, 
    7.479033e-10, 7.494426e-10, 7.496087e-10, 7.505206e-10, 7.490262e-10, 
    7.504616e-10, 7.450317e-10, 7.474582e-10, 7.407994e-10, 7.424201e-10, 
    7.416745e-10, 7.408567e-10, 7.433807e-10, 7.4607e-10, 7.461273e-10, 
    7.469896e-10, 7.494199e-10, 7.452425e-10, 7.581726e-10, 7.501875e-10, 
    7.382682e-10, 7.407158e-10, 7.410652e-10, 7.401171e-10, 7.465508e-10, 
    7.442197e-10, 7.504984e-10, 7.488015e-10, 7.515819e-10, 7.502002e-10, 
    7.49997e-10, 7.482224e-10, 7.471177e-10, 7.443265e-10, 7.420555e-10, 
    7.402546e-10, 7.406734e-10, 7.426517e-10, 7.462345e-10, 7.496238e-10, 
    7.488813e-10, 7.513706e-10, 7.447818e-10, 7.475446e-10, 7.464768e-10, 
    7.492611e-10, 7.431603e-10, 7.483558e-10, 7.418323e-10, 7.424042e-10, 
    7.441734e-10, 7.477321e-10, 7.485193e-10, 7.4936e-10, 7.488412e-10, 
    7.463254e-10, 7.459132e-10, 7.441304e-10, 7.436382e-10, 7.422797e-10, 
    7.411551e-10, 7.421826e-10, 7.432618e-10, 7.463264e-10, 7.490882e-10, 
    7.520994e-10, 7.528362e-10, 7.563548e-10, 7.534907e-10, 7.582171e-10, 
    7.54199e-10, 7.611545e-10, 7.486567e-10, 7.540806e-10, 7.442538e-10, 
    7.453125e-10, 7.472273e-10, 7.51619e-10, 7.49248e-10, 7.520209e-10, 
    7.45897e-10, 7.427199e-10, 7.418978e-10, 7.403641e-10, 7.419328e-10, 
    7.418053e-10, 7.433064e-10, 7.42824e-10, 7.464281e-10, 7.444922e-10, 
    7.499919e-10, 7.51999e-10, 7.576668e-10, 7.611415e-10, 7.646783e-10, 
    7.662398e-10, 7.667151e-10, 7.669138e-10 ;

 SOIL2C =
  5.784045, 5.784051, 5.78405, 5.784055, 5.784052, 5.784055, 5.784046, 
    5.784051, 5.784048, 5.784045, 5.784065, 5.784055, 5.784075, 5.784069, 
    5.784084, 5.784074, 5.784086, 5.784084, 5.784091, 5.784089, 5.784098, 
    5.784092, 5.784103, 5.784097, 5.784098, 5.784092, 5.784057, 5.784063, 
    5.784057, 5.784058, 5.784057, 5.784052, 5.78405, 5.784044, 5.784045, 
    5.784049, 5.784058, 5.784055, 5.784062, 5.784062, 5.784071, 5.784067, 
    5.784081, 5.784077, 5.784089, 5.784086, 5.784089, 5.784088, 5.784089, 
    5.784085, 5.784086, 5.784082, 5.784068, 5.784072, 5.784059, 5.784051, 
    5.784046, 5.784042, 5.784043, 5.784044, 5.784049, 5.784054, 5.784058, 
    5.78406, 5.784062, 5.78407, 5.784073, 5.784082, 5.784081, 5.784083, 
    5.784086, 5.78409, 5.784089, 5.784091, 5.784083, 5.784089, 5.78408, 
    5.784082, 5.784063, 5.784056, 5.784053, 5.78405, 5.784043, 5.784048, 
    5.784046, 5.78405, 5.784053, 5.784052, 5.78406, 5.784057, 5.784074, 
    5.784067, 5.784085, 5.784081, 5.784087, 5.784084, 5.784089, 5.784084, 
    5.784092, 5.784093, 5.784092, 5.784097, 5.784084, 5.784089, 5.784052, 
    5.784052, 5.784053, 5.784049, 5.784048, 5.784044, 5.784048, 5.78405, 
    5.784053, 5.784056, 5.784058, 5.784063, 5.784068, 5.784076, 5.784081, 
    5.784085, 5.784082, 5.784085, 5.784082, 5.784081, 5.784093, 5.784086, 
    5.784096, 5.784096, 5.784091, 5.784096, 5.784052, 5.784051, 5.784047, 
    5.78405, 5.784044, 5.784047, 5.784049, 5.784057, 5.784059, 5.78406, 
    5.784063, 5.784067, 5.784074, 5.784081, 5.784086, 5.784086, 5.784086, 
    5.784087, 5.784084, 5.784087, 5.784088, 5.784086, 5.784096, 5.784093, 
    5.784096, 5.784094, 5.784051, 5.784053, 5.784052, 5.784054, 5.784053, 
    5.78406, 5.784061, 5.784071, 5.784067, 5.784073, 5.784068, 5.784069, 
    5.784073, 5.784068, 5.78408, 5.784072, 5.784087, 5.784079, 5.784088, 
    5.784086, 5.784089, 5.784091, 5.784094, 5.784099, 5.784098, 5.784102, 
    5.784057, 5.784059, 5.784059, 5.784062, 5.784064, 5.784069, 5.784076, 
    5.784073, 5.784078, 5.78408, 5.784071, 5.784076, 5.784061, 5.784064, 
    5.784062, 5.784057, 5.784074, 5.784065, 5.784081, 5.784077, 5.784091, 
    5.784083, 5.784097, 5.784103, 5.784108, 5.784115, 5.784061, 5.784059, 
    5.784062, 5.784067, 5.784071, 5.784077, 5.784078, 5.784079, 5.784081, 
    5.784083, 5.784079, 5.784084, 5.784064, 5.784075, 5.784058, 5.784063, 
    5.784067, 5.784065, 5.784073, 5.784075, 5.784082, 5.784079, 5.784101, 
    5.784091, 5.78412, 5.784111, 5.784058, 5.784061, 5.78407, 5.784065, 
    5.784077, 5.78408, 5.784082, 5.784086, 5.784086, 5.784088, 5.784085, 
    5.784088, 5.784077, 5.784081, 5.784069, 5.784072, 5.78407, 5.784069, 
    5.784074, 5.784079, 5.784079, 5.784081, 5.784086, 5.784077, 5.784103, 
    5.784087, 5.784063, 5.784068, 5.784069, 5.784067, 5.78408, 5.784075, 
    5.784088, 5.784084, 5.78409, 5.784087, 5.784087, 5.784083, 5.784081, 
    5.784075, 5.784071, 5.784068, 5.784068, 5.784072, 5.784079, 5.784086, 
    5.784084, 5.78409, 5.784076, 5.784082, 5.78408, 5.784085, 5.784073, 
    5.784083, 5.78407, 5.784071, 5.784075, 5.784082, 5.784084, 5.784085, 
    5.784084, 5.78408, 5.784079, 5.784075, 5.784074, 5.784071, 5.784069, 
    5.784071, 5.784073, 5.78408, 5.784085, 5.784091, 5.784092, 5.784099, 
    5.784093, 5.784103, 5.784095, 5.784109, 5.784084, 5.784095, 5.784075, 
    5.784078, 5.784081, 5.78409, 5.784085, 5.784091, 5.784079, 5.784072, 
    5.78407, 5.784068, 5.784071, 5.78407, 5.784073, 5.784072, 5.78408, 
    5.784076, 5.784087, 5.784091, 5.784102, 5.784109, 5.784116, 5.784119, 
    5.78412, 5.78412 ;

 SOIL2C_TO_SOIL1C =
  1.086416e-09, 1.091196e-09, 1.090267e-09, 1.094122e-09, 1.091984e-09, 
    1.094508e-09, 1.087385e-09, 1.091386e-09, 1.088832e-09, 1.086846e-09, 
    1.101604e-09, 1.094294e-09, 1.109197e-09, 1.104535e-09, 1.116245e-09, 
    1.108471e-09, 1.117813e-09, 1.116021e-09, 1.121414e-09, 1.119869e-09, 
    1.126767e-09, 1.122127e-09, 1.130342e-09, 1.125659e-09, 1.126391e-09, 
    1.121974e-09, 1.095765e-09, 1.100694e-09, 1.095473e-09, 1.096176e-09, 
    1.095861e-09, 1.092028e-09, 1.090096e-09, 1.086051e-09, 1.086785e-09, 
    1.089756e-09, 1.096492e-09, 1.094206e-09, 1.099968e-09, 1.099838e-09, 
    1.106253e-09, 1.10336e-09, 1.114142e-09, 1.111078e-09, 1.119933e-09, 
    1.117706e-09, 1.119829e-09, 1.119185e-09, 1.119837e-09, 1.116571e-09, 
    1.11797e-09, 1.115096e-09, 1.103902e-09, 1.107192e-09, 1.09738e-09, 
    1.09148e-09, 1.087561e-09, 1.08478e-09, 1.085173e-09, 1.085922e-09, 
    1.089774e-09, 1.093395e-09, 1.096154e-09, 1.098e-09, 1.099819e-09, 
    1.105324e-09, 1.108238e-09, 1.114762e-09, 1.113585e-09, 1.115579e-09, 
    1.117485e-09, 1.120684e-09, 1.120157e-09, 1.121567e-09, 1.115526e-09, 
    1.119541e-09, 1.112914e-09, 1.114726e-09, 1.100314e-09, 1.094822e-09, 
    1.092489e-09, 1.090445e-09, 1.085475e-09, 1.088908e-09, 1.087554e-09, 
    1.090773e-09, 1.092819e-09, 1.091807e-09, 1.098051e-09, 1.095623e-09, 
    1.108411e-09, 1.102903e-09, 1.117262e-09, 1.113826e-09, 1.118086e-09, 
    1.115912e-09, 1.119637e-09, 1.116285e-09, 1.122091e-09, 1.123356e-09, 
    1.122492e-09, 1.125811e-09, 1.116099e-09, 1.119829e-09, 1.091779e-09, 
    1.091944e-09, 1.092712e-09, 1.089334e-09, 1.089127e-09, 1.086031e-09, 
    1.088786e-09, 1.089959e-09, 1.092937e-09, 1.094699e-09, 1.096374e-09, 
    1.100056e-09, 1.104168e-09, 1.109918e-09, 1.114049e-09, 1.116818e-09, 
    1.11512e-09, 1.116619e-09, 1.114943e-09, 1.114158e-09, 1.122882e-09, 
    1.117983e-09, 1.125333e-09, 1.124926e-09, 1.1216e-09, 1.124972e-09, 
    1.09206e-09, 1.09111e-09, 1.087814e-09, 1.090394e-09, 1.085693e-09, 
    1.088324e-09, 1.089837e-09, 1.095674e-09, 1.096957e-09, 1.098146e-09, 
    1.100494e-09, 1.103508e-09, 1.108796e-09, 1.113396e-09, 1.117595e-09, 
    1.117288e-09, 1.117396e-09, 1.118334e-09, 1.11601e-09, 1.118716e-09, 
    1.11917e-09, 1.117983e-09, 1.124872e-09, 1.122904e-09, 1.124918e-09, 
    1.123636e-09, 1.091419e-09, 1.093016e-09, 1.092153e-09, 1.093777e-09, 
    1.092633e-09, 1.097718e-09, 1.099243e-09, 1.106377e-09, 1.103449e-09, 
    1.108109e-09, 1.103922e-09, 1.104664e-09, 1.108261e-09, 1.104148e-09, 
    1.113142e-09, 1.107045e-09, 1.118371e-09, 1.112282e-09, 1.118752e-09, 
    1.117577e-09, 1.119523e-09, 1.121265e-09, 1.123457e-09, 1.127501e-09, 
    1.126565e-09, 1.129947e-09, 1.095398e-09, 1.09747e-09, 1.097288e-09, 
    1.099456e-09, 1.10106e-09, 1.104536e-09, 1.110111e-09, 1.108014e-09, 
    1.111863e-09, 1.112635e-09, 1.106788e-09, 1.110378e-09, 1.098857e-09, 
    1.100719e-09, 1.09961e-09, 1.095562e-09, 1.108497e-09, 1.101859e-09, 
    1.114117e-09, 1.110521e-09, 1.121017e-09, 1.115797e-09, 1.126049e-09, 
    1.130432e-09, 1.134557e-09, 1.139377e-09, 1.098601e-09, 1.097193e-09, 
    1.099714e-09, 1.103202e-09, 1.106438e-09, 1.11074e-09, 1.11118e-09, 
    1.111987e-09, 1.114074e-09, 1.115829e-09, 1.112241e-09, 1.11627e-09, 
    1.101151e-09, 1.109074e-09, 1.096661e-09, 1.100399e-09, 1.102996e-09, 
    1.101857e-09, 1.107775e-09, 1.109169e-09, 1.114837e-09, 1.111907e-09, 
    1.129351e-09, 1.121633e-09, 1.143048e-09, 1.137063e-09, 1.096701e-09, 
    1.098596e-09, 1.105191e-09, 1.102053e-09, 1.111027e-09, 1.113236e-09, 
    1.115032e-09, 1.117328e-09, 1.117575e-09, 1.118935e-09, 1.116707e-09, 
    1.118847e-09, 1.110749e-09, 1.114368e-09, 1.104438e-09, 1.106855e-09, 
    1.105743e-09, 1.104523e-09, 1.108287e-09, 1.112298e-09, 1.112383e-09, 
    1.113669e-09, 1.117294e-09, 1.111064e-09, 1.130347e-09, 1.118438e-09, 
    1.100663e-09, 1.104313e-09, 1.104834e-09, 1.10342e-09, 1.113015e-09, 
    1.109538e-09, 1.118902e-09, 1.116372e-09, 1.120518e-09, 1.118458e-09, 
    1.118154e-09, 1.115508e-09, 1.11386e-09, 1.109698e-09, 1.106311e-09, 
    1.103625e-09, 1.10425e-09, 1.1072e-09, 1.112543e-09, 1.117598e-09, 
    1.116491e-09, 1.120203e-09, 1.110377e-09, 1.114497e-09, 1.112905e-09, 
    1.117057e-09, 1.107959e-09, 1.115707e-09, 1.105978e-09, 1.106831e-09, 
    1.109469e-09, 1.114777e-09, 1.115951e-09, 1.117204e-09, 1.116431e-09, 
    1.112679e-09, 1.112064e-09, 1.109405e-09, 1.108671e-09, 1.106645e-09, 
    1.104968e-09, 1.1065e-09, 1.10811e-09, 1.11268e-09, 1.116799e-09, 
    1.12129e-09, 1.122389e-09, 1.127636e-09, 1.123365e-09, 1.130413e-09, 
    1.124421e-09, 1.134794e-09, 1.116156e-09, 1.124244e-09, 1.109589e-09, 
    1.111168e-09, 1.114024e-09, 1.120574e-09, 1.117037e-09, 1.121173e-09, 
    1.11204e-09, 1.107302e-09, 1.106076e-09, 1.103788e-09, 1.106128e-09, 
    1.105938e-09, 1.108176e-09, 1.107457e-09, 1.112832e-09, 1.109945e-09, 
    1.118147e-09, 1.12114e-09, 1.129593e-09, 1.134774e-09, 1.140049e-09, 
    1.142378e-09, 1.143086e-09, 1.143382e-09 ;

 SOIL2C_TO_SOIL3C =
  7.760115e-11, 7.794258e-11, 7.78762e-11, 7.815158e-11, 7.799882e-11, 
    7.817914e-11, 7.767037e-11, 7.795613e-11, 7.77737e-11, 7.763189e-11, 
    7.8686e-11, 7.816386e-11, 7.922832e-11, 7.889533e-11, 7.97318e-11, 
    7.917651e-11, 7.984376e-11, 7.971577e-11, 8.010097e-11, 7.999062e-11, 
    8.048335e-11, 8.015191e-11, 8.073875e-11, 8.040419e-11, 8.045653e-11, 
    8.014098e-11, 7.826893e-11, 7.862101e-11, 7.824807e-11, 7.829828e-11, 
    7.827575e-11, 7.800198e-11, 7.786402e-11, 7.757506e-11, 7.762752e-11, 
    7.783975e-11, 7.832086e-11, 7.815754e-11, 7.856912e-11, 7.855983e-11, 
    7.901805e-11, 7.881144e-11, 7.958159e-11, 7.93627e-11, 7.999523e-11, 
    7.983616e-11, 7.998776e-11, 7.994178e-11, 7.998836e-11, 7.975506e-11, 
    7.985502e-11, 7.964972e-11, 7.885014e-11, 7.908514e-11, 7.838426e-11, 
    7.796284e-11, 7.768291e-11, 7.748427e-11, 7.751235e-11, 7.756588e-11, 
    7.784098e-11, 7.809963e-11, 7.829673e-11, 7.842858e-11, 7.855849e-11, 
    7.895174e-11, 7.915986e-11, 7.962586e-11, 7.954176e-11, 7.968423e-11, 
    7.982033e-11, 8.004884e-11, 8.001123e-11, 8.011191e-11, 7.968046e-11, 
    7.996721e-11, 7.949384e-11, 7.962331e-11, 7.859385e-11, 7.820159e-11, 
    7.80349e-11, 7.788896e-11, 7.753394e-11, 7.777912e-11, 7.768246e-11, 
    7.791238e-11, 7.805849e-11, 7.798623e-11, 7.843218e-11, 7.825881e-11, 
    7.91722e-11, 7.877878e-11, 7.980445e-11, 7.955901e-11, 7.986328e-11, 
    7.970802e-11, 7.997406e-11, 7.973463e-11, 8.014937e-11, 8.023969e-11, 
    8.017798e-11, 8.041504e-11, 7.972135e-11, 7.998776e-11, 7.79842e-11, 
    7.799599e-11, 7.805089e-11, 7.780956e-11, 7.779479e-11, 7.757362e-11, 
    7.777042e-11, 7.785422e-11, 7.806696e-11, 7.819279e-11, 7.831241e-11, 
    7.857542e-11, 7.886914e-11, 7.927986e-11, 7.957492e-11, 7.977272e-11, 
    7.965143e-11, 7.975851e-11, 7.963881e-11, 7.95827e-11, 8.020585e-11, 
    7.985595e-11, 8.038094e-11, 8.035189e-11, 8.01143e-11, 8.035516e-11, 
    7.800426e-11, 7.793645e-11, 7.770099e-11, 7.788525e-11, 7.754953e-11, 
    7.773746e-11, 7.784552e-11, 7.826245e-11, 7.835404e-11, 7.843898e-11, 
    7.860673e-11, 7.882202e-11, 7.919969e-11, 7.952829e-11, 7.982825e-11, 
    7.980627e-11, 7.9814e-11, 7.988102e-11, 7.971503e-11, 7.990827e-11, 
    7.994071e-11, 7.985591e-11, 8.0348e-11, 8.020741e-11, 8.035127e-11, 
    8.025973e-11, 7.795849e-11, 7.80726e-11, 7.801094e-11, 7.812689e-11, 
    7.804521e-11, 7.840845e-11, 7.851735e-11, 7.902692e-11, 7.881779e-11, 
    7.915062e-11, 7.885159e-11, 7.890458e-11, 7.91615e-11, 7.886775e-11, 
    7.951018e-11, 7.907464e-11, 7.988363e-11, 7.944872e-11, 7.991088e-11, 
    7.982695e-11, 7.99659e-11, 8.009036e-11, 8.024692e-11, 8.053581e-11, 
    8.046892e-11, 8.071051e-11, 7.824272e-11, 7.839073e-11, 7.837769e-11, 
    7.853258e-11, 7.864714e-11, 7.889541e-11, 7.929361e-11, 7.914387e-11, 
    7.941877e-11, 7.947396e-11, 7.905632e-11, 7.931275e-11, 7.848978e-11, 
    7.862275e-11, 7.854358e-11, 7.82544e-11, 7.917839e-11, 7.87042e-11, 
    7.95798e-11, 7.932293e-11, 8.007262e-11, 7.969979e-11, 8.043209e-11, 
    8.074516e-11, 8.103977e-11, 8.138411e-11, 7.847151e-11, 7.837093e-11, 
    7.8551e-11, 7.880015e-11, 7.903129e-11, 7.93386e-11, 7.937003e-11, 
    7.942761e-11, 7.957672e-11, 7.970211e-11, 7.944582e-11, 7.973353e-11, 
    7.86536e-11, 7.921954e-11, 7.833292e-11, 7.859991e-11, 7.878546e-11, 
    7.870406e-11, 7.912675e-11, 7.922638e-11, 7.963123e-11, 7.942194e-11, 
    8.06679e-11, 8.011666e-11, 8.164626e-11, 8.121881e-11, 7.83358e-11, 
    7.847115e-11, 7.894225e-11, 7.87181e-11, 7.935911e-11, 7.951689e-11, 
    7.964515e-11, 7.980912e-11, 7.982681e-11, 7.992396e-11, 7.976476e-11, 
    7.991767e-11, 7.933925e-11, 7.959773e-11, 7.88884e-11, 7.906105e-11, 
    7.898162e-11, 7.88945e-11, 7.916338e-11, 7.944985e-11, 7.945596e-11, 
    7.954782e-11, 7.98067e-11, 7.93617e-11, 8.073907e-11, 7.988846e-11, 
    7.861876e-11, 7.887949e-11, 7.891671e-11, 7.881572e-11, 7.950107e-11, 
    7.925274e-11, 7.992159e-11, 7.974083e-11, 8.0037e-11, 7.988983e-11, 
    7.986817e-11, 7.967915e-11, 7.956146e-11, 7.926414e-11, 7.902221e-11, 
    7.883037e-11, 7.887497e-11, 7.908571e-11, 7.946737e-11, 7.982842e-11, 
    7.974933e-11, 8.00145e-11, 7.931263e-11, 7.960694e-11, 7.949319e-11, 
    7.978979e-11, 7.91399e-11, 7.969335e-11, 7.899843e-11, 7.905936e-11, 
    7.924782e-11, 7.962691e-11, 7.971077e-11, 7.980032e-11, 7.974506e-11, 
    7.947706e-11, 7.943315e-11, 7.924324e-11, 7.919081e-11, 7.904609e-11, 
    7.892628e-11, 7.903575e-11, 7.915071e-11, 7.947717e-11, 7.977137e-11, 
    8.009213e-11, 8.017062e-11, 8.054542e-11, 8.024034e-11, 8.074381e-11, 
    8.031579e-11, 8.10567e-11, 7.97254e-11, 8.030317e-11, 7.925639e-11, 
    7.936916e-11, 7.957314e-11, 8.004097e-11, 7.978839e-11, 8.008377e-11, 
    7.943143e-11, 7.909299e-11, 7.900541e-11, 7.884203e-11, 7.900914e-11, 
    7.899555e-11, 7.915546e-11, 7.910407e-11, 7.948801e-11, 7.928178e-11, 
    7.986763e-11, 8.008143e-11, 8.068519e-11, 8.105532e-11, 8.143206e-11, 
    8.159839e-11, 8.164902e-11, 8.167018e-11 ;

 SOIL2C_vr =
  20.00645, 20.00647, 20.00646, 20.00648, 20.00647, 20.00648, 20.00645, 
    20.00647, 20.00646, 20.00645, 20.0065, 20.00648, 20.00653, 20.00651, 
    20.00655, 20.00653, 20.00656, 20.00655, 20.00657, 20.00657, 20.00659, 
    20.00657, 20.0066, 20.00659, 20.00659, 20.00657, 20.00648, 20.0065, 
    20.00648, 20.00648, 20.00648, 20.00647, 20.00646, 20.00645, 20.00645, 
    20.00646, 20.00648, 20.00648, 20.0065, 20.0065, 20.00652, 20.00651, 
    20.00655, 20.00654, 20.00657, 20.00656, 20.00657, 20.00657, 20.00657, 
    20.00656, 20.00656, 20.00655, 20.00651, 20.00652, 20.00649, 20.00647, 
    20.00645, 20.00644, 20.00644, 20.00645, 20.00646, 20.00647, 20.00648, 
    20.00649, 20.0065, 20.00652, 20.00653, 20.00655, 20.00654, 20.00655, 
    20.00656, 20.00657, 20.00657, 20.00657, 20.00655, 20.00657, 20.00654, 
    20.00655, 20.0065, 20.00648, 20.00647, 20.00646, 20.00645, 20.00646, 
    20.00645, 20.00646, 20.00647, 20.00647, 20.00649, 20.00648, 20.00653, 
    20.00651, 20.00656, 20.00655, 20.00656, 20.00655, 20.00657, 20.00655, 
    20.00657, 20.00658, 20.00658, 20.00659, 20.00655, 20.00657, 20.00647, 
    20.00647, 20.00647, 20.00646, 20.00646, 20.00645, 20.00646, 20.00646, 
    20.00647, 20.00648, 20.00648, 20.0065, 20.00651, 20.00653, 20.00655, 
    20.00656, 20.00655, 20.00656, 20.00655, 20.00655, 20.00658, 20.00656, 
    20.00659, 20.00658, 20.00657, 20.00658, 20.00647, 20.00647, 20.00645, 
    20.00646, 20.00645, 20.00646, 20.00646, 20.00648, 20.00649, 20.00649, 
    20.0065, 20.00651, 20.00653, 20.00654, 20.00656, 20.00656, 20.00656, 
    20.00656, 20.00655, 20.00656, 20.00657, 20.00656, 20.00658, 20.00658, 
    20.00658, 20.00658, 20.00647, 20.00647, 20.00647, 20.00648, 20.00647, 
    20.00649, 20.00649, 20.00652, 20.00651, 20.00653, 20.00651, 20.00651, 
    20.00653, 20.00651, 20.00654, 20.00652, 20.00656, 20.00654, 20.00656, 
    20.00656, 20.00657, 20.00657, 20.00658, 20.00659, 20.00659, 20.0066, 
    20.00648, 20.00649, 20.00649, 20.00649, 20.0065, 20.00651, 20.00653, 
    20.00653, 20.00654, 20.00654, 20.00652, 20.00653, 20.00649, 20.0065, 
    20.0065, 20.00648, 20.00653, 20.0065, 20.00655, 20.00653, 20.00657, 
    20.00655, 20.00659, 20.0066, 20.00662, 20.00664, 20.00649, 20.00649, 
    20.0065, 20.00651, 20.00652, 20.00653, 20.00654, 20.00654, 20.00655, 
    20.00655, 20.00654, 20.00655, 20.0065, 20.00653, 20.00648, 20.0065, 
    20.00651, 20.0065, 20.00653, 20.00653, 20.00655, 20.00654, 20.0066, 
    20.00657, 20.00665, 20.00663, 20.00648, 20.00649, 20.00652, 20.0065, 
    20.00654, 20.00654, 20.00655, 20.00656, 20.00656, 20.00656, 20.00656, 
    20.00656, 20.00653, 20.00655, 20.00651, 20.00652, 20.00652, 20.00651, 
    20.00653, 20.00654, 20.00654, 20.00655, 20.00656, 20.00654, 20.0066, 
    20.00656, 20.0065, 20.00651, 20.00651, 20.00651, 20.00654, 20.00653, 
    20.00656, 20.00656, 20.00657, 20.00656, 20.00656, 20.00655, 20.00655, 
    20.00653, 20.00652, 20.00651, 20.00651, 20.00652, 20.00654, 20.00656, 
    20.00656, 20.00657, 20.00653, 20.00655, 20.00654, 20.00656, 20.00653, 
    20.00655, 20.00652, 20.00652, 20.00653, 20.00655, 20.00655, 20.00656, 
    20.00656, 20.00654, 20.00654, 20.00653, 20.00653, 20.00652, 20.00652, 
    20.00652, 20.00653, 20.00654, 20.00656, 20.00657, 20.00658, 20.00659, 
    20.00658, 20.0066, 20.00658, 20.00662, 20.00655, 20.00658, 20.00653, 
    20.00654, 20.00655, 20.00657, 20.00656, 20.00657, 20.00654, 20.00652, 
    20.00652, 20.00651, 20.00652, 20.00652, 20.00653, 20.00652, 20.00654, 
    20.00653, 20.00656, 20.00657, 20.0066, 20.00662, 20.00664, 20.00665, 
    20.00665, 20.00665,
  20.00607, 20.0061, 20.00609, 20.00611, 20.0061, 20.00611, 20.00608, 
    20.0061, 20.00608, 20.00607, 20.00615, 20.00611, 20.00618, 20.00616, 
    20.00621, 20.00618, 20.00622, 20.00621, 20.00624, 20.00623, 20.00626, 
    20.00624, 20.00628, 20.00626, 20.00626, 20.00624, 20.00612, 20.00614, 
    20.00611, 20.00612, 20.00612, 20.0061, 20.00609, 20.00607, 20.00607, 
    20.00609, 20.00612, 20.00611, 20.00614, 20.00614, 20.00617, 20.00615, 
    20.0062, 20.00619, 20.00623, 20.00622, 20.00623, 20.00623, 20.00623, 
    20.00622, 20.00622, 20.00621, 20.00616, 20.00617, 20.00612, 20.0061, 
    20.00608, 20.00607, 20.00607, 20.00607, 20.00609, 20.00611, 20.00612, 
    20.00613, 20.00614, 20.00616, 20.00618, 20.00621, 20.0062, 20.00621, 
    20.00622, 20.00624, 20.00623, 20.00624, 20.00621, 20.00623, 20.0062, 
    20.00621, 20.00614, 20.00611, 20.0061, 20.00609, 20.00607, 20.00608, 
    20.00608, 20.00609, 20.0061, 20.0061, 20.00613, 20.00612, 20.00618, 
    20.00615, 20.00622, 20.0062, 20.00622, 20.00621, 20.00623, 20.00621, 
    20.00624, 20.00625, 20.00624, 20.00626, 20.00621, 20.00623, 20.0061, 
    20.0061, 20.0061, 20.00609, 20.00609, 20.00607, 20.00608, 20.00609, 
    20.0061, 20.00611, 20.00612, 20.00614, 20.00616, 20.00618, 20.0062, 
    20.00622, 20.00621, 20.00622, 20.00621, 20.0062, 20.00624, 20.00622, 
    20.00626, 20.00625, 20.00624, 20.00625, 20.0061, 20.00609, 20.00608, 
    20.00609, 20.00607, 20.00608, 20.00609, 20.00612, 20.00612, 20.00613, 
    20.00614, 20.00615, 20.00618, 20.0062, 20.00622, 20.00622, 20.00622, 
    20.00622, 20.00621, 20.00623, 20.00623, 20.00622, 20.00625, 20.00624, 
    20.00625, 20.00625, 20.0061, 20.0061, 20.0061, 20.00611, 20.0061, 
    20.00613, 20.00613, 20.00617, 20.00615, 20.00618, 20.00616, 20.00616, 
    20.00618, 20.00616, 20.0062, 20.00617, 20.00622, 20.0062, 20.00623, 
    20.00622, 20.00623, 20.00624, 20.00625, 20.00627, 20.00626, 20.00628, 
    20.00611, 20.00612, 20.00612, 20.00613, 20.00614, 20.00616, 20.00619, 
    20.00617, 20.00619, 20.0062, 20.00617, 20.00619, 20.00613, 20.00614, 
    20.00614, 20.00612, 20.00618, 20.00615, 20.0062, 20.00619, 20.00624, 
    20.00621, 20.00626, 20.00628, 20.0063, 20.00632, 20.00613, 20.00612, 
    20.00614, 20.00615, 20.00617, 20.00619, 20.00619, 20.00619, 20.0062, 
    20.00621, 20.0062, 20.00621, 20.00614, 20.00618, 20.00612, 20.00614, 
    20.00615, 20.00615, 20.00617, 20.00618, 20.00621, 20.00619, 20.00628, 
    20.00624, 20.00634, 20.00631, 20.00612, 20.00613, 20.00616, 20.00615, 
    20.00619, 20.0062, 20.00621, 20.00622, 20.00622, 20.00623, 20.00622, 
    20.00623, 20.00619, 20.0062, 20.00616, 20.00617, 20.00616, 20.00616, 
    20.00618, 20.0062, 20.0062, 20.0062, 20.00622, 20.00619, 20.00628, 
    20.00622, 20.00614, 20.00616, 20.00616, 20.00615, 20.0062, 20.00618, 
    20.00623, 20.00621, 20.00623, 20.00622, 20.00622, 20.00621, 20.0062, 
    20.00618, 20.00617, 20.00616, 20.00616, 20.00617, 20.0062, 20.00622, 
    20.00621, 20.00623, 20.00619, 20.00621, 20.0062, 20.00622, 20.00617, 
    20.00621, 20.00616, 20.00617, 20.00618, 20.00621, 20.00621, 20.00622, 
    20.00621, 20.0062, 20.00619, 20.00618, 20.00618, 20.00617, 20.00616, 
    20.00617, 20.00618, 20.0062, 20.00622, 20.00624, 20.00624, 20.00627, 
    20.00625, 20.00628, 20.00625, 20.0063, 20.00621, 20.00625, 20.00618, 
    20.00619, 20.0062, 20.00624, 20.00622, 20.00624, 20.00619, 20.00617, 
    20.00617, 20.00616, 20.00617, 20.00616, 20.00618, 20.00617, 20.0062, 
    20.00618, 20.00622, 20.00624, 20.00628, 20.0063, 20.00633, 20.00634, 
    20.00634, 20.00634,
  20.00552, 20.00554, 20.00554, 20.00556, 20.00555, 20.00556, 20.00553, 
    20.00555, 20.00553, 20.00552, 20.0056, 20.00556, 20.00564, 20.00561, 
    20.00567, 20.00563, 20.00568, 20.00567, 20.0057, 20.00569, 20.00573, 
    20.0057, 20.00574, 20.00572, 20.00572, 20.0057, 20.00557, 20.00559, 
    20.00557, 20.00557, 20.00557, 20.00555, 20.00554, 20.00552, 20.00552, 
    20.00554, 20.00557, 20.00556, 20.00559, 20.00559, 20.00562, 20.00561, 
    20.00566, 20.00565, 20.00569, 20.00568, 20.00569, 20.00569, 20.00569, 
    20.00567, 20.00568, 20.00567, 20.00561, 20.00563, 20.00558, 20.00555, 
    20.00553, 20.00551, 20.00551, 20.00552, 20.00554, 20.00556, 20.00557, 
    20.00558, 20.00559, 20.00562, 20.00563, 20.00566, 20.00566, 20.00567, 
    20.00568, 20.0057, 20.00569, 20.0057, 20.00567, 20.00569, 20.00566, 
    20.00566, 20.00559, 20.00556, 20.00555, 20.00554, 20.00552, 20.00553, 
    20.00553, 20.00554, 20.00555, 20.00555, 20.00558, 20.00557, 20.00563, 
    20.0056, 20.00568, 20.00566, 20.00568, 20.00567, 20.00569, 20.00567, 
    20.0057, 20.00571, 20.0057, 20.00572, 20.00567, 20.00569, 20.00555, 
    20.00555, 20.00555, 20.00554, 20.00554, 20.00552, 20.00553, 20.00554, 
    20.00555, 20.00556, 20.00557, 20.00559, 20.00561, 20.00564, 20.00566, 
    20.00567, 20.00567, 20.00567, 20.00566, 20.00566, 20.0057, 20.00568, 
    20.00572, 20.00572, 20.0057, 20.00572, 20.00555, 20.00554, 20.00553, 
    20.00554, 20.00552, 20.00553, 20.00554, 20.00557, 20.00558, 20.00558, 
    20.00559, 20.00561, 20.00563, 20.00566, 20.00568, 20.00568, 20.00568, 
    20.00568, 20.00567, 20.00568, 20.00569, 20.00568, 20.00572, 20.0057, 
    20.00572, 20.00571, 20.00555, 20.00555, 20.00555, 20.00556, 20.00555, 
    20.00558, 20.00559, 20.00562, 20.00561, 20.00563, 20.00561, 20.00561, 
    20.00563, 20.00561, 20.00566, 20.00562, 20.00568, 20.00565, 20.00568, 
    20.00568, 20.00569, 20.0057, 20.00571, 20.00573, 20.00572, 20.00574, 
    20.00557, 20.00558, 20.00558, 20.00559, 20.0056, 20.00561, 20.00564, 
    20.00563, 20.00565, 20.00565, 20.00562, 20.00564, 20.00558, 20.00559, 
    20.00559, 20.00557, 20.00563, 20.0056, 20.00566, 20.00564, 20.0057, 
    20.00567, 20.00572, 20.00574, 20.00576, 20.00579, 20.00558, 20.00558, 
    20.00559, 20.00561, 20.00562, 20.00564, 20.00565, 20.00565, 20.00566, 
    20.00567, 20.00565, 20.00567, 20.0056, 20.00564, 20.00557, 20.00559, 
    20.00561, 20.0056, 20.00563, 20.00564, 20.00566, 20.00565, 20.00574, 
    20.0057, 20.00581, 20.00578, 20.00557, 20.00558, 20.00562, 20.0056, 
    20.00565, 20.00566, 20.00567, 20.00568, 20.00568, 20.00569, 20.00567, 
    20.00569, 20.00564, 20.00566, 20.00561, 20.00562, 20.00562, 20.00561, 
    20.00563, 20.00565, 20.00565, 20.00566, 20.00568, 20.00565, 20.00574, 
    20.00568, 20.00559, 20.00561, 20.00562, 20.00561, 20.00566, 20.00564, 
    20.00569, 20.00567, 20.00569, 20.00568, 20.00568, 20.00567, 20.00566, 
    20.00564, 20.00562, 20.00561, 20.00561, 20.00563, 20.00565, 20.00568, 
    20.00567, 20.00569, 20.00564, 20.00566, 20.00566, 20.00568, 20.00563, 
    20.00567, 20.00562, 20.00562, 20.00564, 20.00566, 20.00567, 20.00568, 
    20.00567, 20.00565, 20.00565, 20.00564, 20.00563, 20.00562, 20.00562, 
    20.00562, 20.00563, 20.00565, 20.00567, 20.0057, 20.0057, 20.00573, 
    20.00571, 20.00574, 20.00571, 20.00577, 20.00567, 20.00571, 20.00564, 
    20.00565, 20.00566, 20.00569, 20.00568, 20.0057, 20.00565, 20.00563, 
    20.00562, 20.00561, 20.00562, 20.00562, 20.00563, 20.00563, 20.00566, 
    20.00564, 20.00568, 20.0057, 20.00574, 20.00577, 20.00579, 20.0058, 
    20.00581, 20.00581,
  20.00508, 20.00511, 20.0051, 20.00512, 20.00511, 20.00512, 20.00509, 
    20.00511, 20.00509, 20.00508, 20.00516, 20.00512, 20.0052, 20.00517, 
    20.00523, 20.00519, 20.00524, 20.00523, 20.00526, 20.00525, 20.00528, 
    20.00526, 20.0053, 20.00528, 20.00528, 20.00526, 20.00513, 20.00515, 
    20.00513, 20.00513, 20.00513, 20.00511, 20.0051, 20.00508, 20.00508, 
    20.0051, 20.00513, 20.00512, 20.00515, 20.00515, 20.00518, 20.00517, 
    20.00522, 20.00521, 20.00525, 20.00524, 20.00525, 20.00525, 20.00525, 
    20.00523, 20.00524, 20.00522, 20.00517, 20.00519, 20.00514, 20.00511, 
    20.00509, 20.00507, 20.00508, 20.00508, 20.0051, 20.00512, 20.00513, 
    20.00514, 20.00515, 20.00518, 20.00519, 20.00522, 20.00522, 20.00523, 
    20.00524, 20.00525, 20.00525, 20.00526, 20.00523, 20.00525, 20.00521, 
    20.00522, 20.00515, 20.00512, 20.00511, 20.0051, 20.00508, 20.00509, 
    20.00509, 20.0051, 20.00511, 20.00511, 20.00514, 20.00513, 20.00519, 
    20.00516, 20.00524, 20.00522, 20.00524, 20.00523, 20.00525, 20.00523, 
    20.00526, 20.00527, 20.00526, 20.00528, 20.00523, 20.00525, 20.00511, 
    20.00511, 20.00511, 20.0051, 20.00509, 20.00508, 20.00509, 20.0051, 
    20.00511, 20.00512, 20.00513, 20.00515, 20.00517, 20.0052, 20.00522, 
    20.00523, 20.00522, 20.00523, 20.00522, 20.00522, 20.00526, 20.00524, 
    20.00528, 20.00527, 20.00526, 20.00527, 20.00511, 20.0051, 20.00509, 
    20.0051, 20.00508, 20.00509, 20.0051, 20.00513, 20.00513, 20.00514, 
    20.00515, 20.00517, 20.00519, 20.00522, 20.00524, 20.00524, 20.00524, 
    20.00524, 20.00523, 20.00524, 20.00525, 20.00524, 20.00527, 20.00526, 
    20.00527, 20.00527, 20.00511, 20.00511, 20.00511, 20.00512, 20.00511, 
    20.00514, 20.00515, 20.00518, 20.00517, 20.00519, 20.00517, 20.00517, 
    20.00519, 20.00517, 20.00521, 20.00518, 20.00524, 20.00521, 20.00524, 
    20.00524, 20.00525, 20.00526, 20.00527, 20.00529, 20.00528, 20.0053, 
    20.00513, 20.00514, 20.00514, 20.00515, 20.00516, 20.00517, 20.0052, 
    20.00519, 20.00521, 20.00521, 20.00518, 20.0052, 20.00514, 20.00515, 
    20.00515, 20.00513, 20.00519, 20.00516, 20.00522, 20.0052, 20.00525, 
    20.00523, 20.00528, 20.0053, 20.00532, 20.00535, 20.00514, 20.00513, 
    20.00515, 20.00517, 20.00518, 20.0052, 20.00521, 20.00521, 20.00522, 
    20.00523, 20.00521, 20.00523, 20.00516, 20.0052, 20.00513, 20.00515, 
    20.00517, 20.00516, 20.00519, 20.0052, 20.00522, 20.00521, 20.0053, 
    20.00526, 20.00537, 20.00533, 20.00513, 20.00514, 20.00517, 20.00516, 
    20.00521, 20.00522, 20.00522, 20.00524, 20.00524, 20.00524, 20.00523, 
    20.00524, 20.0052, 20.00522, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00519, 20.00521, 20.00521, 20.00522, 20.00524, 20.00521, 20.0053, 
    20.00524, 20.00515, 20.00517, 20.00517, 20.00517, 20.00521, 20.0052, 
    20.00524, 20.00523, 20.00525, 20.00524, 20.00524, 20.00523, 20.00522, 
    20.0052, 20.00518, 20.00517, 20.00517, 20.00519, 20.00521, 20.00524, 
    20.00523, 20.00525, 20.0052, 20.00522, 20.00521, 20.00524, 20.00519, 
    20.00523, 20.00518, 20.00518, 20.0052, 20.00522, 20.00523, 20.00524, 
    20.00523, 20.00521, 20.00521, 20.0052, 20.00519, 20.00518, 20.00517, 
    20.00518, 20.00519, 20.00521, 20.00523, 20.00526, 20.00526, 20.00529, 
    20.00527, 20.0053, 20.00527, 20.00532, 20.00523, 20.00527, 20.0052, 
    20.00521, 20.00522, 20.00525, 20.00524, 20.00525, 20.00521, 20.00519, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00519, 20.00519, 20.00521, 
    20.0052, 20.00524, 20.00525, 20.0053, 20.00532, 20.00535, 20.00536, 
    20.00537, 20.00537,
  20.00437, 20.00439, 20.00439, 20.0044, 20.00439, 20.00441, 20.00438, 
    20.00439, 20.00438, 20.00437, 20.00444, 20.0044, 20.00447, 20.00445, 
    20.0045, 20.00447, 20.00451, 20.0045, 20.00452, 20.00451, 20.00454, 
    20.00452, 20.00456, 20.00454, 20.00454, 20.00452, 20.00441, 20.00443, 
    20.00441, 20.00441, 20.00441, 20.00439, 20.00439, 20.00437, 20.00437, 
    20.00438, 20.00441, 20.0044, 20.00443, 20.00443, 20.00446, 20.00444, 
    20.00449, 20.00448, 20.00451, 20.00451, 20.00451, 20.00451, 20.00451, 
    20.0045, 20.00451, 20.00449, 20.00445, 20.00446, 20.00442, 20.00439, 
    20.00438, 20.00436, 20.00437, 20.00437, 20.00438, 20.0044, 20.00441, 
    20.00442, 20.00443, 20.00445, 20.00447, 20.00449, 20.00449, 20.0045, 
    20.0045, 20.00452, 20.00451, 20.00452, 20.0045, 20.00451, 20.00448, 
    20.00449, 20.00443, 20.00441, 20.0044, 20.00439, 20.00437, 20.00438, 
    20.00438, 20.00439, 20.0044, 20.00439, 20.00442, 20.00441, 20.00447, 
    20.00444, 20.0045, 20.00449, 20.00451, 20.0045, 20.00451, 20.0045, 
    20.00452, 20.00453, 20.00452, 20.00454, 20.0045, 20.00451, 20.00439, 
    20.00439, 20.0044, 20.00438, 20.00438, 20.00437, 20.00438, 20.00439, 
    20.0044, 20.00441, 20.00441, 20.00443, 20.00445, 20.00447, 20.00449, 
    20.0045, 20.00449, 20.0045, 20.00449, 20.00449, 20.00453, 20.00451, 
    20.00454, 20.00454, 20.00452, 20.00454, 20.00439, 20.00439, 20.00438, 
    20.00439, 20.00437, 20.00438, 20.00439, 20.00441, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00447, 20.00449, 20.0045, 20.0045, 20.0045, 
    20.00451, 20.0045, 20.00451, 20.00451, 20.00451, 20.00454, 20.00453, 
    20.00454, 20.00453, 20.00439, 20.0044, 20.0044, 20.0044, 20.0044, 
    20.00442, 20.00443, 20.00446, 20.00444, 20.00446, 20.00445, 20.00445, 
    20.00447, 20.00445, 20.00449, 20.00446, 20.00451, 20.00448, 20.00451, 
    20.0045, 20.00451, 20.00452, 20.00453, 20.00455, 20.00454, 20.00456, 
    20.00441, 20.00442, 20.00442, 20.00443, 20.00443, 20.00445, 20.00447, 
    20.00446, 20.00448, 20.00448, 20.00446, 20.00447, 20.00443, 20.00443, 
    20.00443, 20.00441, 20.00447, 20.00444, 20.00449, 20.00447, 20.00452, 
    20.0045, 20.00454, 20.00456, 20.00458, 20.0046, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00446, 20.00447, 20.00448, 20.00448, 20.00449, 
    20.0045, 20.00448, 20.0045, 20.00443, 20.00447, 20.00442, 20.00443, 
    20.00444, 20.00444, 20.00446, 20.00447, 20.00449, 20.00448, 20.00455, 
    20.00452, 20.00461, 20.00459, 20.00442, 20.00442, 20.00445, 20.00444, 
    20.00448, 20.00449, 20.00449, 20.0045, 20.0045, 20.00451, 20.0045, 
    20.00451, 20.00447, 20.00449, 20.00445, 20.00446, 20.00445, 20.00445, 
    20.00447, 20.00448, 20.00448, 20.00449, 20.0045, 20.00448, 20.00456, 
    20.00451, 20.00443, 20.00445, 20.00445, 20.00444, 20.00448, 20.00447, 
    20.00451, 20.0045, 20.00452, 20.00451, 20.00451, 20.0045, 20.00449, 
    20.00447, 20.00446, 20.00444, 20.00445, 20.00446, 20.00448, 20.0045, 
    20.0045, 20.00451, 20.00447, 20.00449, 20.00448, 20.0045, 20.00446, 
    20.0045, 20.00446, 20.00446, 20.00447, 20.00449, 20.0045, 20.0045, 
    20.0045, 20.00448, 20.00448, 20.00447, 20.00447, 20.00446, 20.00445, 
    20.00446, 20.00446, 20.00448, 20.0045, 20.00452, 20.00452, 20.00455, 
    20.00453, 20.00456, 20.00453, 20.00458, 20.0045, 20.00453, 20.00447, 
    20.00448, 20.00449, 20.00452, 20.0045, 20.00452, 20.00448, 20.00446, 
    20.00446, 20.00445, 20.00446, 20.00445, 20.00446, 20.00446, 20.00448, 
    20.00447, 20.00451, 20.00452, 20.00455, 20.00458, 20.0046, 20.00461, 
    20.00461, 20.00461,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258222, 0.5258228, 0.5258227, 0.5258232, 0.5258229, 0.5258232, 
    0.5258223, 0.5258228, 0.5258225, 0.5258223, 0.5258241, 0.5258232, 
    0.525825, 0.5258244, 0.5258259, 0.5258249, 0.525826, 0.5258258, 
    0.5258265, 0.5258263, 0.5258271, 0.5258265, 0.5258275, 0.525827, 
    0.5258271, 0.5258265, 0.5258234, 0.525824, 0.5258234, 0.5258234, 
    0.5258234, 0.5258229, 0.5258227, 0.5258222, 0.5258223, 0.5258226, 
    0.5258235, 0.5258232, 0.5258239, 0.5258238, 0.5258246, 0.5258243, 
    0.5258256, 0.5258252, 0.5258263, 0.525826, 0.5258263, 0.5258262, 
    0.5258263, 0.5258259, 0.525826, 0.5258257, 0.5258244, 0.5258247, 
    0.5258235, 0.5258229, 0.5258224, 0.525822, 0.5258221, 0.5258222, 
    0.5258226, 0.5258231, 0.5258234, 0.5258237, 0.5258238, 0.5258245, 
    0.5258248, 0.5258257, 0.5258255, 0.5258257, 0.525826, 0.5258263, 
    0.5258263, 0.5258265, 0.5258257, 0.5258262, 0.5258254, 0.5258256, 
    0.5258239, 0.5258232, 0.525823, 0.5258227, 0.5258221, 0.5258225, 
    0.5258224, 0.5258228, 0.525823, 0.5258229, 0.5258237, 0.5258234, 
    0.5258249, 0.5258242, 0.525826, 0.5258256, 0.525826, 0.5258258, 
    0.5258262, 0.5258259, 0.5258265, 0.5258267, 0.5258266, 0.525827, 
    0.5258258, 0.5258263, 0.5258229, 0.5258229, 0.525823, 0.5258226, 
    0.5258226, 0.5258222, 0.5258225, 0.5258226, 0.525823, 0.5258232, 
    0.5258234, 0.5258239, 0.5258244, 0.5258251, 0.5258256, 0.5258259, 
    0.5258257, 0.5258259, 0.5258257, 0.5258256, 0.5258266, 0.525826, 
    0.5258269, 0.5258269, 0.5258265, 0.5258269, 0.5258229, 0.5258228, 
    0.5258224, 0.5258227, 0.5258222, 0.5258225, 0.5258226, 0.5258234, 
    0.5258235, 0.5258237, 0.525824, 0.5258243, 0.5258249, 0.5258255, 
    0.525826, 0.525826, 0.525826, 0.5258261, 0.5258258, 0.5258262, 0.5258262, 
    0.525826, 0.5258269, 0.5258266, 0.5258269, 0.5258267, 0.5258228, 
    0.5258231, 0.5258229, 0.5258231, 0.525823, 0.5258236, 0.5258238, 
    0.5258247, 0.5258243, 0.5258248, 0.5258244, 0.5258244, 0.5258248, 
    0.5258244, 0.5258254, 0.5258247, 0.5258261, 0.5258254, 0.5258262, 
    0.525826, 0.5258262, 0.5258265, 0.5258267, 0.5258272, 0.5258271, 
    0.5258275, 0.5258233, 0.5258236, 0.5258235, 0.5258238, 0.525824, 
    0.5258244, 0.5258251, 0.5258248, 0.5258253, 0.5258254, 0.5258247, 
    0.5258251, 0.5258237, 0.525824, 0.5258238, 0.5258234, 0.5258249, 
    0.5258241, 0.5258256, 0.5258251, 0.5258264, 0.5258258, 0.525827, 
    0.5258275, 0.525828, 0.5258286, 0.5258237, 0.5258235, 0.5258238, 
    0.5258242, 0.5258247, 0.5258251, 0.5258252, 0.5258253, 0.5258256, 
    0.5258258, 0.5258253, 0.5258259, 0.525824, 0.525825, 0.5258235, 0.525824, 
    0.5258242, 0.5258241, 0.5258248, 0.525825, 0.5258257, 0.5258253, 
    0.5258274, 0.5258265, 0.5258291, 0.5258284, 0.5258235, 0.5258237, 
    0.5258245, 0.5258241, 0.5258252, 0.5258254, 0.5258257, 0.525826, 
    0.525826, 0.5258262, 0.5258259, 0.5258262, 0.5258251, 0.5258256, 
    0.5258244, 0.5258247, 0.5258245, 0.5258244, 0.5258248, 0.5258254, 
    0.5258254, 0.5258255, 0.525826, 0.5258252, 0.5258275, 0.5258261, 
    0.525824, 0.5258244, 0.5258244, 0.5258243, 0.5258254, 0.525825, 
    0.5258262, 0.5258259, 0.5258263, 0.5258261, 0.525826, 0.5258257, 
    0.5258256, 0.525825, 0.5258246, 0.5258243, 0.5258244, 0.5258247, 
    0.5258254, 0.525826, 0.5258259, 0.5258263, 0.5258251, 0.5258256, 
    0.5258254, 0.5258259, 0.5258248, 0.5258257, 0.5258246, 0.5258247, 
    0.525825, 0.5258257, 0.5258258, 0.5258259, 0.5258259, 0.5258254, 
    0.5258253, 0.525825, 0.5258249, 0.5258247, 0.5258245, 0.5258247, 
    0.5258248, 0.5258254, 0.5258259, 0.5258265, 0.5258266, 0.5258272, 
    0.5258267, 0.5258275, 0.5258268, 0.5258281, 0.5258258, 0.5258268, 
    0.525825, 0.5258252, 0.5258256, 0.5258263, 0.5258259, 0.5258264, 
    0.5258253, 0.5258247, 0.5258246, 0.5258243, 0.5258246, 0.5258246, 
    0.5258248, 0.5258248, 0.5258254, 0.5258251, 0.525826, 0.5258264, 
    0.5258274, 0.5258281, 0.5258287, 0.525829, 0.5258291, 0.5258291 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  2.569961e-21, 7.709882e-21, -1.28498e-20, 1.003089e-36, 5.139921e-21, 
    2.569961e-21, 2.569961e-20, -1.28498e-20, -1.003089e-36, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, 0, 
    -2.569961e-21, -2.055969e-20, 5.139921e-21, 5.139921e-21, -1.003089e-36, 
    5.139921e-21, 7.709882e-21, 7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -1.541976e-20, 1.798972e-20, 2.569961e-21, 5.139921e-21, 1.541976e-20, 
    1.28498e-20, -1.541976e-20, 0, -7.709882e-21, -1.28498e-20, 2.569961e-21, 
    1.541976e-20, 1.027984e-20, 1.541976e-20, -1.003089e-36, -2.569961e-21, 
    -7.709882e-21, 7.709882e-21, -2.055969e-20, -7.709882e-21, -1.28498e-20, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, -1.027984e-20, 1.28498e-20, 
    5.139921e-21, 1.027984e-20, -1.027984e-20, 2.055969e-20, 5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -1.28498e-20, 7.709882e-21, 1.003089e-36, 
    5.139921e-21, -7.709882e-21, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, -1.541976e-20, 5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 1.027984e-20, 2.055969e-20, 5.139921e-21, 
    1.798972e-20, -1.027984e-20, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    1.027984e-20, -5.139921e-21, 2.569961e-21, -2.055969e-20, -1.28498e-20, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, -7.709882e-21, 7.709882e-21, 
    1.027984e-20, 1.003089e-36, -1.027984e-20, 2.569961e-21, 1.003089e-36, 
    -1.027984e-20, -5.139921e-21, -5.139921e-21, -2.569961e-21, 1.541976e-20, 
    1.28498e-20, -5.139921e-21, 7.709882e-21, -2.569961e-21, 7.709882e-21, 
    -1.003089e-36, -1.027984e-20, -2.055969e-20, -1.541976e-20, 
    -2.055969e-20, 5.139921e-21, 1.027984e-20, 1.027984e-20, -1.28498e-20, 
    -7.709882e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, -7.709882e-21, 1.003089e-36, 1.541976e-20, 7.709882e-21, 
    5.139921e-21, 1.541976e-20, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    7.709882e-21, -1.003089e-36, 2.569961e-21, 2.569961e-21, -2.055969e-20, 
    -1.027984e-20, 0, 5.139921e-21, -1.027984e-20, 1.003089e-36, 
    -1.28498e-20, 0, 2.569961e-21, 2.569961e-21, 2.569961e-21, -1.027984e-20, 
    -7.709882e-21, -1.541976e-20, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    2.312965e-20, -7.709882e-21, 7.709882e-21, 0, 7.709882e-21, 1.541976e-20, 
    -1.798972e-20, -1.027984e-20, -1.541976e-20, -2.569961e-21, 5.139921e-21, 
    -1.28498e-20, 7.709882e-21, 1.003089e-36, 2.569961e-21, 5.139921e-21, 
    -1.027984e-20, -1.541976e-20, -2.569961e-21, 5.139921e-21, 7.709882e-21, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, -1.28498e-20, 
    -1.28498e-20, 2.569961e-21, -1.003089e-36, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, -1.28498e-20, -1.027984e-20, 
    -2.312965e-20, -1.28498e-20, 2.569961e-21, -5.139921e-21, -1.027984e-20, 
    -2.569961e-21, 1.027984e-20, 1.003089e-36, -1.027984e-20, -2.569961e-21, 
    1.541976e-20, -5.139921e-21, 2.569961e-21, -1.003089e-36, -5.139921e-21, 
    0, -2.569961e-21, 1.28498e-20, 2.569961e-21, -1.798972e-20, 
    -2.569961e-21, 2.055969e-20, -7.709882e-21, 7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 1.027984e-20, -7.709882e-21, -1.027984e-20, -7.709882e-21, 
    -1.28498e-20, 1.027984e-20, -1.798972e-20, 5.139921e-21, -1.027984e-20, 
    2.569961e-21, -2.055969e-20, 5.139921e-21, -2.569961e-21, 0, 
    7.709882e-21, 1.541976e-20, -3.009266e-36, -2.569961e-21, 1.003089e-36, 
    7.709882e-21, 2.569961e-21, 1.798972e-20, 1.003089e-36, -1.541976e-20, 
    5.139921e-21, -5.139921e-21, -7.709882e-21, 0, -7.709882e-21, 
    7.709882e-21, 0, 1.027984e-20, -7.709882e-21, 1.003089e-36, 
    -1.541976e-20, 2.055969e-20, -5.139921e-21, 7.709882e-21, 1.28498e-20, 
    -1.027984e-20, 5.139921e-21, 0, 1.027984e-20, 1.541976e-20, 
    -7.709882e-21, 1.28498e-20, -1.541976e-20, -2.569961e-21, -2.569961e-21, 
    -1.798972e-20, -5.139921e-21, -1.003089e-36, 2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -2.312965e-20, -5.139921e-21, -1.027984e-20, 
    -1.003089e-36, -1.541976e-20, 2.569961e-21, 2.826957e-20, -1.541976e-20, 
    2.569961e-21, -1.28498e-20, 5.139921e-21, -5.139921e-21, -1.28498e-20, 
    -1.28498e-20, -7.709882e-21, -1.027984e-20, -1.027984e-20, -2.569961e-21, 
    2.569961e-21, 7.709882e-21, -2.569961e-21, -2.312965e-20, 3.009266e-36, 
    7.709882e-21, -1.28498e-20, 1.003089e-36, -7.709882e-21, -1.003089e-36, 
    2.569961e-21, 7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -2.055969e-20, -5.139921e-21, 7.709882e-21, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -1.027984e-20, -1.28498e-20, -1.027984e-20, 
    1.798972e-20, 5.139921e-21, -2.569961e-21, 0, 1.003089e-36, 5.139921e-21, 
    -2.569961e-21, 1.541976e-20, 2.569961e-21, 7.709882e-21, 1.027984e-20, 0, 
    5.139921e-21, -7.709882e-21, -2.569961e-21, -1.28498e-20, -5.139921e-21, 
    0, -5.139921e-21, -7.709882e-21, -7.709882e-21, 2.569961e-21, 
    -1.28498e-20, 5.139921e-21, -2.569961e-21, 2.569961e-21,
  -7.709882e-21, 1.027984e-20, -7.709882e-21, -1.027984e-20, 5.139921e-21, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, 7.709882e-21, 7.709882e-21, 
    2.569961e-21, 0, -5.139921e-21, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -1.541976e-20, -1.003089e-36, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 0, 7.709882e-21, -2.569961e-21, -7.709882e-21, 0, 
    -2.569961e-21, 1.027984e-20, 2.055969e-20, 2.569961e-21, -1.027984e-20, 
    0, -5.139921e-21, 0, -1.541976e-20, -5.139921e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, 5.139921e-21, -7.709882e-21, 1.027984e-20, 
    -1.541976e-20, -2.569961e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    -7.709882e-21, 1.027984e-20, 1.28498e-20, 1.003089e-36, 5.139921e-21, 0, 
    7.709882e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, -1.541976e-20, 
    1.28498e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, -1.798972e-20, 2.569961e-21, 
    0, -2.569961e-21, 7.709882e-21, 1.541976e-20, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 0, 1.28498e-20, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, -5.139921e-21, 
    1.027984e-20, 2.569961e-21, 1.003089e-36, 1.798972e-20, 0, -1.027984e-20, 
    -7.709882e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, -1.003089e-36, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, 1.027984e-20, -7.709882e-21, 
    -7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, -1.28498e-20, 
    7.709882e-21, -5.139921e-21, 7.709882e-21, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, 7.709882e-21, -1.28498e-20, -1.798972e-20, 0, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, -7.709882e-21, 1.027984e-20, 7.709882e-21, 5.139921e-21, 
    1.027984e-20, -1.003089e-36, 2.569961e-21, 2.569961e-21, -1.003089e-36, 
    7.709882e-21, 0, 5.139921e-21, 1.28498e-20, -5.139921e-21, 1.28498e-20, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, 1.541976e-20, 5.139921e-21, -2.055969e-20, 0, 7.709882e-21, 
    0, 2.312965e-20, 2.569961e-21, -5.139921e-21, -7.709882e-21, 0, 
    -7.709882e-21, -2.569961e-21, -7.709882e-21, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    0, 5.139921e-21, 2.569961e-21, -2.569961e-21, 0, 2.569961e-21, 
    -1.798972e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, 
    1.28498e-20, 0, 7.709882e-21, -1.28498e-20, 0, -2.569961e-21, 
    -5.139921e-21, 1.798972e-20, 7.709882e-21, 2.569961e-21, -1.541976e-20, 
    1.027984e-20, 7.709882e-21, 5.139921e-21, 0, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, -1.003089e-36, -5.139921e-21, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, -1.28498e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -2.569961e-21, -1.003089e-36, -2.569961e-21, 5.139921e-21, 7.709882e-21, 
    0, -2.569961e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 7.709882e-21, 0, -1.027984e-20, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, 0, 0, 7.709882e-21, 2.569961e-21, 
    1.28498e-20, 5.139921e-21, -7.709882e-21, 7.709882e-21, 0, 7.709882e-21, 
    -7.709882e-21, -1.28498e-20, 0, -1.027984e-20, 7.709882e-21, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 0, -7.709882e-21, 5.139921e-21, 0, 
    -5.139921e-21, 7.709882e-21, -2.569961e-21, 0, 0, -5.139921e-21, 
    1.28498e-20, 2.569961e-21, 1.027984e-20, -7.709882e-21, 1.541976e-20, 
    1.798972e-20, 7.709882e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, 
    -1.027984e-20, -1.003089e-36, -2.569961e-21, -2.569961e-21, 1.027984e-20, 
    0, 2.055969e-20, 0, -1.798972e-20, 1.027984e-20, 2.569961e-21, 
    -1.541976e-20, 1.28498e-20, -5.139921e-21, 1.28498e-20, -7.709882e-21, 
    2.569961e-21, -5.139921e-21, 1.027984e-20, 0, -7.709882e-21, 
    5.139921e-21, 1.28498e-20, -7.709882e-21, 5.139921e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, 7.709882e-21, 5.139921e-21, 1.027984e-20, 
    -1.541976e-20, -1.003089e-36, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, 0,
  1.027984e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 1.28498e-20, 
    -1.28498e-20, -1.003089e-36, -1.003089e-36, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, 1.003089e-36, -5.139921e-21, -2.569961e-21, 7.709882e-21, 
    -1.003089e-36, 1.541976e-20, 7.709882e-21, 1.027984e-20, 1.28498e-20, 
    2.569961e-21, 1.541976e-20, -2.569961e-21, -5.139921e-21, 0, 1.28498e-20, 
    -7.709882e-21, 0, 0, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    2.569961e-21, -1.28498e-20, 2.569961e-21, 2.569961e-21, -2.569961e-20, 
    2.569961e-21, 1.027984e-20, 0, 1.027984e-20, -7.709882e-21, 0, 
    7.709882e-21, -2.569961e-21, -1.027984e-20, 0, 5.139921e-21, 
    1.003089e-36, 2.312965e-20, 1.003089e-36, -1.28498e-20, 0, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -2.055969e-20, 0, 1.027984e-20, 
    -1.027984e-20, 7.709882e-21, -1.541976e-20, -7.709882e-21, -5.139921e-21, 
    -5.139921e-21, -7.709882e-21, -7.709882e-21, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, -7.709882e-21, 
    -1.798972e-20, 1.28498e-20, 5.139921e-21, 2.569961e-21, 1.027984e-20, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, -5.139921e-21, -1.541976e-20, 
    7.709882e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 1.003089e-36, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, 1.798972e-20, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    2.569961e-21, -1.027984e-20, -1.798972e-20, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, -1.798972e-20, -1.027984e-20, -1.003089e-36, 0, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 1.003089e-36, 2.569961e-21, 1.027984e-20, 
    -2.569961e-21, 2.569961e-21, 0, 1.28498e-20, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 1.28498e-20, -1.003089e-36, 7.709882e-21, 
    0, -1.541976e-20, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -1.003089e-36, -7.709882e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 1.541976e-20, 5.139921e-21, 5.139921e-21, 
    -1.003089e-36, 0, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, -5.139921e-21, -1.003089e-36, 
    -5.139921e-21, 5.139921e-21, 7.709882e-21, 1.027984e-20, -1.003089e-36, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, -1.28498e-20, 
    -1.798972e-20, 7.709882e-21, 0, -7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    1.28498e-20, -1.027984e-20, 2.569961e-21, 1.28498e-20, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, -1.28498e-20, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, 1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -2.055969e-20, 1.027984e-20, 0, -1.003089e-36, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 7.709882e-21, 
    2.569961e-20, -1.027984e-20, 7.709882e-21, -2.569961e-21, -1.28498e-20, 
    -2.055969e-20, 5.139921e-21, 1.28498e-20, -1.027984e-20, -2.569961e-21, 
    1.798972e-20, -2.569961e-21, 5.139921e-21, 0, -3.340949e-20, 0, 
    1.003089e-36, -5.139921e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, 
    1.003089e-36, 2.569961e-21, -1.003089e-36, 7.709882e-21, 1.541976e-20, 0, 
    -1.027984e-20, -7.709882e-21, -2.569961e-21, -7.709882e-21, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, -2.569961e-21, 5.139921e-21, 7.709882e-21, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, -7.709882e-21, 0, 
    -1.28498e-20, -1.541976e-20, -1.541976e-20, -1.541976e-20, -1.541976e-20, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, 0, 0, 
    -5.139921e-21, -7.709882e-21, 1.28498e-20, 1.003089e-36, 2.569961e-21, 
    -2.569961e-21, -1.541976e-20, 7.709882e-21, 5.139921e-21, 2.055969e-20, 
    7.709882e-21, -2.569961e-21, -1.798972e-20, -1.28498e-20, 5.139921e-21, 
    7.709882e-21, -7.709882e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    1.003089e-36, 0, -1.541976e-20, -2.569961e-21, 1.003089e-36, 
    1.003089e-36, 1.027984e-20, 7.709882e-21, -5.139921e-21, 5.139921e-21, 
    -1.28498e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -1.541976e-20, 1.541976e-20, 0, 
    -1.027984e-20, 0, -1.027984e-20, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, -7.709882e-21, -5.139921e-21, 
    2.569961e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, 7.709882e-21, -1.003089e-36, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 0, 1.027984e-20, 1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 2.569961e-21, -5.139921e-21, -2.055969e-20, 
    -2.569961e-21, 5.139921e-21, 1.003089e-36, 1.003089e-36, 5.139921e-21, 
    5.139921e-21,
  1.28498e-20, 2.055969e-20, -5.139921e-21, 1.541976e-20, -1.541976e-20, 
    1.003089e-36, -1.28498e-20, 1.027984e-20, 1.003089e-36, 0, -1.541976e-20, 
    1.541976e-20, -1.027984e-20, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, 7.709882e-21, 1.027984e-20, 2.569961e-21, 
    -1.027984e-20, -2.312965e-20, -2.569961e-21, 5.139921e-21, 1.027984e-20, 
    -7.709882e-21, 5.139921e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, 
    -1.28498e-20, 1.28498e-20, 1.027984e-20, -5.139921e-21, -2.569961e-21, 
    2.569961e-20, -5.139921e-21, -7.709882e-21, -2.569961e-21, 1.027984e-20, 
    -7.709882e-21, -5.139921e-21, 1.28498e-20, 2.569961e-21, 7.709882e-21, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, 1.28498e-20, -1.28498e-20, 
    1.027984e-20, 1.003089e-36, -1.28498e-20, 5.139921e-21, 1.541976e-20, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, -2.569961e-21, -1.28498e-20, 
    2.055969e-20, 2.569961e-21, 2.312965e-20, -5.139921e-21, 1.798972e-20, 
    1.541976e-20, -5.139921e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, -5.139921e-21, -5.139921e-21, -1.28498e-20, 
    2.569961e-21, 1.541976e-20, -5.139921e-21, -1.541976e-20, -2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 1.003089e-36, 1.798972e-20, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 1.798972e-20, -1.003089e-36, -7.709882e-21, 
    1.28498e-20, -2.569961e-21, -7.709882e-21, -7.709882e-21, -2.569961e-21, 
    -7.709882e-21, -1.28498e-20, -2.569961e-21, -5.139921e-21, 1.798972e-20, 
    -1.798972e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, -1.541976e-20, 
    1.027984e-20, 7.709882e-21, 0, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    -1.003089e-36, -2.569961e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, 7.709882e-21, -1.541976e-20, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, 0, 
    -2.569961e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 1.28498e-20, 
    -7.709882e-21, 2.312965e-20, -7.709882e-21, 2.569961e-21, 1.003089e-36, 
    7.709882e-21, 5.139921e-21, -1.003089e-36, -7.709882e-21, 0, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, -1.28498e-20, 
    7.709882e-21, -2.055969e-20, -1.027984e-20, 2.569961e-21, -1.541976e-20, 
    -2.569961e-21, 0, -7.709882e-21, 1.003089e-36, 0, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, 2.569961e-21, 1.003089e-36, 
    0, -1.027984e-20, 2.569961e-21, 2.569961e-21, 7.709882e-21, 1.003089e-36, 
    1.027984e-20, 7.709882e-21, -5.139921e-21, -2.569961e-21, 1.798972e-20, 
    1.027984e-20, -1.027984e-20, 1.541976e-20, 1.798972e-20, 1.003089e-36, 
    -5.139921e-21, -7.709882e-21, 1.798972e-20, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, -1.027984e-20, -2.569961e-21, 0, 2.312965e-20, 
    -1.28498e-20, 2.569961e-21, -1.003089e-36, -7.709882e-21, -5.139921e-21, 
    -1.28498e-20, 1.027984e-20, -1.541976e-20, -1.28498e-20, -2.055969e-20, 
    0, 2.569961e-21, -1.28498e-20, -2.569961e-21, 2.569961e-21, 1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 1.28498e-20, 1.003089e-36, -7.709882e-21, 
    -7.709882e-21, -2.569961e-21, 7.709882e-21, -1.28498e-20, -5.139921e-21, 
    1.798972e-20, -7.709882e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 1.541976e-20, 7.709882e-21, -2.569961e-21, -1.003089e-36, 
    1.541976e-20, -2.569961e-21, -7.709882e-21, 0, 1.541976e-20, 
    2.569961e-21, -1.003089e-36, -1.798972e-20, 1.027984e-20, 5.139921e-21, 
    2.569961e-21, 1.28498e-20, 5.139921e-21, -7.709882e-21, 2.312965e-20, 
    1.28498e-20, -2.569961e-21, 1.28498e-20, 5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, -5.139921e-21, 0, 
    1.027984e-20, 2.569961e-21, 2.569961e-21, -1.541976e-20, -2.569961e-21, 
    -7.709882e-21, -1.027984e-20, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, -5.139921e-21, -1.541976e-20, 5.139921e-21, 2.569961e-21, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    5.139921e-21, -1.28498e-20, 1.28498e-20, 2.055969e-20, 5.139921e-21, 
    -1.003089e-36, 1.28498e-20, -7.709882e-21, -1.541976e-20, 0, 
    5.139921e-21, 2.569961e-21, -1.027984e-20, 7.709882e-21, 5.139921e-21, 
    -7.709882e-21, 1.28498e-20, -7.709882e-21, -1.28498e-20, -1.027984e-20, 
    -1.027984e-20, 7.709882e-21, -7.709882e-21, -2.569961e-21, 1.28498e-20, 
    1.28498e-20, 1.027984e-20, -2.569961e-21, -1.003089e-36, -1.003089e-36, 
    2.569961e-21, -5.139921e-21, -2.569961e-21, 1.003089e-36, 7.709882e-21, 
    7.709882e-21, 0, -1.003089e-36, -5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 2.569961e-21, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -1.003089e-36, -7.709882e-21, -1.027984e-20, 2.569961e-20, 0, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, 1.541976e-20, -1.027984e-20, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, -1.027984e-20, 0, -1.541976e-20,
  -7.709882e-21, 1.798972e-20, 2.569961e-21, -2.569961e-21, 1.798972e-20, 
    -2.569961e-21, 2.569961e-21, 7.709882e-21, 1.027984e-20, -1.28498e-20, 
    -2.569961e-21, -1.28498e-20, -1.541976e-20, 2.569961e-21, 2.055969e-20, 
    5.139921e-21, 5.139921e-21, -1.541976e-20, -2.569961e-21, 1.003089e-36, 
    -1.28498e-20, 2.569961e-21, 1.003089e-36, -1.003089e-36, 2.569961e-21, 
    1.003089e-36, -1.541976e-20, 1.027984e-20, -1.798972e-20, 7.709882e-21, 
    1.541976e-20, 5.139921e-21, 1.003089e-36, -1.28498e-20, -1.541976e-20, 
    -1.28498e-20, -1.504633e-36, -1.28498e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, -1.541976e-20, 7.709882e-21, 
    1.003089e-36, -7.709882e-21, 5.139921e-21, -2.569961e-21, 1.798972e-20, 
    1.798972e-20, -2.569961e-21, 1.027984e-20, -2.569961e-21, 1.027984e-20, 
    -7.709882e-21, 2.055969e-20, 0, 7.709882e-21, -7.709882e-21, 
    1.541976e-20, -1.798972e-20, 7.709882e-21, -5.139921e-21, -1.541976e-20, 
    1.027984e-20, -1.027984e-20, -2.569961e-21, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, 0, -1.798972e-20, -5.139921e-21, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, -1.541976e-20, -1.003089e-36, 
    2.569961e-21, -7.709882e-21, 0, -7.709882e-21, 7.709882e-21, 
    -7.709882e-21, 1.28498e-20, -5.139921e-21, 7.709882e-21, -5.139921e-21, 
    1.798972e-20, 1.003089e-36, -2.569961e-21, 1.28498e-20, -1.541976e-20, 
    2.569961e-21, 7.709882e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, -1.027984e-20, 2.569961e-21, -2.569961e-21, 
    1.28498e-20, 2.569961e-21, -5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -7.709882e-21, 0, -1.28498e-20, 5.139921e-21, -5.139921e-21, 0, 
    -2.569961e-21, 5.139921e-21, 1.28498e-20, 2.312965e-20, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, -2.055969e-20, 2.569961e-20, -5.139921e-21, 7.709882e-21, 
    1.027984e-20, 1.541976e-20, 1.027984e-20, -1.798972e-20, 1.798972e-20, 
    -1.541976e-20, -1.541976e-20, 2.312965e-20, -5.139921e-21, 2.312965e-20, 
    -2.826957e-20, 3.009266e-36, 1.798972e-20, -1.28498e-20, -7.709882e-21, 
    -1.003089e-36, -2.569961e-21, 5.139921e-21, -5.139921e-21, 1.027984e-20, 
    1.798972e-20, -3.083953e-20, -1.541976e-20, 7.709882e-21, -1.003089e-36, 
    -2.569961e-21, -1.28498e-20, 5.139921e-21, 1.027984e-20, -7.709882e-21, 
    -1.541976e-20, 1.027984e-20, -2.312965e-20, -1.28498e-20, -1.027984e-20, 
    -1.003089e-36, -1.798972e-20, 1.027984e-20, 2.569961e-20, -5.139921e-21, 
    2.312965e-20, 1.798972e-20, 2.569961e-21, 5.139921e-21, 0, 0, 
    -5.139921e-21, 0, -1.027984e-20, 7.709882e-21, -1.541976e-20, 
    -5.139921e-21, 7.709882e-21, 1.027984e-20, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, -2.312965e-20, 1.027984e-20, -1.798972e-20, 
    -2.055969e-20, -1.027984e-20, -2.055969e-20, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, -1.027984e-20, 1.28498e-20, -2.569961e-21, 
    -2.569961e-20, 5.139921e-21, 0, -7.709882e-21, -1.027984e-20, 
    1.541976e-20, -7.709882e-21, 1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 1.541976e-20, 
    1.027984e-20, 2.569961e-21, 2.312965e-20, 2.055969e-20, 1.027984e-20, 
    -1.28498e-20, -1.798972e-20, 1.28498e-20, -2.569961e-21, 1.541976e-20, 
    1.28498e-20, 1.027984e-20, -1.541976e-20, 7.709882e-21, -5.139921e-21, 
    1.003089e-36, 7.709882e-21, -2.569961e-21, 0, -7.709882e-21, 
    2.312965e-20, 1.027984e-20, 2.569961e-21, -2.312965e-20, -1.027984e-20, 
    7.709882e-21, 1.003089e-36, 1.541976e-20, 7.709882e-21, -1.541976e-20, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, -7.709882e-21, 0, 
    -5.139921e-21, 2.055969e-20, -5.139921e-21, -1.28498e-20, -2.569961e-21, 
    -2.312965e-20, 7.709882e-21, 0, 2.569961e-21, -5.139921e-21, 
    -1.541976e-20, -1.027984e-20, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    1.28498e-20, 1.027984e-20, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.541976e-20, -5.139921e-21, 1.541976e-20, 7.709882e-21, 
    -7.709882e-21, 2.569961e-21, -1.003089e-36, 7.709882e-21, -5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -7.709882e-21, 1.003089e-36, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 2.569961e-21, 1.798972e-20, 5.139921e-21, 
    -1.003089e-36, 7.709882e-21, 1.541976e-20, 1.003089e-36, -7.709882e-21, 
    1.28498e-20, -1.28498e-20, 7.709882e-21, 2.569961e-21, -1.28498e-20, 
    7.709882e-21, 2.569961e-21, 7.709882e-21, 7.709882e-21, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 0, 7.709882e-21, 7.709882e-21, -5.139921e-21, 
    2.569961e-20, -5.139921e-21, 1.28498e-20, 5.139921e-21, -2.055969e-20, 0, 
    1.28498e-20,
  6.259414e-29, 6.25942e-29, 6.259419e-29, 6.259425e-29, 6.259422e-29, 
    6.259425e-29, 6.259416e-29, 6.259421e-29, 6.259417e-29, 6.259415e-29, 
    6.259434e-29, 6.259425e-29, 6.259444e-29, 6.259438e-29, 6.259454e-29, 
    6.259443e-29, 6.259456e-29, 6.259453e-29, 6.259461e-29, 6.259459e-29, 
    6.259468e-29, 6.259462e-29, 6.259473e-29, 6.259467e-29, 6.259467e-29, 
    6.259461e-29, 6.259426e-29, 6.259433e-29, 6.259426e-29, 6.259427e-29, 
    6.259427e-29, 6.259422e-29, 6.259419e-29, 6.259414e-29, 6.259414e-29, 
    6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259432e-29, 6.259432e-29, 
    6.259441e-29, 6.259437e-29, 6.259451e-29, 6.259447e-29, 6.259459e-29, 
    6.259456e-29, 6.259459e-29, 6.259458e-29, 6.259459e-29, 6.259454e-29, 
    6.259456e-29, 6.259452e-29, 6.259437e-29, 6.259442e-29, 6.259429e-29, 
    6.259421e-29, 6.259416e-29, 6.259412e-29, 6.259413e-29, 6.259414e-29, 
    6.259419e-29, 6.259423e-29, 6.259427e-29, 6.259429e-29, 6.259432e-29, 
    6.259439e-29, 6.259443e-29, 6.259452e-29, 6.25945e-29, 6.259453e-29, 
    6.259455e-29, 6.25946e-29, 6.259459e-29, 6.259461e-29, 6.259453e-29, 
    6.259458e-29, 6.259449e-29, 6.259452e-29, 6.259432e-29, 6.259425e-29, 
    6.259422e-29, 6.25942e-29, 6.259413e-29, 6.259417e-29, 6.259416e-29, 
    6.25942e-29, 6.259423e-29, 6.259422e-29, 6.259429e-29, 6.259426e-29, 
    6.259443e-29, 6.259436e-29, 6.259455e-29, 6.25945e-29, 6.259456e-29, 
    6.259453e-29, 6.259458e-29, 6.259454e-29, 6.259462e-29, 6.259463e-29, 
    6.259463e-29, 6.259467e-29, 6.259453e-29, 6.259459e-29, 6.259422e-29, 
    6.259422e-29, 6.259423e-29, 6.259418e-29, 6.259418e-29, 6.259414e-29, 
    6.259417e-29, 6.259419e-29, 6.259423e-29, 6.259425e-29, 6.259428e-29, 
    6.259432e-29, 6.259438e-29, 6.259446e-29, 6.259451e-29, 6.259455e-29, 
    6.259452e-29, 6.259455e-29, 6.259452e-29, 6.259451e-29, 6.259463e-29, 
    6.259456e-29, 6.259466e-29, 6.259466e-29, 6.259461e-29, 6.259466e-29, 
    6.259422e-29, 6.25942e-29, 6.259416e-29, 6.259419e-29, 6.259413e-29, 
    6.259417e-29, 6.259419e-29, 6.259426e-29, 6.259428e-29, 6.25943e-29, 
    6.259433e-29, 6.259437e-29, 6.259444e-29, 6.25945e-29, 6.259456e-29, 
    6.259455e-29, 6.259455e-29, 6.259456e-29, 6.259453e-29, 6.259457e-29, 
    6.259458e-29, 6.259456e-29, 6.259466e-29, 6.259463e-29, 6.259466e-29, 
    6.259464e-29, 6.259421e-29, 6.259423e-29, 6.259422e-29, 6.259424e-29, 
    6.259422e-29, 6.259429e-29, 6.259431e-29, 6.259441e-29, 6.259437e-29, 
    6.259443e-29, 6.259437e-29, 6.259438e-29, 6.259443e-29, 6.259438e-29, 
    6.25945e-29, 6.259441e-29, 6.259456e-29, 6.259449e-29, 6.259457e-29, 
    6.259456e-29, 6.259458e-29, 6.259461e-29, 6.259464e-29, 6.259469e-29, 
    6.259468e-29, 6.259472e-29, 6.259426e-29, 6.259429e-29, 6.259429e-29, 
    6.259432e-29, 6.259434e-29, 6.259438e-29, 6.259446e-29, 6.259443e-29, 
    6.259448e-29, 6.259449e-29, 6.259441e-29, 6.259446e-29, 6.259431e-29, 
    6.259433e-29, 6.259432e-29, 6.259426e-29, 6.259444e-29, 6.259435e-29, 
    6.259451e-29, 6.259446e-29, 6.25946e-29, 6.259453e-29, 6.259467e-29, 
    6.259473e-29, 6.259478e-29, 6.259485e-29, 6.259431e-29, 6.259428e-29, 
    6.259432e-29, 6.259437e-29, 6.259441e-29, 6.259446e-29, 6.259447e-29, 
    6.259448e-29, 6.259451e-29, 6.259453e-29, 6.259449e-29, 6.259454e-29, 
    6.259434e-29, 6.259444e-29, 6.259428e-29, 6.259433e-29, 6.259436e-29, 
    6.259435e-29, 6.259443e-29, 6.259444e-29, 6.259452e-29, 6.259448e-29, 
    6.259472e-29, 6.259461e-29, 6.25949e-29, 6.259482e-29, 6.259428e-29, 
    6.259431e-29, 6.259439e-29, 6.259435e-29, 6.259447e-29, 6.25945e-29, 
    6.259452e-29, 6.259455e-29, 6.259456e-29, 6.259458e-29, 6.259455e-29, 
    6.259457e-29, 6.259447e-29, 6.259452e-29, 6.259438e-29, 6.259441e-29, 
    6.25944e-29, 6.259438e-29, 6.259443e-29, 6.259449e-29, 6.259449e-29, 
    6.25945e-29, 6.259455e-29, 6.259447e-29, 6.259473e-29, 6.259457e-29, 
    6.259433e-29, 6.259438e-29, 6.259438e-29, 6.259437e-29, 6.25945e-29, 
    6.259445e-29, 6.259458e-29, 6.259454e-29, 6.259459e-29, 6.259457e-29, 
    6.259456e-29, 6.259453e-29, 6.25945e-29, 6.259445e-29, 6.259441e-29, 
    6.259437e-29, 6.259438e-29, 6.259442e-29, 6.259449e-29, 6.259456e-29, 
    6.259454e-29, 6.259459e-29, 6.259446e-29, 6.259452e-29, 6.259449e-29, 
    6.259455e-29, 6.259443e-29, 6.259453e-29, 6.25944e-29, 6.259441e-29, 
    6.259445e-29, 6.259452e-29, 6.259453e-29, 6.259455e-29, 6.259454e-29, 
    6.259449e-29, 6.259448e-29, 6.259445e-29, 6.259444e-29, 6.259441e-29, 
    6.259439e-29, 6.259441e-29, 6.259443e-29, 6.259449e-29, 6.259455e-29, 
    6.259461e-29, 6.259462e-29, 6.259469e-29, 6.259463e-29, 6.259473e-29, 
    6.259465e-29, 6.259479e-29, 6.259453e-29, 6.259464e-29, 6.259445e-29, 
    6.259447e-29, 6.259451e-29, 6.259459e-29, 6.259455e-29, 6.259461e-29, 
    6.259448e-29, 6.259442e-29, 6.25944e-29, 6.259437e-29, 6.25944e-29, 
    6.25944e-29, 6.259443e-29, 6.259442e-29, 6.259449e-29, 6.259446e-29, 
    6.259456e-29, 6.259461e-29, 6.259472e-29, 6.259479e-29, 6.259486e-29, 
    6.259489e-29, 6.25949e-29, 6.25949e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.19478e-10, 2.204436e-10, 2.202559e-10, 2.210348e-10, 2.206027e-10, 
    2.211127e-10, 2.196738e-10, 2.20482e-10, 2.19966e-10, 2.195649e-10, 
    2.225463e-10, 2.210695e-10, 2.240801e-10, 2.231383e-10, 2.255041e-10, 
    2.239336e-10, 2.258208e-10, 2.254587e-10, 2.265482e-10, 2.262361e-10, 
    2.276297e-10, 2.266923e-10, 2.28352e-10, 2.274058e-10, 2.275538e-10, 
    2.266613e-10, 2.213667e-10, 2.223624e-10, 2.213077e-10, 2.214497e-10, 
    2.21386e-10, 2.206117e-10, 2.202215e-10, 2.194042e-10, 2.195526e-10, 
    2.201528e-10, 2.215135e-10, 2.210516e-10, 2.222157e-10, 2.221894e-10, 
    2.234854e-10, 2.229011e-10, 2.250793e-10, 2.244602e-10, 2.262491e-10, 
    2.257992e-10, 2.26228e-10, 2.26098e-10, 2.262297e-10, 2.255699e-10, 
    2.258526e-10, 2.252719e-10, 2.230105e-10, 2.236751e-10, 2.216929e-10, 
    2.20501e-10, 2.197092e-10, 2.191474e-10, 2.192268e-10, 2.193783e-10, 
    2.201563e-10, 2.208878e-10, 2.214453e-10, 2.218182e-10, 2.221856e-10, 
    2.232979e-10, 2.238865e-10, 2.252045e-10, 2.249666e-10, 2.253695e-10, 
    2.257545e-10, 2.264008e-10, 2.262944e-10, 2.265791e-10, 2.253589e-10, 
    2.261699e-10, 2.248311e-10, 2.251973e-10, 2.222856e-10, 2.211762e-10, 
    2.207048e-10, 2.20292e-10, 2.192879e-10, 2.199813e-10, 2.19708e-10, 
    2.203583e-10, 2.207715e-10, 2.205671e-10, 2.218284e-10, 2.213381e-10, 
    2.239214e-10, 2.228086e-10, 2.257096e-10, 2.250154e-10, 2.25876e-10, 
    2.254368e-10, 2.261892e-10, 2.255121e-10, 2.266851e-10, 2.269405e-10, 
    2.26766e-10, 2.274365e-10, 2.254745e-10, 2.26228e-10, 2.205614e-10, 
    2.205947e-10, 2.2075e-10, 2.200674e-10, 2.200257e-10, 2.194001e-10, 
    2.199567e-10, 2.201938e-10, 2.207954e-10, 2.211513e-10, 2.214896e-10, 
    2.222335e-10, 2.230642e-10, 2.242259e-10, 2.250604e-10, 2.256198e-10, 
    2.252768e-10, 2.255796e-10, 2.252411e-10, 2.250824e-10, 2.268448e-10, 
    2.258552e-10, 2.2734e-10, 2.272579e-10, 2.265859e-10, 2.272671e-10, 
    2.206181e-10, 2.204263e-10, 2.197604e-10, 2.202815e-10, 2.19332e-10, 
    2.198635e-10, 2.201691e-10, 2.213483e-10, 2.216074e-10, 2.218476e-10, 
    2.223221e-10, 2.22931e-10, 2.239991e-10, 2.249285e-10, 2.257769e-10, 
    2.257147e-10, 2.257366e-10, 2.259261e-10, 2.254566e-10, 2.260032e-10, 
    2.260949e-10, 2.258551e-10, 2.272469e-10, 2.268492e-10, 2.272561e-10, 
    2.269972e-10, 2.204887e-10, 2.208114e-10, 2.20637e-10, 2.20965e-10, 
    2.207339e-10, 2.217613e-10, 2.220693e-10, 2.235105e-10, 2.22919e-10, 
    2.238603e-10, 2.230146e-10, 2.231645e-10, 2.238911e-10, 2.230603e-10, 
    2.248773e-10, 2.236455e-10, 2.259335e-10, 2.247035e-10, 2.260106e-10, 
    2.257732e-10, 2.261662e-10, 2.265182e-10, 2.26961e-10, 2.277781e-10, 
    2.275889e-10, 2.282721e-10, 2.212925e-10, 2.217112e-10, 2.216743e-10, 
    2.221124e-10, 2.224363e-10, 2.231385e-10, 2.242648e-10, 2.238413e-10, 
    2.246187e-10, 2.247748e-10, 2.235936e-10, 2.243189e-10, 2.219913e-10, 
    2.223674e-10, 2.221435e-10, 2.213256e-10, 2.239389e-10, 2.225977e-10, 
    2.250742e-10, 2.243477e-10, 2.26468e-10, 2.254135e-10, 2.274847e-10, 
    2.283702e-10, 2.292034e-10, 2.301773e-10, 2.219396e-10, 2.216552e-10, 
    2.221645e-10, 2.228691e-10, 2.235228e-10, 2.24392e-10, 2.244809e-10, 
    2.246437e-10, 2.250655e-10, 2.254201e-10, 2.246952e-10, 2.25509e-10, 
    2.224547e-10, 2.240553e-10, 2.215476e-10, 2.223028e-10, 2.228276e-10, 
    2.225973e-10, 2.237928e-10, 2.240746e-10, 2.252196e-10, 2.246277e-10, 
    2.281516e-10, 2.265926e-10, 2.309187e-10, 2.297098e-10, 2.215558e-10, 
    2.219386e-10, 2.23271e-10, 2.226371e-10, 2.2445e-10, 2.248963e-10, 
    2.25259e-10, 2.257227e-10, 2.257728e-10, 2.260476e-10, 2.255973e-10, 
    2.260298e-10, 2.243938e-10, 2.251249e-10, 2.231187e-10, 2.23607e-10, 
    2.233824e-10, 2.23136e-10, 2.238964e-10, 2.247067e-10, 2.247239e-10, 
    2.249837e-10, 2.257159e-10, 2.244573e-10, 2.283529e-10, 2.259472e-10, 
    2.223561e-10, 2.230935e-10, 2.231988e-10, 2.229131e-10, 2.248515e-10, 
    2.241492e-10, 2.260409e-10, 2.255296e-10, 2.263673e-10, 2.25951e-10, 
    2.258898e-10, 2.253552e-10, 2.250223e-10, 2.241814e-10, 2.234972e-10, 
    2.229546e-10, 2.230807e-10, 2.236768e-10, 2.247562e-10, 2.257774e-10, 
    2.255537e-10, 2.263036e-10, 2.243185e-10, 2.251509e-10, 2.248292e-10, 
    2.256681e-10, 2.2383e-10, 2.253953e-10, 2.234299e-10, 2.236022e-10, 
    2.241352e-10, 2.252074e-10, 2.254446e-10, 2.256979e-10, 2.255416e-10, 
    2.247836e-10, 2.246594e-10, 2.241223e-10, 2.23974e-10, 2.235647e-10, 
    2.232259e-10, 2.235355e-10, 2.238606e-10, 2.247839e-10, 2.25616e-10, 
    2.265232e-10, 2.267452e-10, 2.278052e-10, 2.269424e-10, 2.283663e-10, 
    2.271558e-10, 2.292513e-10, 2.25486e-10, 2.271201e-10, 2.241595e-10, 
    2.244784e-10, 2.250553e-10, 2.263785e-10, 2.256641e-10, 2.264996e-10, 
    2.246545e-10, 2.236973e-10, 2.234496e-10, 2.229876e-10, 2.234602e-10, 
    2.234218e-10, 2.23874e-10, 2.237287e-10, 2.248146e-10, 2.242313e-10, 
    2.258883e-10, 2.264929e-10, 2.282005e-10, 2.292474e-10, 2.303129e-10, 
    2.307833e-10, 2.309265e-10, 2.309864e-10 ;

 SOIL2N_TO_SOIL3N =
  1.5677e-11, 1.574598e-11, 1.573257e-11, 1.57882e-11, 1.575734e-11, 
    1.579377e-11, 1.569098e-11, 1.574871e-11, 1.571186e-11, 1.568321e-11, 
    1.589616e-11, 1.579068e-11, 1.600572e-11, 1.593845e-11, 1.610743e-11, 
    1.599525e-11, 1.613005e-11, 1.61042e-11, 1.618202e-11, 1.615972e-11, 
    1.625926e-11, 1.61923e-11, 1.631086e-11, 1.624327e-11, 1.625384e-11, 
    1.61901e-11, 1.581191e-11, 1.588303e-11, 1.580769e-11, 1.581783e-11, 
    1.581328e-11, 1.575797e-11, 1.57301e-11, 1.567173e-11, 1.568233e-11, 
    1.57252e-11, 1.58224e-11, 1.57894e-11, 1.587255e-11, 1.587067e-11, 
    1.596324e-11, 1.59215e-11, 1.607709e-11, 1.603287e-11, 1.616065e-11, 
    1.612852e-11, 1.615914e-11, 1.614986e-11, 1.615926e-11, 1.611213e-11, 
    1.613233e-11, 1.609085e-11, 1.592932e-11, 1.59768e-11, 1.58352e-11, 
    1.575007e-11, 1.569352e-11, 1.565339e-11, 1.565906e-11, 1.566988e-11, 
    1.572545e-11, 1.57777e-11, 1.581752e-11, 1.584416e-11, 1.58704e-11, 
    1.594985e-11, 1.599189e-11, 1.608603e-11, 1.606904e-11, 1.609782e-11, 
    1.612532e-11, 1.617148e-11, 1.616388e-11, 1.618422e-11, 1.609706e-11, 
    1.615499e-11, 1.605936e-11, 1.608552e-11, 1.587754e-11, 1.57983e-11, 
    1.576463e-11, 1.573514e-11, 1.566342e-11, 1.571295e-11, 1.569343e-11, 
    1.573988e-11, 1.576939e-11, 1.575479e-11, 1.584489e-11, 1.580986e-11, 
    1.599438e-11, 1.59149e-11, 1.612211e-11, 1.607253e-11, 1.6134e-11, 
    1.610263e-11, 1.615637e-11, 1.610801e-11, 1.619179e-11, 1.621004e-11, 
    1.619757e-11, 1.624546e-11, 1.610532e-11, 1.615914e-11, 1.575439e-11, 
    1.575677e-11, 1.576786e-11, 1.57191e-11, 1.571612e-11, 1.567144e-11, 
    1.571119e-11, 1.572813e-11, 1.57711e-11, 1.579652e-11, 1.582069e-11, 
    1.587382e-11, 1.593316e-11, 1.601613e-11, 1.607574e-11, 1.61157e-11, 
    1.60912e-11, 1.611283e-11, 1.608865e-11, 1.607731e-11, 1.62032e-11, 
    1.613252e-11, 1.623857e-11, 1.62327e-11, 1.618471e-11, 1.623337e-11, 
    1.575844e-11, 1.574474e-11, 1.569717e-11, 1.573439e-11, 1.566657e-11, 
    1.570454e-11, 1.572637e-11, 1.581059e-11, 1.58291e-11, 1.584626e-11, 
    1.588015e-11, 1.592364e-11, 1.599994e-11, 1.606632e-11, 1.612692e-11, 
    1.612248e-11, 1.612404e-11, 1.613758e-11, 1.610405e-11, 1.614309e-11, 
    1.614964e-11, 1.613251e-11, 1.623192e-11, 1.620352e-11, 1.623258e-11, 
    1.621409e-11, 1.574919e-11, 1.577224e-11, 1.575979e-11, 1.578321e-11, 
    1.576671e-11, 1.584009e-11, 1.586209e-11, 1.596503e-11, 1.592279e-11, 
    1.599003e-11, 1.592962e-11, 1.594032e-11, 1.599222e-11, 1.593288e-11, 
    1.606266e-11, 1.597468e-11, 1.613811e-11, 1.605025e-11, 1.614361e-11, 
    1.612666e-11, 1.615473e-11, 1.617987e-11, 1.62115e-11, 1.626986e-11, 
    1.625635e-11, 1.630515e-11, 1.580661e-11, 1.583651e-11, 1.583388e-11, 
    1.586517e-11, 1.588831e-11, 1.593847e-11, 1.601891e-11, 1.598866e-11, 
    1.60442e-11, 1.605534e-11, 1.597097e-11, 1.602278e-11, 1.585652e-11, 
    1.588338e-11, 1.586739e-11, 1.580897e-11, 1.599563e-11, 1.589984e-11, 
    1.607673e-11, 1.602483e-11, 1.617629e-11, 1.610097e-11, 1.624891e-11, 
    1.631215e-11, 1.637167e-11, 1.644123e-11, 1.585283e-11, 1.583251e-11, 
    1.586889e-11, 1.591922e-11, 1.596592e-11, 1.6028e-11, 1.603435e-11, 
    1.604598e-11, 1.607611e-11, 1.610144e-11, 1.604966e-11, 1.610779e-11, 
    1.588962e-11, 1.600395e-11, 1.582483e-11, 1.587877e-11, 1.591625e-11, 
    1.589981e-11, 1.59852e-11, 1.600533e-11, 1.608712e-11, 1.604484e-11, 
    1.629655e-11, 1.618518e-11, 1.649419e-11, 1.640784e-11, 1.582541e-11, 
    1.585276e-11, 1.594793e-11, 1.590265e-11, 1.603214e-11, 1.606402e-11, 
    1.608993e-11, 1.612305e-11, 1.612663e-11, 1.614625e-11, 1.611409e-11, 
    1.614498e-11, 1.602813e-11, 1.608035e-11, 1.593705e-11, 1.597193e-11, 
    1.595588e-11, 1.593828e-11, 1.59926e-11, 1.605048e-11, 1.605171e-11, 
    1.607027e-11, 1.612257e-11, 1.603267e-11, 1.631092e-11, 1.613908e-11, 
    1.588258e-11, 1.593525e-11, 1.594277e-11, 1.592237e-11, 1.606082e-11, 
    1.601066e-11, 1.614578e-11, 1.610926e-11, 1.616909e-11, 1.613936e-11, 
    1.613499e-11, 1.60968e-11, 1.607302e-11, 1.601296e-11, 1.596408e-11, 
    1.592533e-11, 1.593434e-11, 1.597691e-11, 1.605401e-11, 1.612695e-11, 
    1.611098e-11, 1.616455e-11, 1.602275e-11, 1.608221e-11, 1.605923e-11, 
    1.611915e-11, 1.598786e-11, 1.609967e-11, 1.595928e-11, 1.597159e-11, 
    1.600966e-11, 1.608625e-11, 1.610318e-11, 1.612128e-11, 1.611011e-11, 
    1.605597e-11, 1.60471e-11, 1.600873e-11, 1.599814e-11, 1.596891e-11, 
    1.59447e-11, 1.596682e-11, 1.599004e-11, 1.605599e-11, 1.611543e-11, 
    1.618023e-11, 1.619609e-11, 1.62718e-11, 1.621017e-11, 1.631188e-11, 
    1.622541e-11, 1.637509e-11, 1.610614e-11, 1.622286e-11, 1.601139e-11, 
    1.603417e-11, 1.607538e-11, 1.616989e-11, 1.611887e-11, 1.617854e-11, 
    1.604675e-11, 1.597838e-11, 1.596069e-11, 1.592768e-11, 1.596144e-11, 
    1.59587e-11, 1.5991e-11, 1.598062e-11, 1.605818e-11, 1.601652e-11, 
    1.613488e-11, 1.617807e-11, 1.630004e-11, 1.637481e-11, 1.645092e-11, 
    1.648452e-11, 1.649475e-11, 1.649903e-11 ;

 SOIL2N_vr =
  1.818768, 1.81877, 1.818769, 1.818771, 1.81877, 1.818771, 1.818769, 
    1.81877, 1.818769, 1.818768, 1.818773, 1.818771, 1.818775, 1.818774, 
    1.818778, 1.818775, 1.818778, 1.818778, 1.818779, 1.818779, 1.818781, 
    1.81878, 1.818782, 1.818781, 1.818781, 1.818779, 1.818771, 1.818773, 
    1.818771, 1.818771, 1.818771, 1.81877, 1.818769, 1.818768, 1.818768, 
    1.818769, 1.818771, 1.818771, 1.818772, 1.818772, 1.818774, 1.818774, 
    1.818777, 1.818776, 1.818779, 1.818778, 1.818779, 1.818779, 1.818779, 
    1.818778, 1.818778, 1.818777, 1.818774, 1.818775, 1.818772, 1.81877, 
    1.818769, 1.818768, 1.818768, 1.818768, 1.818769, 1.81877, 1.818771, 
    1.818772, 1.818772, 1.818774, 1.818775, 1.818777, 1.818777, 1.818777, 
    1.818778, 1.818779, 1.818779, 1.818779, 1.818777, 1.818779, 1.818777, 
    1.818777, 1.818773, 1.818771, 1.81877, 1.818769, 1.818768, 1.818769, 
    1.818769, 1.81877, 1.81877, 1.81877, 1.818772, 1.818771, 1.818775, 
    1.818773, 1.818778, 1.818777, 1.818778, 1.818778, 1.818779, 1.818778, 
    1.818779, 1.81878, 1.81878, 1.818781, 1.818778, 1.818779, 1.81877, 
    1.81877, 1.81877, 1.818769, 1.818769, 1.818768, 1.818769, 1.818769, 
    1.81877, 1.818771, 1.818771, 1.818773, 1.818774, 1.818776, 1.818777, 
    1.818778, 1.818777, 1.818778, 1.818777, 1.818777, 1.81878, 1.818778, 
    1.818781, 1.81878, 1.818779, 1.81878, 1.81877, 1.81877, 1.818769, 
    1.818769, 1.818768, 1.818769, 1.818769, 1.818771, 1.818771, 1.818772, 
    1.818773, 1.818774, 1.818775, 1.818777, 1.818778, 1.818778, 1.818778, 
    1.818778, 1.818778, 1.818778, 1.818779, 1.818778, 1.81878, 1.81878, 
    1.81878, 1.81878, 1.81877, 1.81877, 1.81877, 1.818771, 1.81877, 1.818772, 
    1.818772, 1.818775, 1.818774, 1.818775, 1.818774, 1.818774, 1.818775, 
    1.818774, 1.818777, 1.818775, 1.818778, 1.818776, 1.818779, 1.818778, 
    1.818779, 1.818779, 1.81878, 1.818781, 1.818781, 1.818782, 1.818771, 
    1.818772, 1.818772, 1.818772, 1.818773, 1.818774, 1.818776, 1.818775, 
    1.818776, 1.818776, 1.818775, 1.818776, 1.818772, 1.818773, 1.818772, 
    1.818771, 1.818775, 1.818773, 1.818777, 1.818776, 1.818779, 1.818778, 
    1.818781, 1.818782, 1.818784, 1.818785, 1.818772, 1.818772, 1.818772, 
    1.818774, 1.818775, 1.818776, 1.818776, 1.818776, 1.818777, 1.818778, 
    1.818776, 1.818778, 1.818773, 1.818775, 1.818771, 1.818773, 1.818773, 
    1.818773, 1.818775, 1.818775, 1.818777, 1.818776, 1.818782, 1.818779, 
    1.818786, 1.818784, 1.818771, 1.818772, 1.818774, 1.818773, 1.818776, 
    1.818777, 1.818777, 1.818778, 1.818778, 1.818779, 1.818778, 1.818779, 
    1.818776, 1.818777, 1.818774, 1.818775, 1.818774, 1.818774, 1.818775, 
    1.818776, 1.818776, 1.818777, 1.818778, 1.818776, 1.818782, 1.818778, 
    1.818773, 1.818774, 1.818774, 1.818774, 1.818777, 1.818776, 1.818779, 
    1.818778, 1.818779, 1.818778, 1.818778, 1.818777, 1.818777, 1.818776, 
    1.818774, 1.818774, 1.818774, 1.818775, 1.818776, 1.818778, 1.818778, 
    1.818779, 1.818776, 1.818777, 1.818777, 1.818778, 1.818775, 1.818777, 
    1.818774, 1.818775, 1.818776, 1.818777, 1.818778, 1.818778, 1.818778, 
    1.818776, 1.818776, 1.818776, 1.818775, 1.818775, 1.818774, 1.818775, 
    1.818775, 1.818776, 1.818778, 1.818779, 1.81878, 1.818781, 1.81878, 
    1.818782, 1.81878, 1.818784, 1.818778, 1.81878, 1.818776, 1.818776, 
    1.818777, 1.818779, 1.818778, 1.818779, 1.818776, 1.818775, 1.818774, 
    1.818774, 1.818774, 1.818774, 1.818775, 1.818775, 1.818777, 1.818776, 
    1.818778, 1.818779, 1.818782, 1.818784, 1.818785, 1.818786, 1.818786, 
    1.818786,
  1.818734, 1.818736, 1.818735, 1.818737, 1.818736, 1.818737, 1.818734, 
    1.818736, 1.818735, 1.818734, 1.81874, 1.818737, 1.818744, 1.818742, 
    1.818747, 1.818743, 1.818747, 1.818747, 1.818749, 1.818748, 1.818751, 
    1.818749, 1.818753, 1.818751, 1.818751, 1.818749, 1.818738, 1.81874, 
    1.818738, 1.818738, 1.818738, 1.818736, 1.818735, 1.818734, 1.818734, 
    1.818735, 1.818738, 1.818737, 1.81874, 1.81874, 1.818742, 1.818741, 
    1.818746, 1.818745, 1.818748, 1.818747, 1.818748, 1.818748, 1.818748, 
    1.818747, 1.818747, 1.818746, 1.818741, 1.818743, 1.818739, 1.818736, 
    1.818734, 1.818733, 1.818733, 1.818734, 1.818735, 1.818737, 1.818738, 
    1.818739, 1.81874, 1.818742, 1.818743, 1.818746, 1.818746, 1.818746, 
    1.818747, 1.818749, 1.818748, 1.818749, 1.818746, 1.818748, 1.818745, 
    1.818746, 1.81874, 1.818738, 1.818736, 1.818736, 1.818733, 1.818735, 
    1.818734, 1.818736, 1.818737, 1.818736, 1.818739, 1.818738, 1.818743, 
    1.818741, 1.818747, 1.818746, 1.818748, 1.818747, 1.818748, 1.818747, 
    1.818749, 1.81875, 1.818749, 1.818751, 1.818747, 1.818748, 1.818736, 
    1.818736, 1.818737, 1.818735, 1.818735, 1.818734, 1.818735, 1.818735, 
    1.818737, 1.818737, 1.818738, 1.81874, 1.818742, 1.818744, 1.818746, 
    1.818747, 1.818746, 1.818747, 1.818746, 1.818746, 1.81875, 1.818747, 
    1.818751, 1.81875, 1.818749, 1.818751, 1.818736, 1.818736, 1.818735, 
    1.818736, 1.818734, 1.818735, 1.818735, 1.818738, 1.818738, 1.818739, 
    1.81874, 1.818741, 1.818743, 1.818745, 1.818747, 1.818747, 1.818747, 
    1.818748, 1.818747, 1.818748, 1.818748, 1.818747, 1.81875, 1.81875, 
    1.81875, 1.81875, 1.818736, 1.818737, 1.818736, 1.818737, 1.818737, 
    1.818739, 1.818739, 1.818743, 1.818741, 1.818743, 1.818741, 1.818742, 
    1.818743, 1.818742, 1.818745, 1.818743, 1.818748, 1.818745, 1.818748, 
    1.818747, 1.818748, 1.818749, 1.81875, 1.818752, 1.818751, 1.818753, 
    1.818738, 1.818739, 1.818739, 1.81874, 1.81874, 1.818742, 1.818744, 
    1.818743, 1.818745, 1.818745, 1.818743, 1.818744, 1.818739, 1.81874, 
    1.81874, 1.818738, 1.818743, 1.81874, 1.818746, 1.818744, 1.818749, 
    1.818747, 1.818751, 1.818753, 1.818755, 1.818757, 1.818739, 1.818738, 
    1.81874, 1.818741, 1.818743, 1.818744, 1.818745, 1.818745, 1.818746, 
    1.818747, 1.818745, 1.818747, 1.81874, 1.818744, 1.818738, 1.81874, 
    1.818741, 1.81874, 1.818743, 1.818744, 1.818746, 1.818745, 1.818752, 
    1.818749, 1.818758, 1.818756, 1.818738, 1.818739, 1.818742, 1.818741, 
    1.818744, 1.818745, 1.818746, 1.818747, 1.818747, 1.818748, 1.818747, 
    1.818748, 1.818744, 1.818746, 1.818742, 1.818743, 1.818742, 1.818742, 
    1.818743, 1.818745, 1.818745, 1.818746, 1.818747, 1.818745, 1.818753, 
    1.818748, 1.81874, 1.818742, 1.818742, 1.818741, 1.818745, 1.818744, 
    1.818748, 1.818747, 1.818749, 1.818748, 1.818748, 1.818746, 1.818746, 
    1.818744, 1.818742, 1.818741, 1.818742, 1.818743, 1.818745, 1.818747, 
    1.818747, 1.818748, 1.818744, 1.818746, 1.818745, 1.818747, 1.818743, 
    1.818746, 1.818742, 1.818743, 1.818744, 1.818746, 1.818747, 1.818747, 
    1.818747, 1.818745, 1.818745, 1.818744, 1.818743, 1.818743, 1.818742, 
    1.818743, 1.818743, 1.818745, 1.818747, 1.818749, 1.818749, 1.818752, 
    1.81875, 1.818753, 1.81875, 1.818755, 1.818747, 1.81875, 1.818744, 
    1.818745, 1.818746, 1.818749, 1.818747, 1.818749, 1.818745, 1.818743, 
    1.818742, 1.818741, 1.818742, 1.818742, 1.818743, 1.818743, 1.818745, 
    1.818744, 1.818748, 1.818749, 1.818752, 1.818755, 1.818757, 1.818758, 
    1.818758, 1.818758,
  1.818684, 1.818686, 1.818686, 1.818687, 1.818686, 1.818687, 1.818684, 
    1.818686, 1.818685, 1.818684, 1.818691, 1.818687, 1.818694, 1.818692, 
    1.818697, 1.818694, 1.818698, 1.818697, 1.8187, 1.818699, 1.818702, 
    1.8187, 1.818704, 1.818702, 1.818702, 1.8187, 1.818688, 1.81869, 
    1.818688, 1.818688, 1.818688, 1.818686, 1.818685, 1.818684, 1.818684, 
    1.818685, 1.818688, 1.818687, 1.81869, 1.81869, 1.818693, 1.818691, 
    1.818696, 1.818695, 1.818699, 1.818698, 1.818699, 1.818699, 1.818699, 
    1.818698, 1.818698, 1.818697, 1.818692, 1.818693, 1.818689, 1.818686, 
    1.818684, 1.818683, 1.818683, 1.818684, 1.818685, 1.818687, 1.818688, 
    1.818689, 1.81869, 1.818692, 1.818694, 1.818697, 1.818696, 1.818697, 
    1.818698, 1.818699, 1.818699, 1.8187, 1.818697, 1.818699, 1.818696, 
    1.818697, 1.81869, 1.818688, 1.818686, 1.818686, 1.818683, 1.818685, 
    1.818684, 1.818686, 1.818687, 1.818686, 1.818689, 1.818688, 1.818694, 
    1.818691, 1.818698, 1.818696, 1.818698, 1.818697, 1.818699, 1.818697, 
    1.8187, 1.818701, 1.8187, 1.818702, 1.818697, 1.818699, 1.818686, 
    1.818686, 1.818687, 1.818685, 1.818685, 1.818684, 1.818685, 1.818685, 
    1.818687, 1.818688, 1.818688, 1.81869, 1.818692, 1.818695, 1.818696, 
    1.818698, 1.818697, 1.818698, 1.818697, 1.818696, 1.818701, 1.818698, 
    1.818702, 1.818701, 1.8187, 1.818702, 1.818686, 1.818686, 1.818684, 
    1.818686, 1.818683, 1.818685, 1.818685, 1.818688, 1.818689, 1.818689, 
    1.81869, 1.818692, 1.818694, 1.818696, 1.818698, 1.818698, 1.818698, 
    1.818698, 1.818697, 1.818699, 1.818699, 1.818698, 1.818701, 1.818701, 
    1.818701, 1.818701, 1.818686, 1.818687, 1.818686, 1.818687, 1.818687, 
    1.818689, 1.81869, 1.818693, 1.818692, 1.818694, 1.818692, 1.818692, 
    1.818694, 1.818692, 1.818696, 1.818693, 1.818698, 1.818696, 1.818699, 
    1.818698, 1.818699, 1.8187, 1.818701, 1.818703, 1.818702, 1.818704, 
    1.818688, 1.818689, 1.818689, 1.81869, 1.818691, 1.818692, 1.818695, 
    1.818694, 1.818695, 1.818696, 1.818693, 1.818695, 1.818689, 1.81869, 
    1.81869, 1.818688, 1.818694, 1.818691, 1.818696, 1.818695, 1.8187, 
    1.818697, 1.818702, 1.818704, 1.818706, 1.818708, 1.818689, 1.818689, 
    1.81869, 1.818691, 1.818693, 1.818695, 1.818695, 1.818696, 1.818696, 
    1.818697, 1.818696, 1.818697, 1.818691, 1.818694, 1.818689, 1.81869, 
    1.818691, 1.818691, 1.818694, 1.818694, 1.818697, 1.818695, 1.818703, 
    1.8187, 1.81871, 1.818707, 1.818689, 1.818689, 1.818692, 1.818691, 
    1.818695, 1.818696, 1.818697, 1.818698, 1.818698, 1.818699, 1.818698, 
    1.818699, 1.818695, 1.818697, 1.818692, 1.818693, 1.818693, 1.818692, 
    1.818694, 1.818696, 1.818696, 1.818696, 1.818698, 1.818695, 1.818704, 
    1.818698, 1.81869, 1.818692, 1.818692, 1.818692, 1.818696, 1.818694, 
    1.818699, 1.818698, 1.818699, 1.818699, 1.818698, 1.818697, 1.818696, 
    1.818694, 1.818693, 1.818692, 1.818692, 1.818693, 1.818696, 1.818698, 
    1.818698, 1.818699, 1.818695, 1.818697, 1.818696, 1.818698, 1.818694, 
    1.818697, 1.818693, 1.818693, 1.818694, 1.818697, 1.818697, 1.818698, 
    1.818698, 1.818696, 1.818696, 1.818694, 1.818694, 1.818693, 1.818692, 
    1.818693, 1.818694, 1.818696, 1.818698, 1.8187, 1.8187, 1.818703, 
    1.818701, 1.818704, 1.818701, 1.818706, 1.818697, 1.818701, 1.818694, 
    1.818695, 1.818696, 1.818699, 1.818698, 1.8187, 1.818696, 1.818693, 
    1.818693, 1.818692, 1.818693, 1.818693, 1.818694, 1.818693, 1.818696, 
    1.818695, 1.818698, 1.8187, 1.818704, 1.818706, 1.818708, 1.818709, 
    1.81871, 1.81871,
  1.818644, 1.818646, 1.818645, 1.818647, 1.818646, 1.818647, 1.818644, 
    1.818646, 1.818645, 1.818644, 1.818651, 1.818647, 1.818654, 1.818652, 
    1.818657, 1.818654, 1.818658, 1.818657, 1.81866, 1.818659, 1.818662, 
    1.81866, 1.818664, 1.818662, 1.818662, 1.81866, 1.818648, 1.81865, 
    1.818648, 1.818648, 1.818648, 1.818646, 1.818645, 1.818644, 1.818644, 
    1.818645, 1.818648, 1.818647, 1.81865, 1.81865, 1.818653, 1.818651, 
    1.818656, 1.818655, 1.818659, 1.818658, 1.818659, 1.818659, 1.818659, 
    1.818658, 1.818658, 1.818657, 1.818652, 1.818653, 1.818649, 1.818646, 
    1.818644, 1.818643, 1.818643, 1.818644, 1.818645, 1.818647, 1.818648, 
    1.818649, 1.81865, 1.818652, 1.818654, 1.818657, 1.818656, 1.818657, 
    1.818658, 1.818659, 1.818659, 1.81866, 1.818657, 1.818659, 1.818656, 
    1.818657, 1.81865, 1.818648, 1.818647, 1.818646, 1.818643, 1.818645, 
    1.818644, 1.818646, 1.818647, 1.818646, 1.818649, 1.818648, 1.818654, 
    1.818651, 1.818658, 1.818656, 1.818658, 1.818657, 1.818659, 1.818657, 
    1.81866, 1.818661, 1.81866, 1.818662, 1.818657, 1.818659, 1.818646, 
    1.818646, 1.818647, 1.818645, 1.818645, 1.818644, 1.818645, 1.818645, 
    1.818647, 1.818648, 1.818648, 1.81865, 1.818652, 1.818654, 1.818656, 
    1.818658, 1.818657, 1.818658, 1.818657, 1.818656, 1.81866, 1.818658, 
    1.818661, 1.818661, 1.81866, 1.818661, 1.818646, 1.818646, 1.818644, 
    1.818646, 1.818643, 1.818645, 1.818645, 1.818648, 1.818649, 1.818649, 
    1.81865, 1.818652, 1.818654, 1.818656, 1.818658, 1.818658, 1.818658, 
    1.818658, 1.818657, 1.818658, 1.818659, 1.818658, 1.818661, 1.81866, 
    1.818661, 1.818661, 1.818646, 1.818647, 1.818646, 1.818647, 1.818647, 
    1.818649, 1.81865, 1.818653, 1.818652, 1.818654, 1.818652, 1.818652, 
    1.818654, 1.818652, 1.818656, 1.818653, 1.818658, 1.818655, 1.818658, 
    1.818658, 1.818659, 1.81866, 1.818661, 1.818663, 1.818662, 1.818664, 
    1.818648, 1.818649, 1.818649, 1.81865, 1.81865, 1.818652, 1.818655, 
    1.818654, 1.818655, 1.818656, 1.818653, 1.818655, 1.818649, 1.81865, 
    1.81865, 1.818648, 1.818654, 1.818651, 1.818656, 1.818655, 1.81866, 
    1.818657, 1.818662, 1.818664, 1.818666, 1.818668, 1.818649, 1.818649, 
    1.81865, 1.818651, 1.818653, 1.818655, 1.818655, 1.818655, 1.818656, 
    1.818657, 1.818655, 1.818657, 1.81865, 1.818654, 1.818648, 1.81865, 
    1.818651, 1.818651, 1.818653, 1.818654, 1.818657, 1.818655, 1.818663, 
    1.81866, 1.81867, 1.818667, 1.818648, 1.818649, 1.818652, 1.818651, 
    1.818655, 1.818656, 1.818657, 1.818658, 1.818658, 1.818659, 1.818658, 
    1.818658, 1.818655, 1.818656, 1.818652, 1.818653, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818656, 1.818656, 1.818658, 1.818655, 1.818664, 
    1.818658, 1.81865, 1.818652, 1.818652, 1.818652, 1.818656, 1.818654, 
    1.818659, 1.818657, 1.818659, 1.818658, 1.818658, 1.818657, 1.818656, 
    1.818654, 1.818653, 1.818652, 1.818652, 1.818653, 1.818656, 1.818658, 
    1.818657, 1.818659, 1.818655, 1.818657, 1.818656, 1.818658, 1.818654, 
    1.818657, 1.818653, 1.818653, 1.818654, 1.818657, 1.818657, 1.818658, 
    1.818657, 1.818656, 1.818655, 1.818654, 1.818654, 1.818653, 1.818652, 
    1.818653, 1.818654, 1.818656, 1.818658, 1.81866, 1.81866, 1.818663, 
    1.818661, 1.818664, 1.818661, 1.818666, 1.818657, 1.818661, 1.818654, 
    1.818655, 1.818656, 1.818659, 1.818658, 1.81866, 1.818655, 1.818653, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.81866, 1.818663, 1.818666, 1.818668, 1.818669, 
    1.81867, 1.81867,
  1.818579, 1.818581, 1.818581, 1.818582, 1.818581, 1.818582, 1.81858, 
    1.818581, 1.81858, 1.818579, 1.818585, 1.818582, 1.818588, 1.818586, 
    1.818591, 1.818588, 1.818591, 1.818591, 1.818593, 1.818592, 1.818595, 
    1.818593, 1.818596, 1.818594, 1.818595, 1.818593, 1.818583, 1.818585, 
    1.818583, 1.818583, 1.818583, 1.818581, 1.818581, 1.818579, 1.818579, 
    1.818581, 1.818583, 1.818582, 1.818584, 1.818584, 1.818587, 1.818586, 
    1.81859, 1.818589, 1.818592, 1.818591, 1.818592, 1.818592, 1.818592, 
    1.818591, 1.818591, 1.81859, 1.818586, 1.818587, 1.818583, 1.818581, 
    1.81858, 1.818579, 1.818579, 1.818579, 1.818581, 1.818582, 1.818583, 
    1.818584, 1.818584, 1.818587, 1.818588, 1.81859, 1.81859, 1.818591, 
    1.818591, 1.818592, 1.818592, 1.818593, 1.818591, 1.818592, 1.818589, 
    1.81859, 1.818585, 1.818582, 1.818582, 1.818581, 1.818579, 1.81858, 
    1.81858, 1.818581, 1.818582, 1.818581, 1.818584, 1.818583, 1.818588, 
    1.818586, 1.818591, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818593, 1.818594, 1.818593, 1.818594, 1.818591, 1.818592, 1.818581, 
    1.818581, 1.818582, 1.81858, 1.81858, 1.818579, 1.81858, 1.818581, 
    1.818582, 1.818582, 1.818583, 1.818584, 1.818586, 1.818588, 1.81859, 
    1.818591, 1.81859, 1.818591, 1.81859, 1.81859, 1.818593, 1.818591, 
    1.818594, 1.818594, 1.818593, 1.818594, 1.818581, 1.818581, 1.81858, 
    1.818581, 1.818579, 1.81858, 1.818581, 1.818583, 1.818583, 1.818584, 
    1.818585, 1.818586, 1.818588, 1.81859, 1.818591, 1.818591, 1.818591, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.818594, 1.818593, 
    1.818594, 1.818594, 1.818581, 1.818582, 1.818581, 1.818582, 1.818582, 
    1.818584, 1.818584, 1.818587, 1.818586, 1.818588, 1.818586, 1.818586, 
    1.818588, 1.818586, 1.81859, 1.818587, 1.818592, 1.818589, 1.818592, 
    1.818591, 1.818592, 1.818593, 1.818594, 1.818595, 1.818595, 1.818596, 
    1.818583, 1.818583, 1.818583, 1.818584, 1.818585, 1.818586, 1.818588, 
    1.818588, 1.818589, 1.818589, 1.818587, 1.818588, 1.818584, 1.818585, 
    1.818584, 1.818583, 1.818588, 1.818585, 1.81859, 1.818588, 1.818593, 
    1.818591, 1.818595, 1.818596, 1.818598, 1.8186, 1.818584, 1.818583, 
    1.818584, 1.818586, 1.818587, 1.818589, 1.818589, 1.818589, 1.81859, 
    1.818591, 1.818589, 1.818591, 1.818585, 1.818588, 1.818583, 1.818585, 
    1.818586, 1.818585, 1.818588, 1.818588, 1.81859, 1.818589, 1.818596, 
    1.818593, 1.818601, 1.818599, 1.818583, 1.818584, 1.818586, 1.818585, 
    1.818589, 1.81859, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818592, 1.818589, 1.81859, 1.818586, 1.818587, 1.818587, 1.818586, 
    1.818588, 1.818589, 1.818589, 1.81859, 1.818591, 1.818589, 1.818596, 
    1.818592, 1.818585, 1.818586, 1.818586, 1.818586, 1.81859, 1.818588, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.818591, 1.81859, 
    1.818588, 1.818587, 1.818586, 1.818586, 1.818587, 1.818589, 1.818591, 
    1.818591, 1.818592, 1.818588, 1.81859, 1.818589, 1.818591, 1.818588, 
    1.818591, 1.818587, 1.818587, 1.818588, 1.81859, 1.818591, 1.818591, 
    1.818591, 1.818589, 1.818589, 1.818588, 1.818588, 1.818587, 1.818586, 
    1.818587, 1.818588, 1.818589, 1.818591, 1.818593, 1.818593, 1.818595, 
    1.818594, 1.818596, 1.818594, 1.818598, 1.818591, 1.818594, 1.818588, 
    1.818589, 1.81859, 1.818592, 1.818591, 1.818593, 1.818589, 1.818587, 
    1.818587, 1.818586, 1.818587, 1.818587, 1.818588, 1.818587, 1.818589, 
    1.818588, 1.818591, 1.818593, 1.818596, 1.818598, 1.8186, 1.818601, 
    1.818601, 1.818601,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.327842e-09, 1.333684e-09, 1.332548e-09, 1.33726e-09, 1.334646e-09, 
    1.337732e-09, 1.329026e-09, 1.333916e-09, 1.330795e-09, 1.328368e-09, 
    1.346405e-09, 1.337471e-09, 1.355685e-09, 1.349987e-09, 1.3643e-09, 
    1.354798e-09, 1.366215e-09, 1.364025e-09, 1.370617e-09, 1.368728e-09, 
    1.377159e-09, 1.371488e-09, 1.38153e-09, 1.375805e-09, 1.376701e-09, 
    1.371301e-09, 1.339268e-09, 1.345293e-09, 1.338912e-09, 1.339771e-09, 
    1.339385e-09, 1.3347e-09, 1.33234e-09, 1.327395e-09, 1.328293e-09, 
    1.331925e-09, 1.340157e-09, 1.337362e-09, 1.344405e-09, 1.344246e-09, 
    1.352087e-09, 1.348551e-09, 1.36173e-09, 1.357984e-09, 1.368807e-09, 
    1.366085e-09, 1.368679e-09, 1.367893e-09, 1.36869e-09, 1.364698e-09, 
    1.366408e-09, 1.362895e-09, 1.349214e-09, 1.353235e-09, 1.341242e-09, 
    1.334031e-09, 1.329241e-09, 1.325842e-09, 1.326322e-09, 1.327239e-09, 
    1.331946e-09, 1.336371e-09, 1.339744e-09, 1.342e-09, 1.344223e-09, 
    1.350952e-09, 1.354513e-09, 1.362487e-09, 1.361048e-09, 1.363486e-09, 
    1.365815e-09, 1.369725e-09, 1.369081e-09, 1.370804e-09, 1.363421e-09, 
    1.368328e-09, 1.360228e-09, 1.362443e-09, 1.344828e-09, 1.338116e-09, 
    1.335264e-09, 1.332767e-09, 1.326692e-09, 1.330887e-09, 1.329233e-09, 
    1.333168e-09, 1.335667e-09, 1.334431e-09, 1.342062e-09, 1.339095e-09, 
    1.354724e-09, 1.347992e-09, 1.365543e-09, 1.361343e-09, 1.36655e-09, 
    1.363893e-09, 1.368445e-09, 1.364348e-09, 1.371445e-09, 1.37299e-09, 
    1.371934e-09, 1.375991e-09, 1.364121e-09, 1.368679e-09, 1.334396e-09, 
    1.334598e-09, 1.335537e-09, 1.331408e-09, 1.331155e-09, 1.327371e-09, 
    1.330738e-09, 1.332172e-09, 1.335812e-09, 1.337966e-09, 1.340012e-09, 
    1.344513e-09, 1.349539e-09, 1.356567e-09, 1.361615e-09, 1.365e-09, 
    1.362924e-09, 1.364757e-09, 1.362709e-09, 1.361748e-09, 1.372411e-09, 
    1.366424e-09, 1.375407e-09, 1.37491e-09, 1.370845e-09, 1.374966e-09, 
    1.33474e-09, 1.333579e-09, 1.32955e-09, 1.332703e-09, 1.326959e-09, 
    1.330174e-09, 1.332023e-09, 1.339157e-09, 1.340725e-09, 1.342178e-09, 
    1.345049e-09, 1.348732e-09, 1.355195e-09, 1.360817e-09, 1.36595e-09, 
    1.365574e-09, 1.365706e-09, 1.366853e-09, 1.364013e-09, 1.367319e-09, 
    1.367874e-09, 1.366423e-09, 1.374844e-09, 1.372438e-09, 1.3749e-09, 
    1.373333e-09, 1.333956e-09, 1.335909e-09, 1.334854e-09, 1.336838e-09, 
    1.33544e-09, 1.341656e-09, 1.343519e-09, 1.352238e-09, 1.34866e-09, 
    1.354355e-09, 1.349238e-09, 1.350145e-09, 1.354541e-09, 1.349515e-09, 
    1.360507e-09, 1.353055e-09, 1.366898e-09, 1.359456e-09, 1.367364e-09, 
    1.365928e-09, 1.368305e-09, 1.370435e-09, 1.373114e-09, 1.378057e-09, 
    1.376913e-09, 1.381046e-09, 1.33882e-09, 1.341352e-09, 1.341129e-09, 
    1.34378e-09, 1.34574e-09, 1.349988e-09, 1.356802e-09, 1.35424e-09, 
    1.358943e-09, 1.359888e-09, 1.352741e-09, 1.357129e-09, 1.343047e-09, 
    1.345323e-09, 1.343968e-09, 1.33902e-09, 1.35483e-09, 1.346716e-09, 
    1.361699e-09, 1.357303e-09, 1.370131e-09, 1.363752e-09, 1.376282e-09, 
    1.381639e-09, 1.386681e-09, 1.392573e-09, 1.342735e-09, 1.341014e-09, 
    1.344095e-09, 1.348358e-09, 1.352313e-09, 1.357571e-09, 1.35811e-09, 
    1.359095e-09, 1.361646e-09, 1.363792e-09, 1.359406e-09, 1.364329e-09, 
    1.345851e-09, 1.355534e-09, 1.340363e-09, 1.344932e-09, 1.348107e-09, 
    1.346714e-09, 1.353947e-09, 1.355651e-09, 1.362579e-09, 1.358998e-09, 
    1.380317e-09, 1.370885e-09, 1.397058e-09, 1.389744e-09, 1.340413e-09, 
    1.342729e-09, 1.35079e-09, 1.346954e-09, 1.357923e-09, 1.360622e-09, 
    1.362817e-09, 1.365623e-09, 1.365925e-09, 1.367588e-09, 1.364864e-09, 
    1.36748e-09, 1.357583e-09, 1.362006e-09, 1.349868e-09, 1.352822e-09, 
    1.351463e-09, 1.349973e-09, 1.354573e-09, 1.359475e-09, 1.35958e-09, 
    1.361152e-09, 1.365581e-09, 1.357967e-09, 1.381535e-09, 1.36698e-09, 
    1.345254e-09, 1.349716e-09, 1.350353e-09, 1.348625e-09, 1.360352e-09, 
    1.356103e-09, 1.367547e-09, 1.364454e-09, 1.369522e-09, 1.367004e-09, 
    1.366633e-09, 1.363399e-09, 1.361385e-09, 1.356297e-09, 1.352158e-09, 
    1.348875e-09, 1.349638e-09, 1.353244e-09, 1.359775e-09, 1.365953e-09, 
    1.3646e-09, 1.369137e-09, 1.357127e-09, 1.362163e-09, 1.360217e-09, 
    1.365292e-09, 1.354172e-09, 1.363642e-09, 1.351751e-09, 1.352793e-09, 
    1.356018e-09, 1.362505e-09, 1.36394e-09, 1.365472e-09, 1.364526e-09, 
    1.359941e-09, 1.359189e-09, 1.35594e-09, 1.355043e-09, 1.352566e-09, 
    1.350516e-09, 1.352389e-09, 1.354357e-09, 1.359943e-09, 1.364977e-09, 
    1.370465e-09, 1.371808e-09, 1.378222e-09, 1.373001e-09, 1.381616e-09, 
    1.374292e-09, 1.38697e-09, 1.36419e-09, 1.374077e-09, 1.356165e-09, 
    1.358095e-09, 1.361585e-09, 1.36959e-09, 1.365268e-09, 1.370322e-09, 
    1.35916e-09, 1.353369e-09, 1.35187e-09, 1.349075e-09, 1.351934e-09, 
    1.351702e-09, 1.354438e-09, 1.353559e-09, 1.360128e-09, 1.356599e-09, 
    1.366624e-09, 1.370282e-09, 1.380613e-09, 1.386947e-09, 1.393393e-09, 
    1.396239e-09, 1.397105e-09, 1.397468e-09 ;

 SOIL2_HR_S3 =
  9.484586e-11, 9.526315e-11, 9.518202e-11, 9.55186e-11, 9.533189e-11, 
    9.555228e-11, 9.493045e-11, 9.527972e-11, 9.505675e-11, 9.488342e-11, 
    9.617179e-11, 9.553362e-11, 9.683462e-11, 9.642763e-11, 9.744998e-11, 
    9.677129e-11, 9.758682e-11, 9.743038e-11, 9.790119e-11, 9.776632e-11, 
    9.836854e-11, 9.796344e-11, 9.868069e-11, 9.827179e-11, 9.833576e-11, 
    9.795009e-11, 9.566203e-11, 9.609234e-11, 9.563654e-11, 9.56979e-11, 
    9.567036e-11, 9.533575e-11, 9.516713e-11, 9.481396e-11, 9.487807e-11, 
    9.513747e-11, 9.572549e-11, 9.552587e-11, 9.602893e-11, 9.601757e-11, 
    9.657761e-11, 9.63251e-11, 9.726639e-11, 9.699886e-11, 9.777194e-11, 
    9.757752e-11, 9.776281e-11, 9.770663e-11, 9.776355e-11, 9.747841e-11, 
    9.760057e-11, 9.734966e-11, 9.63724e-11, 9.665961e-11, 9.580299e-11, 
    9.528792e-11, 9.494577e-11, 9.4703e-11, 9.473732e-11, 9.480275e-11, 
    9.513899e-11, 9.54551e-11, 9.569601e-11, 9.585716e-11, 9.601593e-11, 
    9.649657e-11, 9.675094e-11, 9.73205e-11, 9.72177e-11, 9.739184e-11, 
    9.755818e-11, 9.783747e-11, 9.77915e-11, 9.791455e-11, 9.738723e-11, 
    9.77377e-11, 9.715914e-11, 9.731738e-11, 9.605915e-11, 9.557972e-11, 
    9.537598e-11, 9.519762e-11, 9.47637e-11, 9.506336e-11, 9.494523e-11, 
    9.522625e-11, 9.540482e-11, 9.53165e-11, 9.586156e-11, 9.564966e-11, 
    9.676601e-11, 9.628517e-11, 9.753878e-11, 9.723879e-11, 9.761068e-11, 
    9.742091e-11, 9.774607e-11, 9.745343e-11, 9.796035e-11, 9.807073e-11, 
    9.79953e-11, 9.828505e-11, 9.743721e-11, 9.776282e-11, 9.531403e-11, 
    9.532843e-11, 9.539554e-11, 9.510057e-11, 9.508253e-11, 9.48122e-11, 
    9.505273e-11, 9.515516e-11, 9.541517e-11, 9.556897e-11, 9.571517e-11, 
    9.603662e-11, 9.639562e-11, 9.689761e-11, 9.725824e-11, 9.749999e-11, 
    9.735174e-11, 9.748262e-11, 9.733632e-11, 9.726775e-11, 9.802938e-11, 
    9.760172e-11, 9.824337e-11, 9.820787e-11, 9.791748e-11, 9.821187e-11, 
    9.533855e-11, 9.525566e-11, 9.496788e-11, 9.519309e-11, 9.478276e-11, 
    9.501245e-11, 9.514452e-11, 9.56541e-11, 9.576604e-11, 9.586986e-11, 
    9.607489e-11, 9.633803e-11, 9.679962e-11, 9.720123e-11, 9.756786e-11, 
    9.7541e-11, 9.755045e-11, 9.763235e-11, 9.742948e-11, 9.766566e-11, 
    9.770531e-11, 9.760166e-11, 9.820311e-11, 9.803128e-11, 9.820711e-11, 
    9.809523e-11, 9.52826e-11, 9.542207e-11, 9.534671e-11, 9.548843e-11, 
    9.538859e-11, 9.583254e-11, 9.596565e-11, 9.658847e-11, 9.633285e-11, 
    9.673965e-11, 9.637417e-11, 9.643893e-11, 9.675294e-11, 9.639391e-11, 
    9.71791e-11, 9.664679e-11, 9.763554e-11, 9.710399e-11, 9.766885e-11, 
    9.756627e-11, 9.77361e-11, 9.788822e-11, 9.807957e-11, 9.843266e-11, 
    9.83509e-11, 9.864617e-11, 9.562999e-11, 9.581089e-11, 9.579496e-11, 
    9.598427e-11, 9.612428e-11, 9.642772e-11, 9.691442e-11, 9.673139e-11, 
    9.706738e-11, 9.713483e-11, 9.662438e-11, 9.693781e-11, 9.593196e-11, 
    9.609448e-11, 9.599771e-11, 9.564426e-11, 9.677358e-11, 9.619402e-11, 
    9.72642e-11, 9.695025e-11, 9.786653e-11, 9.741085e-11, 9.830588e-11, 
    9.868853e-11, 9.904861e-11, 9.946946e-11, 9.590961e-11, 9.57867e-11, 
    9.600678e-11, 9.631129e-11, 9.65938e-11, 9.69694e-11, 9.700782e-11, 
    9.707819e-11, 9.726044e-11, 9.741368e-11, 9.710045e-11, 9.74521e-11, 
    9.613219e-11, 9.682389e-11, 9.574023e-11, 9.606656e-11, 9.629333e-11, 
    9.619384e-11, 9.671048e-11, 9.683224e-11, 9.732706e-11, 9.707126e-11, 
    9.85941e-11, 9.792036e-11, 9.978987e-11, 9.926743e-11, 9.574375e-11, 
    9.590919e-11, 9.648497e-11, 9.621102e-11, 9.699447e-11, 9.718731e-11, 
    9.734407e-11, 9.754447e-11, 9.756611e-11, 9.768484e-11, 9.749027e-11, 
    9.767715e-11, 9.69702e-11, 9.728612e-11, 9.641915e-11, 9.663017e-11, 
    9.653309e-11, 9.642661e-11, 9.675524e-11, 9.710537e-11, 9.711284e-11, 
    9.722512e-11, 9.754152e-11, 9.699764e-11, 9.868108e-11, 9.764146e-11, 
    9.608959e-11, 9.640826e-11, 9.645376e-11, 9.633032e-11, 9.716798e-11, 
    9.686447e-11, 9.768195e-11, 9.7461e-11, 9.782301e-11, 9.764312e-11, 
    9.761666e-11, 9.738562e-11, 9.724178e-11, 9.687839e-11, 9.65827e-11, 
    9.634822e-11, 9.640275e-11, 9.666031e-11, 9.712679e-11, 9.756807e-11, 
    9.747141e-11, 9.779549e-11, 9.693766e-11, 9.729737e-11, 9.715834e-11, 
    9.752085e-11, 9.672654e-11, 9.740298e-11, 9.655363e-11, 9.66281e-11, 
    9.685844e-11, 9.732178e-11, 9.742427e-11, 9.753372e-11, 9.746618e-11, 
    9.713862e-11, 9.708496e-11, 9.685284e-11, 9.678876e-11, 9.661189e-11, 
    9.646546e-11, 9.659925e-11, 9.673976e-11, 9.713876e-11, 9.749834e-11, 
    9.789038e-11, 9.798632e-11, 9.844441e-11, 9.807152e-11, 9.868688e-11, 
    9.816374e-11, 9.90693e-11, 9.744216e-11, 9.814833e-11, 9.686892e-11, 
    9.700675e-11, 9.725606e-11, 9.782784e-11, 9.751915e-11, 9.788016e-11, 
    9.708286e-11, 9.666921e-11, 9.656217e-11, 9.636248e-11, 9.656673e-11, 
    9.655012e-11, 9.674556e-11, 9.668275e-11, 9.715201e-11, 9.689995e-11, 
    9.7616e-11, 9.787731e-11, 9.861523e-11, 9.906761e-11, 9.952807e-11, 
    9.973137e-11, 9.979324e-11, 9.981911e-11 ;

 SOIL3C =
  5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782611, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782613, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782613, 
    5.782613, 5.782613 ;

 SOIL3C_TO_SOIL1C =
  2.618456e-11, 2.629973e-11, 2.627734e-11, 2.637024e-11, 2.631871e-11, 
    2.637954e-11, 2.620791e-11, 2.630431e-11, 2.624277e-11, 2.619492e-11, 
    2.655053e-11, 2.637439e-11, 2.673348e-11, 2.662115e-11, 2.690333e-11, 
    2.6716e-11, 2.69411e-11, 2.689792e-11, 2.702787e-11, 2.699064e-11, 
    2.715686e-11, 2.704505e-11, 2.724302e-11, 2.713016e-11, 2.714781e-11, 
    2.704136e-11, 2.640983e-11, 2.65286e-11, 2.64028e-11, 2.641973e-11, 
    2.641213e-11, 2.631977e-11, 2.627323e-11, 2.617575e-11, 2.619345e-11, 
    2.626505e-11, 2.642735e-11, 2.637225e-11, 2.65111e-11, 2.650797e-11, 
    2.666255e-11, 2.659285e-11, 2.685266e-11, 2.677882e-11, 2.699219e-11, 
    2.693853e-11, 2.698967e-11, 2.697417e-11, 2.698988e-11, 2.691117e-11, 
    2.694489e-11, 2.687564e-11, 2.66059e-11, 2.668518e-11, 2.644874e-11, 
    2.630657e-11, 2.621214e-11, 2.614512e-11, 2.61546e-11, 2.617266e-11, 
    2.626546e-11, 2.635272e-11, 2.641921e-11, 2.646369e-11, 2.650751e-11, 
    2.664018e-11, 2.671039e-11, 2.686759e-11, 2.683922e-11, 2.688728e-11, 
    2.693319e-11, 2.701028e-11, 2.699759e-11, 2.703156e-11, 2.688601e-11, 
    2.698274e-11, 2.682306e-11, 2.686673e-11, 2.651944e-11, 2.638711e-11, 
    2.633088e-11, 2.628165e-11, 2.616188e-11, 2.624459e-11, 2.621199e-11, 
    2.628955e-11, 2.633884e-11, 2.631446e-11, 2.646491e-11, 2.640642e-11, 
    2.671455e-11, 2.658183e-11, 2.692784e-11, 2.684504e-11, 2.694768e-11, 
    2.689531e-11, 2.698505e-11, 2.690428e-11, 2.70442e-11, 2.707466e-11, 
    2.705384e-11, 2.713382e-11, 2.689981e-11, 2.698968e-11, 2.631378e-11, 
    2.631776e-11, 2.633628e-11, 2.625486e-11, 2.624988e-11, 2.617527e-11, 
    2.624166e-11, 2.626993e-11, 2.634169e-11, 2.638415e-11, 2.64245e-11, 
    2.651322e-11, 2.661231e-11, 2.675087e-11, 2.685041e-11, 2.691713e-11, 
    2.687622e-11, 2.691234e-11, 2.687196e-11, 2.685303e-11, 2.706325e-11, 
    2.694521e-11, 2.712231e-11, 2.711251e-11, 2.703236e-11, 2.711362e-11, 
    2.632055e-11, 2.629767e-11, 2.621824e-11, 2.62804e-11, 2.616714e-11, 
    2.623054e-11, 2.626699e-11, 2.640764e-11, 2.643854e-11, 2.64672e-11, 
    2.652379e-11, 2.659642e-11, 2.672382e-11, 2.683467e-11, 2.693586e-11, 
    2.692845e-11, 2.693106e-11, 2.695367e-11, 2.689767e-11, 2.696286e-11, 
    2.69738e-11, 2.694519e-11, 2.71112e-11, 2.706377e-11, 2.711231e-11, 
    2.708143e-11, 2.63051e-11, 2.63436e-11, 2.63228e-11, 2.636192e-11, 
    2.633436e-11, 2.64569e-11, 2.649364e-11, 2.666554e-11, 2.659499e-11, 
    2.670727e-11, 2.660639e-11, 2.662427e-11, 2.671094e-11, 2.661184e-11, 
    2.682856e-11, 2.668164e-11, 2.695455e-11, 2.680783e-11, 2.696374e-11, 
    2.693543e-11, 2.69823e-11, 2.702429e-11, 2.70771e-11, 2.717456e-11, 
    2.715199e-11, 2.723349e-11, 2.640099e-11, 2.645092e-11, 2.644652e-11, 
    2.649878e-11, 2.653742e-11, 2.662117e-11, 2.675551e-11, 2.670499e-11, 
    2.679773e-11, 2.681634e-11, 2.667546e-11, 2.676196e-11, 2.648434e-11, 
    2.652919e-11, 2.650248e-11, 2.640493e-11, 2.671664e-11, 2.655667e-11, 
    2.685205e-11, 2.67654e-11, 2.70183e-11, 2.689253e-11, 2.713957e-11, 
    2.724518e-11, 2.734457e-11, 2.746073e-11, 2.647817e-11, 2.644424e-11, 
    2.650499e-11, 2.658904e-11, 2.666701e-11, 2.677068e-11, 2.678129e-11, 
    2.680071e-11, 2.685101e-11, 2.689331e-11, 2.680685e-11, 2.690391e-11, 
    2.65396e-11, 2.673052e-11, 2.643142e-11, 2.652149e-11, 2.658408e-11, 
    2.655662e-11, 2.669922e-11, 2.673283e-11, 2.68694e-11, 2.67988e-11, 
    2.721912e-11, 2.703316e-11, 2.754916e-11, 2.740496e-11, 2.643239e-11, 
    2.647805e-11, 2.663698e-11, 2.656136e-11, 2.67776e-11, 2.683083e-11, 
    2.68741e-11, 2.692941e-11, 2.693538e-11, 2.696815e-11, 2.691445e-11, 
    2.696603e-11, 2.67709e-11, 2.68581e-11, 2.661881e-11, 2.667705e-11, 
    2.665026e-11, 2.662087e-11, 2.671157e-11, 2.680821e-11, 2.681027e-11, 
    2.684126e-11, 2.692859e-11, 2.677848e-11, 2.724313e-11, 2.695618e-11, 
    2.652784e-11, 2.66158e-11, 2.662836e-11, 2.659429e-11, 2.682549e-11, 
    2.674172e-11, 2.696736e-11, 2.690637e-11, 2.700629e-11, 2.695664e-11, 
    2.694934e-11, 2.688556e-11, 2.684587e-11, 2.674556e-11, 2.666395e-11, 
    2.659923e-11, 2.661428e-11, 2.668537e-11, 2.681412e-11, 2.693592e-11, 
    2.690924e-11, 2.699869e-11, 2.676192e-11, 2.686121e-11, 2.682283e-11, 
    2.692289e-11, 2.670365e-11, 2.689036e-11, 2.665593e-11, 2.667648e-11, 
    2.674006e-11, 2.686795e-11, 2.689623e-11, 2.692644e-11, 2.69078e-11, 
    2.681739e-11, 2.680258e-11, 2.673851e-11, 2.672083e-11, 2.6672e-11, 
    2.663159e-11, 2.666852e-11, 2.67073e-11, 2.681743e-11, 2.691668e-11, 
    2.702489e-11, 2.705136e-11, 2.71778e-11, 2.707488e-11, 2.724473e-11, 
    2.710034e-11, 2.735028e-11, 2.690117e-11, 2.709608e-11, 2.674295e-11, 
    2.678099e-11, 2.684981e-11, 2.700763e-11, 2.692242e-11, 2.702207e-11, 
    2.6802e-11, 2.668783e-11, 2.665828e-11, 2.660317e-11, 2.665954e-11, 
    2.665496e-11, 2.67089e-11, 2.669157e-11, 2.682109e-11, 2.675151e-11, 
    2.694915e-11, 2.702128e-11, 2.722495e-11, 2.734981e-11, 2.74769e-11, 
    2.753302e-11, 2.755009e-11, 2.755723e-11 ;

 SOIL3C_vr =
  20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00008, 20.00007, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  5.139921e-21, -5.139921e-21, -2.569961e-21, -2.826957e-20, -7.709882e-21, 
    1.541976e-20, 7.709882e-21, 1.027984e-20, 2.569961e-21, 1.003089e-36, 
    -1.027984e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, -2.569961e-20, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 1.28498e-20, 1.28498e-20, 
    1.027984e-20, 1.027984e-20, 1.798972e-20, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, 2.312965e-20, -2.569961e-21, -1.027984e-20, -7.709882e-21, 
    1.28498e-20, -5.139921e-21, -2.569961e-21, 1.541976e-20, -1.28498e-20, 
    -1.798972e-20, 5.139921e-21, 0, 1.28498e-20, -5.139921e-21, 1.541976e-20, 
    -1.798972e-20, -5.139921e-21, -1.541976e-20, -2.569961e-21, 1.027984e-20, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    1.027984e-20, 1.027984e-20, -1.28498e-20, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 1.541976e-20, -1.798972e-20, -1.003089e-36, 
    -1.027984e-20, -1.003089e-36, 1.28498e-20, 7.709882e-21, -7.709882e-21, 
    -1.003089e-36, -2.569961e-21, 1.003089e-36, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 1.003089e-36, 2.569961e-21, -1.003089e-36, 
    -5.139921e-21, 7.709882e-21, -1.027984e-20, 5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21, 1.027984e-20, -7.709882e-21, 
    0, -2.569961e-21, 0, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 7.709882e-21, -5.139921e-21, -1.027984e-20, 
    1.027984e-20, -2.569961e-21, -1.541976e-20, 0, 0, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 2.055969e-20, 2.569961e-21, 0, 
    1.003089e-36, 1.28498e-20, 2.569961e-21, -1.003089e-36, -1.28498e-20, 
    1.027984e-20, 1.003089e-36, -1.28498e-20, 1.027984e-20, -5.139921e-21, 
    2.569961e-21, 1.28498e-20, -2.569961e-21, 5.139921e-21, 1.798972e-20, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, -1.027984e-20, 2.569961e-20, 
    -7.709882e-21, -7.709882e-21, -1.027984e-20, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, 1.28498e-20, 0, 
    -2.569961e-21, 1.28498e-20, 7.709882e-21, -1.28498e-20, 2.569961e-21, 
    -2.312965e-20, -7.709882e-21, -5.139921e-21, 1.798972e-20, 1.28498e-20, 
    -5.139921e-21, -5.139921e-21, -7.709882e-21, 7.709882e-21, -1.027984e-20, 
    -1.28498e-20, 2.569961e-21, 1.003089e-36, 0, 5.139921e-21, 1.28498e-20, 
    5.139921e-21, 5.139921e-21, -1.003089e-36, 0, -1.28498e-20, 0, 
    -1.28498e-20, 5.139921e-21, 1.28498e-20, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 2.569961e-21, 1.027984e-20, 2.569961e-21, 
    2.569961e-21, -1.003089e-36, 7.709882e-21, 7.709882e-21, 7.709882e-21, 
    1.003089e-36, 2.569961e-21, 0, -1.541976e-20, 1.541976e-20, 
    -2.569961e-21, 1.28498e-20, 7.709882e-21, -5.139921e-21, -2.569961e-21, 
    1.28498e-20, -1.541976e-20, -2.569961e-21, -1.28498e-20, -2.569961e-21, 
    1.798972e-20, -1.003089e-36, 1.027984e-20, 1.027984e-20, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, 1.798972e-20, 5.139921e-21, -7.709882e-21, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 1.003089e-36, 
    5.139921e-21, 7.709882e-21, 7.709882e-21, 7.709882e-21, 2.312965e-20, 
    -7.709882e-21, 1.28498e-20, -2.312965e-20, -5.139921e-21, 5.139921e-21, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 0, -2.569961e-21, 
    -1.541976e-20, -2.569961e-21, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, -1.027984e-20, 7.709882e-21, -2.569961e-21, 
    1.003089e-36, -2.569961e-21, 7.709882e-21, -1.541976e-20, -1.003089e-36, 
    1.027984e-20, -1.798972e-20, 5.139921e-21, -5.139921e-21, 7.709882e-21, 
    1.798972e-20, 2.569961e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -7.709882e-21, 1.28498e-20, -1.027984e-20, -1.28498e-20, -1.28498e-20, 
    -1.027984e-20, 0, 7.709882e-21, 2.569961e-21, -1.027984e-20, 
    5.139921e-21, -1.541976e-20, 1.798972e-20, -1.798972e-20, -1.798972e-20, 
    -2.569961e-21, 1.027984e-20, -7.709882e-21, -1.798972e-20, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, 1.003089e-36, -5.139921e-21, 0, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 1.541976e-20, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, 1.027984e-20, 2.569961e-20, 1.798972e-20, 
    -1.28498e-20, -2.569961e-21, 2.569961e-21, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, -1.28498e-20, 2.569961e-21, 7.709882e-21, 
    1.541976e-20, -2.055969e-20, -1.003089e-36, -2.569961e-21, 7.709882e-21, 
    0, -5.139921e-21, -2.569961e-21, -2.569961e-21, -1.28498e-20, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, 7.709882e-21, -1.798972e-20, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, -1.798972e-20, 
    -7.709882e-21, 7.709882e-21, 1.027984e-20, -2.569961e-21, 1.027984e-20, 
    -1.027984e-20, 5.139921e-21, -5.139921e-21, -2.569961e-21, -1.541976e-20, 
    0, 5.139921e-21, -5.139921e-21, -1.027984e-20, -1.798972e-20, 
    1.027984e-20, 5.139921e-21, -2.569961e-21,
  -2.569961e-21, 1.541976e-20, -5.139921e-21, -7.709882e-21, 5.139921e-21, 
    7.709882e-21, 1.28498e-20, -2.569961e-21, 7.709882e-21, 5.139921e-21, 
    -1.027984e-20, -7.709882e-21, -1.28498e-20, -1.027984e-20, 1.003089e-36, 
    7.709882e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, 1.003089e-36, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, 
    -1.003089e-36, -7.709882e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, 0, 0, -5.139921e-21, -1.541976e-20, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 1.027984e-20, 1.28498e-20, 
    1.027984e-20, 5.139921e-21, 1.027984e-20, 2.569961e-21, -2.569961e-21, 
    -1.003089e-36, -2.569961e-21, 7.709882e-21, 0, 1.027984e-20, 
    7.709882e-21, -1.28498e-20, -5.139921e-21, -1.003089e-36, 5.139921e-21, 
    -1.28498e-20, -5.139921e-21, -2.569961e-21, -5.139921e-21, 2.312965e-20, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    -5.139921e-21, 1.28498e-20, 7.709882e-21, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, 0, 2.569961e-21, 7.709882e-21, 1.003089e-36, 1.541976e-20, 
    2.569961e-21, -2.569961e-21, 7.709882e-21, -1.28498e-20, -2.569961e-21, 
    1.003089e-36, 7.709882e-21, -1.28498e-20, 2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 0, 0, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    0, -1.003089e-36, 1.003089e-36, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 0, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    2.569961e-21, -5.139921e-21, -1.541976e-20, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, -7.709882e-21, 
    -1.28498e-20, -1.027984e-20, 1.541976e-20, 0, 5.139921e-21, 5.139921e-21, 
    -1.003089e-36, -2.569961e-21, 1.28498e-20, 0, -1.027984e-20, 
    2.569961e-21, 7.709882e-21, -1.027984e-20, 0, -7.709882e-21, 
    -2.569961e-21, -1.027984e-20, 1.798972e-20, -5.139921e-21, 0, 
    7.709882e-21, 1.541976e-20, -7.709882e-21, -7.709882e-21, 5.139921e-21, 
    2.569961e-21, -1.027984e-20, -1.28498e-20, -1.027984e-20, 1.003089e-36, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, -7.709882e-21, 0, 
    -2.569961e-21, 5.139921e-21, -1.28498e-20, 1.027984e-20, 2.569961e-21, 
    -1.003089e-36, 1.003089e-36, -2.569961e-21, -7.709882e-21, -2.569961e-21, 
    0, -7.709882e-21, 1.28498e-20, -5.139921e-21, 0, -1.003089e-36, 
    2.569961e-21, -2.569961e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    0, -5.139921e-21, 1.28498e-20, -1.541976e-20, 1.027984e-20, 2.569961e-21, 
    2.569961e-21, 5.139921e-21, 1.027984e-20, 5.139921e-21, -1.798972e-20, 
    -7.709882e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, -1.027984e-20, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, 2.569961e-21, 1.027984e-20, -1.28498e-20, 
    -1.541976e-20, -1.003089e-36, -2.569961e-21, 5.139921e-21, 0, 
    1.027984e-20, 1.027984e-20, 5.139921e-21, 1.28498e-20, 7.709882e-21, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 
    1.027984e-20, -5.139921e-21, -1.003089e-36, 1.027984e-20, -7.709882e-21, 
    5.139921e-21, 1.027984e-20, -7.709882e-21, 2.569961e-21, 1.541976e-20, 
    5.139921e-21, -1.28498e-20, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, 1.003089e-36, 1.28498e-20, 
    -2.569961e-21, 2.569961e-21, -1.027984e-20, 7.709882e-21, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 0, 2.569961e-21, 0, 1.003089e-36, 
    2.569961e-21, -1.541976e-20, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    2.569961e-21, 1.541976e-20, -1.027984e-20, -2.569961e-21, -7.709882e-21, 
    2.569961e-21, 2.569961e-21, 1.28498e-20, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -5.139921e-21, -5.139921e-21, 2.055969e-20, -5.139921e-21, 
    0, -2.569961e-21, 2.569961e-21, 7.709882e-21, -1.027984e-20, 
    7.709882e-21, 5.139921e-21, -5.139921e-21, -7.709882e-21, -5.139921e-21, 
    1.541976e-20, 2.569961e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    7.709882e-21, 0, 1.027984e-20, -5.139921e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, 2.569961e-21,
  2.569961e-21, -1.003089e-36, 7.709882e-21, -1.003089e-36, 5.139921e-21, 
    1.28498e-20, -1.003089e-36, 7.709882e-21, -1.027984e-20, -5.139921e-21, 
    2.569961e-21, 1.027984e-20, 2.569961e-21, -1.027984e-20, -5.139921e-21, 
    -1.541976e-20, 2.569961e-21, 1.798972e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, 1.541976e-20, -5.139921e-21, 
    2.569961e-21, -1.003089e-36, 0, 0, 1.541976e-20, -7.709882e-21, 
    -5.139921e-21, -1.28498e-20, -5.139921e-21, 0, -7.709882e-21, 
    -7.709882e-21, -7.709882e-21, -1.003089e-36, 5.139921e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    1.28498e-20, -1.027984e-20, -1.027984e-20, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -2.569961e-21, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    2.569961e-21, -2.569961e-21, -1.28498e-20, 2.312965e-20, -1.003089e-36, 
    0, -7.709882e-21, 1.28498e-20, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    -7.709882e-21, 7.709882e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    1.541976e-20, 5.139921e-21, 0, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, 1.28498e-20, 7.709882e-21, 5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, -1.28498e-20, -1.027984e-20, -1.003089e-36, 
    0, 2.569961e-21, 5.139921e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, 5.139921e-21, -1.027984e-20, -7.709882e-21, 
    -1.28498e-20, 0, 5.139921e-21, 1.28498e-20, -1.003089e-36, 5.139921e-21, 
    -7.709882e-21, 7.709882e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    -1.027984e-20, -1.003089e-36, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    7.709882e-21, -1.541976e-20, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    -1.003089e-36, 2.569961e-21, 0, -1.798972e-20, 0, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, -1.541976e-20, 1.003089e-36, 
    1.027984e-20, -7.709882e-21, 7.709882e-21, 1.027984e-20, 1.28498e-20, 
    2.569961e-21, 5.139921e-21, 1.28498e-20, 1.28498e-20, -1.28498e-20, 0, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, 1.003089e-36, 7.709882e-21, 
    1.798972e-20, 1.28498e-20, -2.569961e-21, 5.139921e-21, 2.569961e-21, 0, 
    1.28498e-20, -5.139921e-21, 5.139921e-21, 1.28498e-20, -2.569961e-21, 
    5.139921e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, 1.798972e-20, -1.027984e-20, 
    -1.003089e-36, 5.139921e-21, 5.139921e-21, -1.027984e-20, -7.709882e-21, 
    1.28498e-20, 2.569961e-21, 2.569961e-21, 7.709882e-21, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 1.027984e-20, 1.541976e-20, 7.709882e-21, 
    1.027984e-20, 5.139921e-21, 2.569961e-21, -1.541976e-20, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, -2.055969e-20, 2.569961e-21, 
    1.541976e-20, -5.139921e-21, 7.709882e-21, -1.541976e-20, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, 2.569961e-21, 1.541976e-20, 
    -7.709882e-21, 7.709882e-21, 0, 0, -2.569961e-21, 7.709882e-21, 
    1.28498e-20, -2.569961e-21, 0, 1.003089e-36, -7.709882e-21, 
    -1.541976e-20, 5.139921e-21, 1.798972e-20, -1.003089e-36, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, -7.709882e-21, -1.027984e-20, 
    -7.709882e-21, -2.569961e-21, -1.798972e-20, -2.569961e-21, 
    -5.139921e-21, 1.003089e-36, -1.027984e-20, -1.003089e-36, -1.027984e-20, 
    1.027984e-20, 1.027984e-20, -1.027984e-20, 2.569961e-21, 1.027984e-20, 0, 
    -2.569961e-21, 0, 2.569961e-21, -1.541976e-20, -1.798972e-20, 
    -2.569961e-21, 7.709882e-21, -1.28498e-20, -2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -7.709882e-21, 2.312965e-20, -1.027984e-20, 1.027984e-20, 
    -1.003089e-36, -1.027984e-20, 0, -5.139921e-21, -2.569961e-21, 0, 
    -2.569961e-21, 2.569961e-21, 1.28498e-20, 2.569961e-21, 0, 0, 
    7.709882e-21, 1.798972e-20, -5.139921e-21, -7.709882e-21, -2.569961e-21, 
    0, -1.003089e-36, 5.139921e-21, -7.709882e-21, 7.709882e-21, 
    -1.003089e-36, 2.569961e-21, 7.709882e-21, -5.139921e-21, 1.28498e-20, 
    -5.139921e-21, 1.003089e-36, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, -1.28498e-20, 7.709882e-21, 
    -1.28498e-20, -1.003089e-36, 1.28498e-20, -2.569961e-21, 5.139921e-21, 
    7.709882e-21, -2.055969e-20, -1.027984e-20, -1.28498e-20, -5.139921e-21, 
    2.569961e-21, 0, 1.541976e-20, 1.003089e-36, -1.027984e-20, 
    -1.003089e-36, -5.139921e-21, 1.28498e-20, -2.569961e-21, -2.569961e-21, 
    1.027984e-20, 7.709882e-21, 0, 0, -7.709882e-21,
  -7.709882e-21, 1.798972e-20, -5.139921e-21, -7.709882e-21, -5.139921e-21, 
    1.003089e-36, 5.139921e-21, 2.569961e-21, 2.569961e-21, 1.003089e-36, 
    -2.569961e-21, -2.569961e-20, -5.139921e-21, -7.709882e-21, 
    -2.569961e-20, -1.027984e-20, 1.541976e-20, -1.003089e-36, 1.027984e-20, 
    -7.709882e-21, 1.027984e-20, -7.709882e-21, -2.569961e-21, -2.312965e-20, 
    -5.139921e-21, -1.798972e-20, 1.003089e-36, 1.541976e-20, 1.541976e-20, 
    1.28498e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -7.709882e-21, -1.003089e-36, -2.055969e-20, 
    -1.027984e-20, 1.027984e-20, -1.28498e-20, -1.541976e-20, 5.139921e-21, 
    5.139921e-21, 7.709882e-21, 1.28498e-20, 5.139921e-21, -7.709882e-21, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, 7.709882e-21, 7.709882e-21, 
    0, -5.139921e-21, -1.541976e-20, -5.139921e-21, 1.027984e-20, 
    2.569961e-21, 1.003089e-36, -2.569961e-21, -7.709882e-21, 2.569961e-21, 
    1.027984e-20, 7.709882e-21, 5.139921e-21, -2.569961e-21, 1.28498e-20, 
    -2.569961e-21, 1.798972e-20, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, -1.027984e-20, 1.027984e-20, 
    -1.003089e-36, 7.709882e-21, 0, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, -1.003089e-36, 
    -7.709882e-21, -2.569961e-21, 1.027984e-20, -1.28498e-20, 1.003089e-36, 
    1.027984e-20, 5.139921e-21, -7.709882e-21, 1.28498e-20, -1.798972e-20, 
    -5.139921e-21, -2.569961e-21, -2.055969e-20, 1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 1.798972e-20, 2.569961e-21, -2.569961e-21, 
    0, -2.826957e-20, -5.139921e-21, -1.003089e-36, -1.28498e-20, 
    2.826957e-20, 1.28498e-20, 1.003089e-36, -2.569961e-21, 2.569961e-21, 
    1.28498e-20, -1.027984e-20, -7.709882e-21, -7.709882e-21, 7.709882e-21, 
    -2.569961e-20, 1.28498e-20, 5.139921e-21, -1.28498e-20, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 5.139921e-21, -1.541976e-20, -1.003089e-36, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -1.798972e-20, -2.312965e-20, 7.709882e-21, 2.312965e-20, -1.027984e-20, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 1.28498e-20, 2.569961e-21, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, 0, -1.027984e-20, 5.139921e-21, 
    1.541976e-20, -2.569961e-21, -7.709882e-21, -2.569961e-21, -1.28498e-20, 
    1.28498e-20, -5.139921e-21, 2.569961e-21, 1.541976e-20, -1.003089e-36, 
    1.28498e-20, 2.569961e-21, 1.027984e-20, 1.798972e-20, 0, -1.027984e-20, 
    1.003089e-36, 1.027984e-20, 2.569961e-21, -1.541976e-20, -2.569961e-21, 
    -7.709882e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    1.28498e-20, -2.569961e-21, -1.003089e-36, 5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 1.28498e-20, -2.055969e-20, -1.027984e-20, 7.709882e-21, 
    1.28498e-20, -2.569961e-21, 7.709882e-21, 3.009266e-36, -1.027984e-20, 
    1.28498e-20, -1.798972e-20, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -1.003089e-36, 5.139921e-21, -5.139921e-21, -1.003089e-36, 1.541976e-20, 
    -5.139921e-21, -2.569961e-21, 1.28498e-20, -1.798972e-20, -5.139921e-21, 
    0, -7.709882e-21, 1.541976e-20, 0, -1.798972e-20, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    7.709882e-21, -5.139921e-21, -1.28498e-20, 5.139921e-21, 5.139921e-21, 
    -1.003089e-36, -1.027984e-20, 2.569961e-21, -7.709882e-21, -5.139921e-21, 
    5.139921e-21, -1.003089e-36, 2.569961e-21, 2.569961e-21, -1.28498e-20, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, -1.003089e-36, 1.027984e-20, 
    2.569961e-21, 1.003089e-36, 2.569961e-21, 1.003089e-36, -1.027984e-20, 
    2.569961e-21, -5.139921e-21, 1.003089e-36, 1.003089e-36, -1.003089e-36, 
    -1.027984e-20, 0, 1.003089e-36, 5.139921e-21, -5.139921e-21, 
    -2.312965e-20, 7.709882e-21, -1.027984e-20, 7.709882e-21, 0, 
    1.541976e-20, 1.003089e-36, -5.139921e-21, -1.003089e-36, 7.709882e-21, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, -7.709882e-21, -1.027984e-20, 
    -2.569961e-21, -2.569961e-21, 1.28498e-20, 2.569961e-21, 1.541976e-20, 
    -2.055969e-20, -2.312965e-20, -7.709882e-21, 5.139921e-21, 1.027984e-20, 
    7.709882e-21, 7.709882e-21, 1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -1.541976e-20, 0, 7.709882e-21, -1.003089e-36, -1.798972e-20, 
    2.569961e-21, -1.28498e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, 2.055969e-20, 5.139921e-21, -1.798972e-20, -7.709882e-21, 
    -2.055969e-20, 7.709882e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -1.798972e-20, -5.139921e-21, -7.709882e-21, 2.569961e-21, 
    1.541976e-20, 5.139921e-21, -7.709882e-21, -1.027984e-20, -7.709882e-21, 
    2.569961e-21, 2.569961e-21, 7.709882e-21, -1.003089e-36, 2.569961e-21, 
    -1.28498e-20, 1.003089e-36, 7.709882e-21, -1.541976e-20, 2.569961e-21, 
    -5.139921e-21, 1.003089e-36,
  5.139921e-21, -2.569961e-20, 1.003089e-36, 1.541976e-20, -2.569961e-21, 
    5.139921e-21, -5.139921e-21, -2.569961e-20, 1.003089e-36, -1.027984e-20, 
    5.139921e-21, -2.569961e-20, 1.003089e-36, 5.139921e-21, -2.569961e-21, 
    1.003089e-36, 1.003089e-36, 5.139921e-21, -1.798972e-20, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, -1.28498e-20, 5.139921e-21, 
    1.003089e-36, 5.139921e-21, -1.027984e-20, -2.569961e-21, -7.709882e-21, 
    -2.569961e-21, 1.003089e-36, -5.139921e-21, -2.055969e-20, 2.569961e-21, 
    7.709882e-21, -1.798972e-20, -7.709882e-21, -7.709882e-21, 1.027984e-20, 
    -7.709882e-21, 1.541976e-20, -1.003089e-36, 1.28498e-20, -5.139921e-21, 
    2.569961e-21, 1.027984e-20, -1.027984e-20, -2.569961e-21, 2.569961e-21, 
    2.055969e-20, 1.541976e-20, 2.569961e-21, -1.541976e-20, -5.139921e-21, 
    2.569961e-21, -1.798972e-20, 1.541976e-20, 1.28498e-20, -1.798972e-20, 
    1.027984e-20, -1.003089e-36, 5.139921e-21, 2.569961e-21, 1.28498e-20, 
    -1.541976e-20, 7.709882e-21, 7.709882e-21, 1.28498e-20, -1.798972e-20, 
    1.541976e-20, 2.826957e-20, -1.798972e-20, -2.569961e-21, -5.139921e-21, 
    2.569961e-20, 2.569961e-21, 1.798972e-20, 1.027984e-20, -2.569961e-21, 
    -7.709882e-21, -1.027984e-20, 1.003089e-36, 1.28498e-20, -1.28498e-20, 
    2.569961e-21, -1.541976e-20, 7.709882e-21, -5.139921e-21, 3.340949e-20, 
    5.139921e-21, 1.003089e-36, 1.798972e-20, -7.709882e-21, 0, 1.798972e-20, 
    7.709882e-21, 1.541976e-20, 5.139921e-21, 1.798972e-20, -5.139921e-21, 
    7.709882e-21, 2.055969e-20, 5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -2.055969e-20, 1.541976e-20, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 1.28498e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    1.027984e-20, -1.798972e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, 
    -1.541976e-20, -5.139921e-21, -2.569961e-21, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21, 7.709882e-21, 1.003089e-36, 
    -2.569961e-21, 2.312965e-20, 5.139921e-21, -2.569961e-21, 5.139921e-21, 
    7.709882e-21, 1.027984e-20, -7.709882e-21, -1.541976e-20, 7.709882e-21, 
    -2.569961e-20, 7.709882e-21, -2.569961e-21, 2.569961e-21, -1.027984e-20, 
    2.569961e-21, -7.709882e-21, -2.055969e-20, -1.027984e-20, 1.541976e-20, 
    -5.139921e-21, -1.28498e-20, 1.541976e-20, -2.569961e-21, 2.569961e-21, 
    1.28498e-20, 7.709882e-21, -5.139921e-21, 1.28498e-20, 2.569961e-21, 
    1.28498e-20, -7.709882e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, 
    2.569961e-21, -1.541976e-20, -1.28498e-20, -2.569961e-21, -1.541976e-20, 
    5.139921e-21, 2.569961e-21, -1.28498e-20, 7.709882e-21, 1.003089e-36, 
    -5.139921e-21, -7.709882e-21, -5.139921e-21, 0, 1.003089e-36, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, 0, -2.055969e-20, -5.139921e-21, 
    -5.139921e-21, 1.28498e-20, -1.027984e-20, -1.003089e-36, 1.28498e-20, 
    3.009266e-36, -2.312965e-20, -1.027984e-20, -5.139921e-21, 2.569961e-21, 
    2.569961e-20, 7.709882e-21, -1.027984e-20, 2.569961e-21, -3.083953e-20, 
    2.569961e-21, 5.139921e-21, -1.003089e-36, 7.709882e-21, -1.003089e-36, 
    2.569961e-21, -1.28498e-20, -2.569961e-21, -7.709882e-21, 1.027984e-20, 
    -7.709882e-21, -5.139921e-21, -1.541976e-20, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, 2.055969e-20, -2.569961e-21, 1.027984e-20, 1.798972e-20, 
    -2.569961e-21, -1.28498e-20, 1.003089e-36, 2.569961e-21, 5.139921e-21, 
    -2.826957e-20, 7.709882e-21, 2.569961e-21, 1.027984e-20, 1.003089e-36, 
    -5.139921e-21, -1.541976e-20, -2.055969e-20, 2.312965e-20, -1.027984e-20, 
    1.003089e-36, -2.569961e-21, 1.798972e-20, -1.003089e-36, 1.28498e-20, 0, 
    -1.541976e-20, -1.541976e-20, -1.003089e-36, 7.709882e-21, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, 1.003089e-36, 2.569961e-21, -5.139921e-21, 1.003089e-36, 
    -1.541976e-20, 1.003089e-36, 7.709882e-21, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-20, -2.569961e-21, -2.569961e-21, -1.798972e-20, 
    -7.709882e-21, 7.709882e-21, 7.709882e-21, 1.28498e-20, 7.709882e-21, 
    -1.003089e-36, 1.027984e-20, 1.28498e-20, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, -2.569961e-21, 2.569961e-21, 7.709882e-21, -7.709882e-21, 
    1.027984e-20, -7.709882e-21, -1.003089e-36, 5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -1.027984e-20, 1.798972e-20, -1.28498e-20, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, -7.709882e-21, -1.541976e-20, 
    2.569961e-21, 1.541976e-20, 2.569961e-21, 5.139921e-21, 1.027984e-20, 
    -1.28498e-20, 5.139921e-21, 5.139921e-21, 1.28498e-20, 1.003089e-36, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, -1.798972e-20, -5.139921e-21, 
    -1.28498e-20, 1.003089e-36, 5.139921e-21, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, 1.28498e-20, 5.139921e-21, -2.826957e-20, 7.709882e-21, 
    2.569961e-21, 1.28498e-20, 7.709882e-21, -2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, -5.139921e-21, 1.798972e-20, 
    7.709882e-21, 1.027984e-20,
  6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.28981e-12, 5.313078e-12, 5.308554e-12, 5.327322e-12, 5.316911e-12, 
    5.3292e-12, 5.294527e-12, 5.314002e-12, 5.301569e-12, 5.291904e-12, 
    5.363744e-12, 5.328159e-12, 5.400703e-12, 5.37801e-12, 5.435016e-12, 
    5.397172e-12, 5.442646e-12, 5.433923e-12, 5.460176e-12, 5.452655e-12, 
    5.486234e-12, 5.463647e-12, 5.50364e-12, 5.48084e-12, 5.484407e-12, 
    5.462902e-12, 5.33532e-12, 5.359314e-12, 5.333898e-12, 5.33732e-12, 
    5.335784e-12, 5.317126e-12, 5.307724e-12, 5.288031e-12, 5.291606e-12, 
    5.30607e-12, 5.338858e-12, 5.327727e-12, 5.355778e-12, 5.355145e-12, 
    5.386373e-12, 5.372293e-12, 5.424779e-12, 5.409862e-12, 5.452969e-12, 
    5.442128e-12, 5.45246e-12, 5.449327e-12, 5.4525e-12, 5.436601e-12, 
    5.443413e-12, 5.429422e-12, 5.37493e-12, 5.390945e-12, 5.34318e-12, 
    5.314459e-12, 5.295381e-12, 5.281844e-12, 5.283757e-12, 5.287406e-12, 
    5.306154e-12, 5.323781e-12, 5.337214e-12, 5.3462e-12, 5.355054e-12, 
    5.381854e-12, 5.396037e-12, 5.427796e-12, 5.422064e-12, 5.431774e-12, 
    5.441049e-12, 5.456623e-12, 5.454059e-12, 5.460921e-12, 5.431517e-12, 
    5.451059e-12, 5.418799e-12, 5.427623e-12, 5.357463e-12, 5.33073e-12, 
    5.31937e-12, 5.309424e-12, 5.285229e-12, 5.301938e-12, 5.295351e-12, 
    5.311021e-12, 5.320978e-12, 5.316053e-12, 5.346446e-12, 5.33463e-12, 
    5.396878e-12, 5.370066e-12, 5.439967e-12, 5.42324e-12, 5.443976e-12, 
    5.433395e-12, 5.451526e-12, 5.435209e-12, 5.463474e-12, 5.469629e-12, 
    5.465423e-12, 5.481579e-12, 5.434304e-12, 5.45246e-12, 5.315915e-12, 
    5.316718e-12, 5.32046e-12, 5.304012e-12, 5.303006e-12, 5.287933e-12, 
    5.301345e-12, 5.307056e-12, 5.321554e-12, 5.33013e-12, 5.338283e-12, 
    5.356207e-12, 5.376225e-12, 5.404216e-12, 5.424325e-12, 5.437804e-12, 
    5.429539e-12, 5.436836e-12, 5.428678e-12, 5.424855e-12, 5.467323e-12, 
    5.443477e-12, 5.479256e-12, 5.477275e-12, 5.461084e-12, 5.477499e-12, 
    5.317282e-12, 5.31266e-12, 5.296614e-12, 5.309172e-12, 5.286291e-12, 
    5.299099e-12, 5.306463e-12, 5.334878e-12, 5.341119e-12, 5.346909e-12, 
    5.358341e-12, 5.373013e-12, 5.398752e-12, 5.421146e-12, 5.441589e-12, 
    5.440091e-12, 5.440618e-12, 5.445185e-12, 5.433873e-12, 5.447043e-12, 
    5.449253e-12, 5.443474e-12, 5.47701e-12, 5.467429e-12, 5.477233e-12, 
    5.470995e-12, 5.314163e-12, 5.32194e-12, 5.317737e-12, 5.32564e-12, 
    5.320073e-12, 5.344828e-12, 5.352249e-12, 5.386978e-12, 5.372725e-12, 
    5.395408e-12, 5.375029e-12, 5.37864e-12, 5.396149e-12, 5.37613e-12, 
    5.419912e-12, 5.39023e-12, 5.445363e-12, 5.415724e-12, 5.44722e-12, 
    5.441501e-12, 5.45097e-12, 5.459452e-12, 5.470122e-12, 5.48981e-12, 
    5.485251e-12, 5.501715e-12, 5.333533e-12, 5.343621e-12, 5.342732e-12, 
    5.353288e-12, 5.361095e-12, 5.378015e-12, 5.405153e-12, 5.394948e-12, 
    5.413683e-12, 5.417443e-12, 5.388981e-12, 5.406457e-12, 5.350371e-12, 
    5.359433e-12, 5.354037e-12, 5.334329e-12, 5.3973e-12, 5.364984e-12, 
    5.424657e-12, 5.407151e-12, 5.458243e-12, 5.432834e-12, 5.482741e-12, 
    5.504077e-12, 5.524155e-12, 5.547621e-12, 5.349125e-12, 5.342271e-12, 
    5.354543e-12, 5.371523e-12, 5.387275e-12, 5.408219e-12, 5.410361e-12, 
    5.414285e-12, 5.424447e-12, 5.432992e-12, 5.415526e-12, 5.435134e-12, 
    5.361536e-12, 5.400105e-12, 5.33968e-12, 5.357876e-12, 5.370522e-12, 
    5.364974e-12, 5.393781e-12, 5.400571e-12, 5.428161e-12, 5.413899e-12, 
    5.498812e-12, 5.461244e-12, 5.565487e-12, 5.536357e-12, 5.339877e-12, 
    5.349101e-12, 5.381207e-12, 5.365931e-12, 5.409616e-12, 5.420369e-12, 
    5.42911e-12, 5.440285e-12, 5.441491e-12, 5.448112e-12, 5.437263e-12, 
    5.447683e-12, 5.408263e-12, 5.425879e-12, 5.377537e-12, 5.389304e-12, 
    5.38389e-12, 5.377953e-12, 5.396278e-12, 5.415801e-12, 5.416217e-12, 
    5.422478e-12, 5.44012e-12, 5.409793e-12, 5.503662e-12, 5.445693e-12, 
    5.359161e-12, 5.37693e-12, 5.379467e-12, 5.372584e-12, 5.419291e-12, 
    5.402368e-12, 5.44795e-12, 5.435631e-12, 5.455816e-12, 5.445786e-12, 
    5.44431e-12, 5.431427e-12, 5.423407e-12, 5.403144e-12, 5.386656e-12, 
    5.373582e-12, 5.376622e-12, 5.390984e-12, 5.416995e-12, 5.441601e-12, 
    5.436211e-12, 5.454282e-12, 5.406449e-12, 5.426506e-12, 5.418754e-12, 
    5.438968e-12, 5.394677e-12, 5.432395e-12, 5.385036e-12, 5.389188e-12, 
    5.402032e-12, 5.427868e-12, 5.433582e-12, 5.439686e-12, 5.43592e-12, 
    5.417655e-12, 5.414663e-12, 5.401719e-12, 5.398146e-12, 5.388284e-12, 
    5.380119e-12, 5.387579e-12, 5.395414e-12, 5.417662e-12, 5.437713e-12, 
    5.459573e-12, 5.464922e-12, 5.490465e-12, 5.469673e-12, 5.503985e-12, 
    5.474815e-12, 5.525309e-12, 5.43458e-12, 5.473956e-12, 5.402616e-12, 
    5.410302e-12, 5.424203e-12, 5.456086e-12, 5.438872e-12, 5.459003e-12, 
    5.414545e-12, 5.39148e-12, 5.385511e-12, 5.374377e-12, 5.385766e-12, 
    5.38484e-12, 5.395738e-12, 5.392236e-12, 5.418401e-12, 5.404346e-12, 
    5.444273e-12, 5.458844e-12, 5.49999e-12, 5.525214e-12, 5.55089e-12, 
    5.562225e-12, 5.565676e-12, 5.567118e-12 ;

 SOIL3N_vr =
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818188, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.200335e-11, 3.214412e-11, 3.211675e-11, 3.22303e-11, 3.216731e-11, 
    3.224166e-11, 3.203189e-11, 3.214971e-11, 3.207449e-11, 3.201602e-11, 
    3.245065e-11, 3.223536e-11, 3.267426e-11, 3.253696e-11, 3.288185e-11, 
    3.265289e-11, 3.292801e-11, 3.287524e-11, 3.303406e-11, 3.298856e-11, 
    3.319172e-11, 3.305506e-11, 3.329702e-11, 3.315908e-11, 3.318066e-11, 
    3.305056e-11, 3.227868e-11, 3.242385e-11, 3.227009e-11, 3.229078e-11, 
    3.228149e-11, 3.216861e-11, 3.211173e-11, 3.199259e-11, 3.201422e-11, 
    3.210172e-11, 3.230009e-11, 3.223275e-11, 3.240246e-11, 3.239863e-11, 
    3.258755e-11, 3.250237e-11, 3.281991e-11, 3.272966e-11, 3.299046e-11, 
    3.292487e-11, 3.298738e-11, 3.296843e-11, 3.298763e-11, 3.289144e-11, 
    3.293265e-11, 3.284801e-11, 3.251832e-11, 3.261522e-11, 3.232624e-11, 
    3.215248e-11, 3.203706e-11, 3.195515e-11, 3.196673e-11, 3.19888e-11, 
    3.210223e-11, 3.220888e-11, 3.229015e-11, 3.234451e-11, 3.239807e-11, 
    3.256022e-11, 3.264603e-11, 3.283817e-11, 3.280349e-11, 3.286223e-11, 
    3.291835e-11, 3.301257e-11, 3.299706e-11, 3.303857e-11, 3.286068e-11, 
    3.297891e-11, 3.278373e-11, 3.283711e-11, 3.241265e-11, 3.225092e-11, 
    3.218219e-11, 3.212201e-11, 3.197563e-11, 3.207672e-11, 3.203687e-11, 
    3.213168e-11, 3.219192e-11, 3.216212e-11, 3.2346e-11, 3.227451e-11, 
    3.265111e-11, 3.24889e-11, 3.29118e-11, 3.28106e-11, 3.293606e-11, 
    3.287204e-11, 3.298173e-11, 3.288301e-11, 3.305402e-11, 3.309126e-11, 
    3.306581e-11, 3.316356e-11, 3.287754e-11, 3.298738e-11, 3.216129e-11, 
    3.216614e-11, 3.218878e-11, 3.208928e-11, 3.208319e-11, 3.199199e-11, 
    3.207314e-11, 3.210769e-11, 3.219541e-11, 3.224729e-11, 3.229661e-11, 
    3.240505e-11, 3.252616e-11, 3.269551e-11, 3.281717e-11, 3.289872e-11, 
    3.284871e-11, 3.289286e-11, 3.284351e-11, 3.282037e-11, 3.30773e-11, 
    3.293303e-11, 3.314949e-11, 3.313752e-11, 3.303956e-11, 3.313887e-11, 
    3.216956e-11, 3.214159e-11, 3.204451e-11, 3.212049e-11, 3.198206e-11, 
    3.205955e-11, 3.21041e-11, 3.227601e-11, 3.231377e-11, 3.23488e-11, 
    3.241796e-11, 3.250673e-11, 3.266245e-11, 3.279793e-11, 3.292161e-11, 
    3.291255e-11, 3.291574e-11, 3.294337e-11, 3.287493e-11, 3.295461e-11, 
    3.296798e-11, 3.293301e-11, 3.313591e-11, 3.307795e-11, 3.313726e-11, 
    3.309952e-11, 3.215068e-11, 3.219773e-11, 3.217231e-11, 3.222012e-11, 
    3.218644e-11, 3.233621e-11, 3.238111e-11, 3.259121e-11, 3.250498e-11, 
    3.264222e-11, 3.251893e-11, 3.254077e-11, 3.26467e-11, 3.252559e-11, 
    3.279046e-11, 3.261089e-11, 3.294445e-11, 3.276513e-11, 3.295568e-11, 
    3.292108e-11, 3.297837e-11, 3.302968e-11, 3.309424e-11, 3.321335e-11, 
    3.318577e-11, 3.328538e-11, 3.226788e-11, 3.23289e-11, 3.232353e-11, 
    3.238739e-11, 3.243462e-11, 3.253699e-11, 3.270118e-11, 3.263943e-11, 
    3.275278e-11, 3.277553e-11, 3.260333e-11, 3.270906e-11, 3.236975e-11, 
    3.242457e-11, 3.239193e-11, 3.227269e-11, 3.265367e-11, 3.245815e-11, 
    3.281917e-11, 3.271326e-11, 3.302237e-11, 3.286865e-11, 3.317058e-11, 
    3.329967e-11, 3.342114e-11, 3.356311e-11, 3.236221e-11, 3.232074e-11, 
    3.239499e-11, 3.249771e-11, 3.259302e-11, 3.271972e-11, 3.273268e-11, 
    3.275642e-11, 3.28179e-11, 3.28696e-11, 3.276393e-11, 3.288256e-11, 
    3.243729e-11, 3.267064e-11, 3.230506e-11, 3.241515e-11, 3.249166e-11, 
    3.245809e-11, 3.263238e-11, 3.267345e-11, 3.284038e-11, 3.275409e-11, 
    3.326781e-11, 3.304053e-11, 3.36712e-11, 3.349496e-11, 3.230625e-11, 
    3.236206e-11, 3.25563e-11, 3.246389e-11, 3.272818e-11, 3.279323e-11, 
    3.284612e-11, 3.291372e-11, 3.292102e-11, 3.296108e-11, 3.289544e-11, 
    3.295848e-11, 3.271999e-11, 3.282657e-11, 3.25341e-11, 3.260529e-11, 
    3.257253e-11, 3.253662e-11, 3.264748e-11, 3.27656e-11, 3.276811e-11, 
    3.280599e-11, 3.291273e-11, 3.272925e-11, 3.329716e-11, 3.294644e-11, 
    3.242292e-11, 3.253043e-11, 3.254578e-11, 3.250413e-11, 3.278671e-11, 
    3.268432e-11, 3.29601e-11, 3.288557e-11, 3.300769e-11, 3.2947e-11, 
    3.293808e-11, 3.286013e-11, 3.281161e-11, 3.268902e-11, 3.258927e-11, 
    3.251017e-11, 3.252856e-11, 3.261546e-11, 3.277282e-11, 3.292168e-11, 
    3.288908e-11, 3.299841e-11, 3.270902e-11, 3.283037e-11, 3.278346e-11, 
    3.290575e-11, 3.26378e-11, 3.286599e-11, 3.257947e-11, 3.260459e-11, 
    3.268229e-11, 3.28386e-11, 3.287317e-11, 3.29101e-11, 3.288731e-11, 
    3.277681e-11, 3.275871e-11, 3.26804e-11, 3.265879e-11, 3.259912e-11, 
    3.254972e-11, 3.259485e-11, 3.264225e-11, 3.277686e-11, 3.289816e-11, 
    3.303042e-11, 3.306278e-11, 3.321731e-11, 3.309152e-11, 3.329911e-11, 
    3.312263e-11, 3.342812e-11, 3.287921e-11, 3.311743e-11, 3.268583e-11, 
    3.273232e-11, 3.281643e-11, 3.300932e-11, 3.290518e-11, 3.302697e-11, 
    3.2758e-11, 3.261846e-11, 3.258234e-11, 3.251498e-11, 3.258388e-11, 
    3.257828e-11, 3.264421e-11, 3.262303e-11, 3.278133e-11, 3.269629e-11, 
    3.293785e-11, 3.302601e-11, 3.327494e-11, 3.342755e-11, 3.358288e-11, 
    3.365146e-11, 3.367234e-11, 3.368106e-11 ;

 SOILC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.34459, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34452, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34455, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34452, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.3445, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.34449, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34456, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34455, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34455, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 SOILC_HR =
  6.359073e-08, 6.38703e-08, 6.381595e-08, 6.404144e-08, 6.391635e-08, 
    6.406401e-08, 6.364741e-08, 6.38814e-08, 6.373202e-08, 6.361589e-08, 
    6.447906e-08, 6.405151e-08, 6.492314e-08, 6.465046e-08, 6.533541e-08, 
    6.488071e-08, 6.542709e-08, 6.532228e-08, 6.563771e-08, 6.554734e-08, 
    6.595081e-08, 6.567942e-08, 6.615994e-08, 6.588599e-08, 6.592885e-08, 
    6.567046e-08, 6.413754e-08, 6.442583e-08, 6.412046e-08, 6.416157e-08, 
    6.414312e-08, 6.391894e-08, 6.380597e-08, 6.356935e-08, 6.36123e-08, 
    6.37861e-08, 6.418006e-08, 6.404632e-08, 6.438335e-08, 6.437574e-08, 
    6.475095e-08, 6.458178e-08, 6.521241e-08, 6.503318e-08, 6.555111e-08, 
    6.542086e-08, 6.5545e-08, 6.550735e-08, 6.554549e-08, 6.535446e-08, 
    6.54363e-08, 6.52682e-08, 6.461346e-08, 6.480589e-08, 6.423198e-08, 
    6.388689e-08, 6.365767e-08, 6.349501e-08, 6.3518e-08, 6.356184e-08, 
    6.378711e-08, 6.39989e-08, 6.41603e-08, 6.426826e-08, 6.437465e-08, 
    6.469666e-08, 6.486707e-08, 6.524866e-08, 6.517979e-08, 6.529645e-08, 
    6.54079e-08, 6.559502e-08, 6.556422e-08, 6.564666e-08, 6.529337e-08, 
    6.552817e-08, 6.514056e-08, 6.524657e-08, 6.440359e-08, 6.408239e-08, 
    6.39459e-08, 6.38264e-08, 6.353569e-08, 6.373644e-08, 6.36573e-08, 
    6.384558e-08, 6.396522e-08, 6.390604e-08, 6.427122e-08, 6.412925e-08, 
    6.487718e-08, 6.455502e-08, 6.53949e-08, 6.519392e-08, 6.544307e-08, 
    6.531594e-08, 6.553378e-08, 6.533772e-08, 6.567733e-08, 6.575129e-08, 
    6.570075e-08, 6.589487e-08, 6.532685e-08, 6.5545e-08, 6.390439e-08, 
    6.391404e-08, 6.395899e-08, 6.376138e-08, 6.374928e-08, 6.356817e-08, 
    6.372932e-08, 6.379795e-08, 6.397214e-08, 6.407519e-08, 6.417314e-08, 
    6.43885e-08, 6.462902e-08, 6.496534e-08, 6.520695e-08, 6.536891e-08, 
    6.52696e-08, 6.535728e-08, 6.525926e-08, 6.521332e-08, 6.572358e-08, 
    6.543706e-08, 6.586696e-08, 6.584317e-08, 6.564862e-08, 6.584585e-08, 
    6.392082e-08, 6.386528e-08, 6.367247e-08, 6.382336e-08, 6.354846e-08, 
    6.370234e-08, 6.379082e-08, 6.413222e-08, 6.420723e-08, 6.427678e-08, 
    6.441415e-08, 6.459044e-08, 6.489969e-08, 6.516876e-08, 6.541438e-08, 
    6.539639e-08, 6.540272e-08, 6.54576e-08, 6.532167e-08, 6.547991e-08, 
    6.550647e-08, 6.543703e-08, 6.583998e-08, 6.572486e-08, 6.584266e-08, 
    6.57677e-08, 6.388333e-08, 6.397677e-08, 6.392628e-08, 6.402123e-08, 
    6.395434e-08, 6.425178e-08, 6.434096e-08, 6.475822e-08, 6.458697e-08, 
    6.485951e-08, 6.461465e-08, 6.465804e-08, 6.486842e-08, 6.462788e-08, 
    6.515393e-08, 6.47973e-08, 6.545973e-08, 6.510361e-08, 6.548205e-08, 
    6.541332e-08, 6.55271e-08, 6.562901e-08, 6.575721e-08, 6.599377e-08, 
    6.593899e-08, 6.613681e-08, 6.411607e-08, 6.423728e-08, 6.42266e-08, 
    6.435343e-08, 6.444724e-08, 6.465053e-08, 6.49766e-08, 6.485399e-08, 
    6.507909e-08, 6.512427e-08, 6.478229e-08, 6.499227e-08, 6.431839e-08, 
    6.442727e-08, 6.436243e-08, 6.412564e-08, 6.488224e-08, 6.449396e-08, 
    6.521095e-08, 6.500061e-08, 6.561448e-08, 6.530919e-08, 6.590884e-08, 
    6.616519e-08, 6.640643e-08, 6.668839e-08, 6.430341e-08, 6.422106e-08, 
    6.436851e-08, 6.457253e-08, 6.47618e-08, 6.501344e-08, 6.503917e-08, 
    6.508632e-08, 6.520843e-08, 6.531109e-08, 6.510123e-08, 6.533683e-08, 
    6.445253e-08, 6.491594e-08, 6.418993e-08, 6.440856e-08, 6.45605e-08, 
    6.449384e-08, 6.483997e-08, 6.492154e-08, 6.525305e-08, 6.508168e-08, 
    6.610193e-08, 6.565055e-08, 6.690304e-08, 6.655304e-08, 6.419229e-08, 
    6.430313e-08, 6.468889e-08, 6.450534e-08, 6.503023e-08, 6.515943e-08, 
    6.526445e-08, 6.539872e-08, 6.541321e-08, 6.549276e-08, 6.53624e-08, 
    6.54876e-08, 6.501397e-08, 6.522563e-08, 6.464479e-08, 6.478616e-08, 
    6.472112e-08, 6.464978e-08, 6.486996e-08, 6.510454e-08, 6.510954e-08, 
    6.518476e-08, 6.539673e-08, 6.503235e-08, 6.61602e-08, 6.546369e-08, 
    6.442399e-08, 6.46375e-08, 6.466798e-08, 6.458527e-08, 6.514647e-08, 
    6.494314e-08, 6.549082e-08, 6.53428e-08, 6.558533e-08, 6.546481e-08, 
    6.544708e-08, 6.529229e-08, 6.519593e-08, 6.495246e-08, 6.475436e-08, 
    6.459727e-08, 6.46338e-08, 6.480636e-08, 6.511888e-08, 6.541453e-08, 
    6.534977e-08, 6.556689e-08, 6.499217e-08, 6.523317e-08, 6.514002e-08, 
    6.538289e-08, 6.485072e-08, 6.530392e-08, 6.473489e-08, 6.478478e-08, 
    6.49391e-08, 6.524952e-08, 6.531818e-08, 6.539152e-08, 6.534626e-08, 
    6.512681e-08, 6.509086e-08, 6.493535e-08, 6.489241e-08, 6.477391e-08, 
    6.467581e-08, 6.476544e-08, 6.485958e-08, 6.51269e-08, 6.536781e-08, 
    6.563047e-08, 6.569473e-08, 6.600164e-08, 6.575182e-08, 6.616408e-08, 
    6.58136e-08, 6.642029e-08, 6.533017e-08, 6.580328e-08, 6.494612e-08, 
    6.503846e-08, 6.520549e-08, 6.558857e-08, 6.538175e-08, 6.562362e-08, 
    6.508945e-08, 6.481232e-08, 6.47406e-08, 6.460682e-08, 6.474366e-08, 
    6.473253e-08, 6.486347e-08, 6.482139e-08, 6.513578e-08, 6.49669e-08, 
    6.544663e-08, 6.562171e-08, 6.611609e-08, 6.641916e-08, 6.672765e-08, 
    6.686385e-08, 6.690531e-08, 6.692264e-08 ;

 SOILC_LOSS =
  6.359073e-08, 6.38703e-08, 6.381595e-08, 6.404144e-08, 6.391635e-08, 
    6.406401e-08, 6.364741e-08, 6.38814e-08, 6.373202e-08, 6.361589e-08, 
    6.447906e-08, 6.405151e-08, 6.492314e-08, 6.465046e-08, 6.533541e-08, 
    6.488071e-08, 6.542709e-08, 6.532228e-08, 6.563771e-08, 6.554734e-08, 
    6.595081e-08, 6.567942e-08, 6.615994e-08, 6.588599e-08, 6.592885e-08, 
    6.567046e-08, 6.413754e-08, 6.442583e-08, 6.412046e-08, 6.416157e-08, 
    6.414312e-08, 6.391894e-08, 6.380597e-08, 6.356935e-08, 6.36123e-08, 
    6.37861e-08, 6.418006e-08, 6.404632e-08, 6.438335e-08, 6.437574e-08, 
    6.475095e-08, 6.458178e-08, 6.521241e-08, 6.503318e-08, 6.555111e-08, 
    6.542086e-08, 6.5545e-08, 6.550735e-08, 6.554549e-08, 6.535446e-08, 
    6.54363e-08, 6.52682e-08, 6.461346e-08, 6.480589e-08, 6.423198e-08, 
    6.388689e-08, 6.365767e-08, 6.349501e-08, 6.3518e-08, 6.356184e-08, 
    6.378711e-08, 6.39989e-08, 6.41603e-08, 6.426826e-08, 6.437465e-08, 
    6.469666e-08, 6.486707e-08, 6.524866e-08, 6.517979e-08, 6.529645e-08, 
    6.54079e-08, 6.559502e-08, 6.556422e-08, 6.564666e-08, 6.529337e-08, 
    6.552817e-08, 6.514056e-08, 6.524657e-08, 6.440359e-08, 6.408239e-08, 
    6.39459e-08, 6.38264e-08, 6.353569e-08, 6.373644e-08, 6.36573e-08, 
    6.384558e-08, 6.396522e-08, 6.390604e-08, 6.427122e-08, 6.412925e-08, 
    6.487718e-08, 6.455502e-08, 6.53949e-08, 6.519392e-08, 6.544307e-08, 
    6.531594e-08, 6.553378e-08, 6.533772e-08, 6.567733e-08, 6.575129e-08, 
    6.570075e-08, 6.589487e-08, 6.532685e-08, 6.5545e-08, 6.390439e-08, 
    6.391404e-08, 6.395899e-08, 6.376138e-08, 6.374928e-08, 6.356817e-08, 
    6.372932e-08, 6.379795e-08, 6.397214e-08, 6.407519e-08, 6.417314e-08, 
    6.43885e-08, 6.462902e-08, 6.496534e-08, 6.520695e-08, 6.536891e-08, 
    6.52696e-08, 6.535728e-08, 6.525926e-08, 6.521332e-08, 6.572358e-08, 
    6.543706e-08, 6.586696e-08, 6.584317e-08, 6.564862e-08, 6.584585e-08, 
    6.392082e-08, 6.386528e-08, 6.367247e-08, 6.382336e-08, 6.354846e-08, 
    6.370234e-08, 6.379082e-08, 6.413222e-08, 6.420723e-08, 6.427678e-08, 
    6.441415e-08, 6.459044e-08, 6.489969e-08, 6.516876e-08, 6.541438e-08, 
    6.539639e-08, 6.540272e-08, 6.54576e-08, 6.532167e-08, 6.547991e-08, 
    6.550647e-08, 6.543703e-08, 6.583998e-08, 6.572486e-08, 6.584266e-08, 
    6.57677e-08, 6.388333e-08, 6.397677e-08, 6.392628e-08, 6.402123e-08, 
    6.395434e-08, 6.425178e-08, 6.434096e-08, 6.475822e-08, 6.458697e-08, 
    6.485951e-08, 6.461465e-08, 6.465804e-08, 6.486842e-08, 6.462788e-08, 
    6.515393e-08, 6.47973e-08, 6.545973e-08, 6.510361e-08, 6.548205e-08, 
    6.541332e-08, 6.55271e-08, 6.562901e-08, 6.575721e-08, 6.599377e-08, 
    6.593899e-08, 6.613681e-08, 6.411607e-08, 6.423728e-08, 6.42266e-08, 
    6.435343e-08, 6.444724e-08, 6.465053e-08, 6.49766e-08, 6.485399e-08, 
    6.507909e-08, 6.512427e-08, 6.478229e-08, 6.499227e-08, 6.431839e-08, 
    6.442727e-08, 6.436243e-08, 6.412564e-08, 6.488224e-08, 6.449396e-08, 
    6.521095e-08, 6.500061e-08, 6.561448e-08, 6.530919e-08, 6.590884e-08, 
    6.616519e-08, 6.640643e-08, 6.668839e-08, 6.430341e-08, 6.422106e-08, 
    6.436851e-08, 6.457253e-08, 6.47618e-08, 6.501344e-08, 6.503917e-08, 
    6.508632e-08, 6.520843e-08, 6.531109e-08, 6.510123e-08, 6.533683e-08, 
    6.445253e-08, 6.491594e-08, 6.418993e-08, 6.440856e-08, 6.45605e-08, 
    6.449384e-08, 6.483997e-08, 6.492154e-08, 6.525305e-08, 6.508168e-08, 
    6.610193e-08, 6.565055e-08, 6.690304e-08, 6.655304e-08, 6.419229e-08, 
    6.430313e-08, 6.468889e-08, 6.450534e-08, 6.503023e-08, 6.515943e-08, 
    6.526445e-08, 6.539872e-08, 6.541321e-08, 6.549276e-08, 6.53624e-08, 
    6.54876e-08, 6.501397e-08, 6.522563e-08, 6.464479e-08, 6.478616e-08, 
    6.472112e-08, 6.464978e-08, 6.486996e-08, 6.510454e-08, 6.510954e-08, 
    6.518476e-08, 6.539673e-08, 6.503235e-08, 6.61602e-08, 6.546369e-08, 
    6.442399e-08, 6.46375e-08, 6.466798e-08, 6.458527e-08, 6.514647e-08, 
    6.494314e-08, 6.549082e-08, 6.53428e-08, 6.558533e-08, 6.546481e-08, 
    6.544708e-08, 6.529229e-08, 6.519593e-08, 6.495246e-08, 6.475436e-08, 
    6.459727e-08, 6.46338e-08, 6.480636e-08, 6.511888e-08, 6.541453e-08, 
    6.534977e-08, 6.556689e-08, 6.499217e-08, 6.523317e-08, 6.514002e-08, 
    6.538289e-08, 6.485072e-08, 6.530392e-08, 6.473489e-08, 6.478478e-08, 
    6.49391e-08, 6.524952e-08, 6.531818e-08, 6.539152e-08, 6.534626e-08, 
    6.512681e-08, 6.509086e-08, 6.493535e-08, 6.489241e-08, 6.477391e-08, 
    6.467581e-08, 6.476544e-08, 6.485958e-08, 6.51269e-08, 6.536781e-08, 
    6.563047e-08, 6.569473e-08, 6.600164e-08, 6.575182e-08, 6.616408e-08, 
    6.58136e-08, 6.642029e-08, 6.533017e-08, 6.580328e-08, 6.494612e-08, 
    6.503846e-08, 6.520549e-08, 6.558857e-08, 6.538175e-08, 6.562362e-08, 
    6.508945e-08, 6.481232e-08, 6.47406e-08, 6.460682e-08, 6.474366e-08, 
    6.473253e-08, 6.486347e-08, 6.482139e-08, 6.513578e-08, 6.49669e-08, 
    6.544663e-08, 6.562171e-08, 6.611609e-08, 6.641916e-08, 6.672765e-08, 
    6.686385e-08, 6.690531e-08, 6.692264e-08 ;

 SOILICE =
  57.88735, 58.08074, 58.04312, 58.19937, 58.11268, 58.21503, 57.92654, 
    58.0884, 57.98505, 57.90478, 58.50351, 58.20636, 58.81379, 58.62326, 
    59.10293, 58.78407, 59.16741, 59.09379, 59.31577, 59.25211, 59.53662, 
    59.34517, 59.68464, 59.49089, 59.52114, 59.33885, 58.26613, 58.46642, 
    58.25426, 58.28279, 58.27, 58.11444, 58.03613, 57.87264, 57.90231, 
    58.02243, 58.29562, 58.20281, 58.43708, 58.43179, 58.69345, 58.57535, 
    59.01663, 58.89095, 59.25477, 59.16309, 59.25045, 59.22396, 59.25079, 
    59.11639, 59.17394, 59.05581, 58.59744, 58.73183, 58.33173, 58.09213, 
    57.93362, 57.82131, 57.83717, 57.86742, 58.02313, 58.16991, 58.28196, 
    58.357, 58.43103, 58.65538, 58.77457, 59.04203, 58.99376, 59.07561, 
    59.15398, 59.28567, 59.26399, 59.32205, 59.07349, 59.23857, 58.96625, 
    59.04063, 58.45092, 58.22785, 58.13304, 58.05034, 57.84937, 57.98808, 
    57.93336, 58.06366, 58.14655, 58.10556, 58.35905, 58.26038, 58.78164, 
    58.55665, 59.14484, 59.00367, 59.17873, 59.08936, 59.24253, 59.10466, 
    59.34369, 59.39581, 59.36018, 59.49722, 59.09702, 59.25043, 58.1044, 
    58.11108, 58.14225, 58.00532, 57.99697, 57.87181, 57.98319, 58.03065, 
    58.15138, 58.22284, 58.29086, 58.44065, 58.60826, 58.84338, 59.01281, 
    59.12658, 59.05681, 59.1184, 59.04955, 59.0173, 59.37626, 59.17447, 
    59.47749, 59.4607, 59.32342, 59.46259, 58.11578, 58.07732, 57.94387, 
    58.04828, 57.8582, 57.9645, 58.02568, 58.26239, 58.31456, 58.3629, 
    58.45852, 58.58139, 58.79744, 58.98598, 59.15856, 59.1459, 59.15036, 
    59.18893, 59.09338, 59.20464, 59.2233, 59.17447, 59.45845, 59.37721, 
    59.46034, 59.40744, 58.08982, 58.15457, 58.11957, 58.18539, 58.139, 
    58.34546, 58.40747, 58.69846, 58.57896, 58.76931, 58.59829, 58.62855, 
    58.77543, 58.60754, 58.97552, 58.72575, 59.19043, 58.94017, 59.20614, 
    59.15781, 59.23787, 59.30962, 59.40003, 59.56707, 59.52837, 59.66831, 
    58.25124, 58.3354, 58.32803, 58.41624, 58.48154, 58.62334, 58.8513, 
    58.76551, 58.92313, 58.9548, 58.71539, 58.86225, 58.39182, 58.46757, 
    58.42249, 58.25784, 58.7852, 58.51405, 59.0156, 58.86812, 59.29938, 
    59.08455, 59.50706, 59.68829, 59.85947, 60.05975, 58.38143, 58.32419, 
    58.42676, 58.56883, 58.70103, 58.8771, 58.89516, 58.92819, 59.01386, 
    59.08595, 58.93859, 59.10403, 58.48506, 58.80881, 58.30252, 58.45453, 
    58.56047, 58.51402, 58.75572, 58.81279, 59.04513, 58.92496, 59.64348, 
    59.32472, 60.21274, 59.96351, 58.30419, 58.38126, 58.65007, 58.52205, 
    58.88889, 58.97945, 59.0532, 59.1475, 59.15772, 59.21367, 59.12201, 
    59.21006, 58.87748, 59.02592, 58.61935, 58.71807, 58.67265, 58.62283, 
    58.77669, 58.9409, 58.94448, 58.9972, 59.14584, 58.89038, 59.68459, 
    59.19298, 58.46539, 58.61414, 58.63551, 58.57781, 58.97037, 58.82788, 
    59.21231, 59.10823, 59.27886, 59.19402, 59.18154, 59.07274, 59.00507, 
    58.83439, 58.69583, 58.58619, 58.61167, 58.73217, 58.95097, 59.15862, 
    59.11307, 59.26588, 58.86223, 59.03118, 58.96581, 59.13639, 58.76321, 
    59.08066, 58.68227, 58.71712, 58.82505, 59.0426, 59.09093, 59.14244, 
    59.11066, 58.95655, 58.93136, 58.82244, 58.79236, 58.70954, 58.64101, 
    58.7036, 58.76938, 58.95664, 59.12577, 59.31063, 59.35597, 59.5725, 
    59.39609, 59.68732, 59.4395, 59.86908, 59.09921, 59.43237, 58.82999, 
    58.89466, 59.01171, 59.28104, 59.13559, 59.30575, 58.93038, 58.73629, 
    58.68625, 58.59283, 58.68839, 58.68062, 58.77216, 58.74273, 58.96287, 
    58.84454, 59.18121, 59.30443, 59.6536, 59.86841, 60.08781, 60.18483, 
    60.21439, 60.22675,
  78.10485, 78.40597, 78.34741, 78.58918, 78.45574, 78.61291, 78.16592, 
    78.41786, 78.257, 78.13204, 79.04958, 78.59978, 79.52005, 79.23138, 
    79.95847, 79.47494, 80.0563, 79.94473, 80.28149, 80.18491, 80.61639, 
    80.3261, 80.84117, 80.54712, 80.59297, 80.3165, 78.69035, 78.99339, 
    78.67237, 78.71553, 78.69621, 78.45846, 78.33643, 78.08202, 78.1282, 
    78.31516, 78.73495, 78.59448, 78.94936, 78.94134, 79.33776, 79.15882, 
    79.82771, 79.63719, 80.18894, 80.04987, 80.18237, 80.1422, 80.18289, 
    79.979, 80.06629, 79.88715, 79.19226, 79.39589, 78.78968, 78.42358, 
    78.17691, 78.0021, 78.02679, 78.07384, 78.31625, 78.54466, 78.71438, 
    78.82803, 78.94018, 79.27982, 79.46059, 79.86617, 79.79305, 79.9171, 
    80.03605, 80.23579, 80.20291, 80.29096, 79.91398, 80.16429, 79.75138, 
    79.86412, 78.96989, 78.6324, 78.4873, 78.35863, 78.04577, 78.26168, 
    78.17649, 78.37943, 78.50851, 78.44468, 78.83114, 78.68167, 79.47131, 
    79.13041, 80.02216, 79.80807, 80.07358, 79.93805, 80.17032, 79.96126, 
    80.32382, 80.40285, 80.34882, 80.55679, 79.94966, 80.18229, 78.44286, 
    78.45325, 78.50182, 78.28853, 78.27553, 78.08071, 78.2541, 78.32798, 
    78.51604, 78.62481, 78.72782, 78.9547, 79.2086, 79.56497, 79.82193, 
    79.99451, 79.8887, 79.9821, 79.87766, 79.82879, 80.37318, 80.06706, 
    80.52686, 80.50139, 80.29303, 80.50426, 78.46057, 78.4007, 78.19288, 
    78.35548, 78.05953, 78.22499, 78.32021, 78.68462, 78.76375, 78.83692, 
    78.9818, 79.16796, 79.49534, 79.7812, 80.04301, 80.02381, 80.03056, 
    80.08905, 79.94412, 80.11287, 80.14114, 80.06712, 80.49797, 80.3747, 
    80.50084, 80.42059, 78.42018, 78.521, 78.46649, 78.56807, 78.49671, 
    78.8104, 78.90433, 79.34525, 79.16425, 79.45269, 79.19357, 79.23939, 
    79.46178, 79.20761, 79.76527, 79.38655, 80.09132, 79.71157, 80.11515, 
    80.04187, 80.16331, 80.27212, 80.40932, 80.66273, 80.60403, 80.81644, 
    78.66782, 78.79523, 78.78416, 78.91776, 79.01666, 79.23155, 79.57702, 
    79.44702, 79.68599, 79.73398, 79.37106, 79.59358, 78.88071, 78.99538, 
    78.9272, 78.67778, 79.47675, 79.0658, 79.82615, 79.60255, 80.25658, 
    79.93063, 80.57169, 80.84659, 81.1067, 81.41068, 78.86501, 78.77834, 
    78.93371, 79.14882, 79.34927, 79.61614, 79.64358, 79.69362, 79.82356, 
    79.93288, 79.7093, 79.9603, 79.02169, 79.51257, 78.74545, 78.9756, 
    79.13619, 79.06586, 79.43221, 79.5187, 79.87089, 79.68876, 80.77854, 
    80.29491, 81.64324, 81.26456, 78.74803, 78.86478, 79.27197, 79.07804, 
    79.63406, 79.77135, 79.88322, 80.02617, 80.04173, 80.12655, 79.98757, 
    80.12111, 79.61671, 79.84182, 79.22552, 79.37508, 79.3063, 79.2308, 
    79.46399, 79.71278, 79.71835, 79.79822, 80.02322, 79.63634, 80.84068, 
    80.09478, 78.99223, 79.21746, 79.24997, 79.16257, 79.75757, 79.54153, 
    80.12451, 79.96667, 80.22549, 80.09677, 80.07784, 79.91285, 79.8102, 
    79.55138, 79.34137, 79.17528, 79.21389, 79.39643, 79.72808, 80.04302, 
    79.97392, 80.2058, 79.59364, 79.84974, 79.7506, 80.00936, 79.44351, 
    79.92442, 79.32088, 79.3737, 79.53725, 79.86697, 79.94043, 80.01849, 
    79.97036, 79.73656, 79.69841, 79.53333, 79.48768, 79.36221, 79.25835, 
    79.35318, 79.45283, 79.73676, 79.9932, 80.27363, 80.34248, 80.67075, 
    80.40311, 80.8448, 80.46866, 81.12093, 79.95273, 80.45809, 79.54478, 
    79.64283, 79.82017, 80.22861, 80.00815, 80.26614, 79.69694, 79.40262, 
    79.3269, 79.18533, 79.33015, 79.31837, 79.45712, 79.41253, 79.7462, 
    79.56683, 80.07729, 80.26416, 80.79408, 81.12013, 81.45351, 81.60089, 
    81.64581, 81.66459,
  118.4624, 119.0191, 118.9107, 119.3608, 119.111, 119.4059, 118.5752, 
    119.0412, 118.7435, 118.5125, 120.2376, 119.3809, 121.1325, 120.5825, 
    121.9626, 121.0468, 122.1428, 121.9369, 122.5576, 122.3795, 123.1759, 
    122.6398, 123.5903, 123.0477, 123.1325, 122.6222, 119.553, 120.1307, 
    119.5188, 119.601, 119.5641, 119.1161, 118.8908, 118.42, 118.5054, 
    118.8512, 119.638, 119.3705, 120.0456, 120.0303, 120.785, 120.4443, 
    121.718, 121.355, 122.387, 122.1306, 122.3749, 122.3008, 122.3759, 
    122.0001, 122.161, 121.8307, 120.5081, 120.8958, 119.742, 119.0521, 
    118.5956, 118.2723, 118.318, 118.4051, 118.8532, 119.2758, 119.5985, 
    119.8148, 120.0281, 120.6755, 121.0192, 121.7914, 121.6518, 121.8862, 
    122.1052, 122.4734, 122.4128, 122.5752, 121.8802, 122.3417, 121.5724, 
    121.7872, 120.0861, 119.4427, 119.1699, 118.9315, 118.3531, 118.7523, 
    118.5948, 118.9698, 119.2085, 119.0904, 119.8207, 119.5364, 121.0396, 
    120.3905, 122.0796, 121.6805, 122.1743, 121.9245, 122.3528, 121.9673, 
    122.6357, 122.7816, 122.6819, 123.0653, 121.9459, 122.3749, 119.0871, 
    119.1064, 119.1961, 118.802, 118.7779, 118.4177, 118.7382, 118.8749, 
    119.2224, 119.4283, 119.6242, 120.0559, 120.5394, 121.2178, 121.7069, 
    122.0285, 121.8335, 122.0057, 121.813, 121.7198, 122.7269, 122.1625, 
    123.0101, 122.9631, 122.5791, 122.9684, 119.1199, 119.0091, 118.625, 
    118.9255, 118.3785, 118.6844, 118.8606, 119.5423, 119.6925, 119.8318, 
    120.1074, 120.4617, 121.0851, 121.6295, 122.1179, 122.0825, 122.095, 
    122.2029, 121.9357, 122.2468, 122.299, 122.1624, 122.9568, 122.7295, 
    122.9621, 122.8141, 119.0451, 119.2316, 119.1308, 119.3204, 119.1868, 
    119.7817, 119.9605, 120.7996, 120.4547, 121.004, 120.5105, 120.5978, 
    121.0219, 120.5371, 121.5994, 120.8784, 122.2071, 121.4974, 122.251, 
    122.1158, 122.3397, 122.5404, 122.7933, 123.261, 123.1526, 123.5444, 
    119.51, 119.7526, 119.7313, 119.9855, 120.1738, 120.5827, 121.2406, 
    120.9929, 121.4479, 121.5394, 120.8482, 121.2722, 119.9152, 120.1337, 
    120.0036, 119.5291, 121.0499, 120.2677, 121.715, 121.2891, 122.5118, 
    121.9112, 123.0929, 123.6006, 124.08, 124.6418, 119.8852, 119.7202, 
    120.0158, 120.4256, 120.8069, 121.315, 121.3671, 121.4625, 121.7099, 
    121.915, 121.4927, 121.9655, 120.1844, 121.118, 119.6578, 120.0961, 
    120.4015, 120.2675, 120.9646, 121.1293, 121.8004, 121.4531, 123.4752, 
    122.5828, 125.0709, 124.3718, 119.6626, 119.8847, 120.6599, 120.2906, 
    121.349, 121.6106, 121.8234, 122.0871, 122.1156, 122.2721, 122.0157, 
    122.2619, 121.3161, 121.7448, 120.5711, 120.856, 120.7249, 120.5812, 
    121.0251, 121.4994, 121.5095, 121.6619, 122.083, 121.3533, 123.5906, 
    122.2147, 120.1272, 120.5564, 120.6178, 120.4514, 121.5843, 121.1729, 
    122.2683, 121.9772, 122.4544, 122.2171, 122.1822, 121.878, 121.6845, 
    121.1918, 120.7919, 120.4755, 120.549, 120.8968, 121.5284, 122.1182, 
    121.9909, 122.418, 121.2721, 121.76, 121.5713, 122.056, 120.9863, 
    121.9007, 120.7527, 120.8532, 121.1648, 121.7932, 121.9289, 122.0729, 
    121.984, 121.5445, 121.4717, 121.1572, 121.0704, 120.8313, 120.6336, 
    120.8143, 121.0042, 121.5447, 122.0263, 122.5433, 122.6701, 123.2764, 
    122.7826, 123.5983, 122.9044, 124.1074, 121.9523, 122.8842, 121.179, 
    121.3657, 121.7039, 122.4606, 122.0537, 122.5297, 121.4689, 120.9087, 
    120.7642, 120.4947, 120.7703, 120.7479, 121.012, 120.9271, 121.5627, 
    121.221, 122.1813, 122.526, 123.5033, 124.1053, 124.7203, 124.9925, 
    125.0754, 125.1101,
  187.2937, 188.2959, 188.1007, 188.9114, 188.4613, 188.9927, 187.4965, 
    188.3358, 187.7997, 187.3837, 190.4924, 188.9476, 192.1069, 191.1142, 
    193.6134, 191.9522, 193.9387, 193.5668, 194.6876, 194.366, 195.8053, 
    194.8362, 196.5546, 195.5735, 195.7267, 194.8043, 189.2577, 190.2996, 
    189.1961, 189.3443, 189.2778, 188.4707, 188.065, 187.2172, 187.3709, 
    187.9936, 189.4111, 188.9289, 190.1456, 190.1181, 191.4796, 190.8648, 
    193.1642, 192.5085, 194.3794, 193.9166, 194.3577, 194.2238, 194.3594, 
    193.6809, 193.9714, 193.3687, 190.9798, 191.6796, 189.5985, 188.3556, 
    187.5333, 186.9515, 187.0337, 187.1904, 187.9973, 188.7582, 189.3398, 
    189.7295, 190.1141, 191.2822, 191.9025, 193.2971, 193.0448, 193.4723, 
    193.8706, 194.5357, 194.4261, 194.7195, 193.461, 194.2979, 192.9012, 
    193.2894, 190.2191, 189.0589, 188.5676, 188.1382, 187.0969, 187.8156, 
    187.532, 188.2071, 188.637, 188.4243, 189.7402, 189.2278, 191.9393, 
    190.7677, 193.8244, 193.0965, 193.9955, 193.5437, 194.3178, 193.6216, 
    194.8288, 195.0925, 194.9123, 195.6052, 193.5831, 194.3577, 188.4183, 
    188.453, 188.6147, 187.905, 187.8616, 187.213, 187.79, 188.0361, 188.662, 
    189.0329, 189.3861, 190.1643, 191.0364, 192.2609, 193.1442, 193.7322, 
    193.3738, 193.6909, 193.3359, 193.1676, 194.9937, 193.9741, 195.5054, 
    195.4205, 194.7265, 195.43, 188.4774, 188.2778, 187.5863, 188.1273, 
    187.1425, 187.6933, 188.0106, 189.2385, 189.5091, 189.7603, 190.2571, 
    190.8962, 192.0214, 193.0044, 193.8936, 193.8297, 193.8522, 194.047, 
    193.5647, 194.1263, 194.2207, 193.974, 195.4091, 194.9982, 195.4186, 
    195.151, 188.3427, 188.6786, 188.497, 188.8386, 188.5979, 189.67, 
    189.9923, 191.5061, 190.8837, 191.8749, 190.9841, 191.1418, 191.9074, 
    191.0322, 192.9502, 191.6483, 194.0546, 192.7661, 194.1339, 193.8898, 
    194.2941, 194.6567, 195.1136, 195.959, 195.763, 196.4716, 189.1803, 
    189.6176, 189.579, 190.0374, 190.377, 191.1145, 192.302, 191.8547, 
    192.6763, 192.8416, 191.5936, 192.3592, 189.9107, 190.3047, 190.07, 
    189.2148, 191.9578, 190.5463, 193.1589, 192.3896, 194.6049, 193.519, 
    195.6552, 196.5735, 197.4406, 198.4581, 189.8565, 189.559, 190.0919, 
    190.8313, 191.5191, 192.4364, 192.5305, 192.7028, 193.1496, 193.5259, 
    192.7573, 193.6184, 190.3963, 192.0807, 189.4467, 190.237, 190.7876, 
    190.5459, 191.8036, 192.101, 193.3132, 192.6858, 196.3466, 194.7334, 
    199.2354, 197.9692, 189.4552, 189.8555, 191.2539, 190.5875, 192.4978, 
    192.9702, 193.3549, 193.838, 193.8894, 194.172, 193.7091, 194.1537, 
    192.4384, 193.2126, 191.0936, 191.6077, 191.3711, 191.1117, 191.9129, 
    192.7694, 192.7877, 193.063, 193.8311, 192.5056, 196.5557, 194.0688, 
    190.2928, 191.0672, 191.1779, 190.8775, 192.9228, 192.1798, 194.1651, 
    193.6396, 194.5012, 194.0727, 194.0097, 193.457, 193.1039, 192.2139, 
    191.492, 190.921, 191.0537, 191.6813, 192.8219, 193.8941, 193.6643, 
    194.4356, 192.3588, 193.2403, 192.8992, 193.7818, 191.8429, 193.4998, 
    191.4211, 191.6027, 192.1651, 193.3002, 193.552, 193.8124, 193.6519, 
    192.8509, 192.7194, 192.1514, 191.9948, 191.5631, 191.2063, 191.5323, 
    191.8752, 192.8512, 193.7283, 194.6619, 194.8908, 195.9873, 195.0945, 
    196.5696, 195.315, 197.4907, 193.5949, 195.2781, 192.1907, 192.5278, 
    193.1389, 194.5127, 193.7778, 194.6375, 192.7142, 191.703, 191.4419, 
    190.9557, 191.453, 191.4126, 191.8893, 191.736, 192.8837, 192.2665, 
    194.0081, 194.6307, 196.3973, 197.4865, 198.6001, 199.0933, 199.2436, 
    199.3065,
  314.8134, 316.5515, 316.2129, 317.6201, 316.8387, 317.7612, 315.165, 
    316.6208, 315.6907, 314.9695, 320.3683, 317.683, 323.18, 321.4506, 
    325.8119, 322.9104, 326.3999, 325.7276, 327.7547, 327.1727, 329.768, 
    328.0236, 331.0811, 329.3589, 329.6304, 327.9659, 318.2215, 320.0329, 
    318.1145, 318.3721, 318.2565, 316.8549, 316.1509, 314.6809, 314.9472, 
    316.0271, 318.488, 317.6505, 319.765, 319.7171, 322.0868, 321.0163, 
    325.0244, 323.8803, 327.197, 326.3598, 327.1576, 326.9155, 327.1608, 
    325.9338, 326.459, 325.3813, 321.2166, 322.4352, 318.8137, 316.6552, 
    315.2288, 314.2204, 314.3628, 314.6344, 316.0334, 317.3541, 318.3641, 
    319.0414, 319.7102, 321.7431, 322.8237, 325.2563, 324.8159, 325.5623, 
    326.2766, 327.4796, 327.2813, 327.8124, 325.5424, 327.0494, 324.5653, 
    325.2429, 319.8928, 317.8762, 317.0232, 316.278, 314.4723, 315.7182, 
    315.2265, 316.3974, 317.1436, 316.7743, 319.06, 318.1696, 322.8879, 
    320.8474, 326.1932, 324.9062, 326.5024, 325.687, 327.0855, 325.8265, 
    328.0102, 328.4877, 328.1613, 329.4164, 325.7569, 327.1577, 316.764, 
    316.8242, 317.1048, 315.8733, 315.7981, 314.6736, 315.6739, 316.1009, 
    317.1869, 317.8311, 318.4446, 319.7975, 321.315, 323.4485, 324.9895, 
    326.0265, 325.3902, 325.9519, 325.3241, 325.0302, 328.3087, 326.4639, 
    329.2356, 329.0816, 327.8251, 329.0989, 316.8665, 316.5202, 315.3207, 
    316.259, 314.5514, 315.5062, 316.0565, 318.1883, 318.6583, 319.095, 
    319.9589, 321.071, 323.0309, 324.7455, 326.3182, 326.2027, 326.2434, 
    326.5957, 325.7237, 326.7391, 326.9099, 326.4636, 329.061, 328.3169, 
    329.0783, 328.5936, 316.6327, 317.2158, 316.9006, 317.4937, 317.0758, 
    318.938, 319.4984, 322.133, 321.0491, 322.7756, 321.224, 321.4985, 
    322.8324, 321.3076, 324.6508, 322.3809, 326.6094, 324.3297, 326.7528, 
    326.3114, 327.0425, 327.6987, 328.5258, 330.0373, 329.6938, 330.9356, 
    318.087, 318.847, 318.7798, 319.5768, 320.1674, 321.4509, 323.5201, 
    322.7404, 324.173, 324.4613, 322.2854, 323.6198, 319.3564, 320.0417, 
    319.6334, 318.1469, 322.9201, 320.462, 325.015, 323.6729, 327.605, 
    325.6439, 329.5049, 331.1143, 332.6356, 334.423, 319.2623, 318.7451, 
    319.6716, 320.9579, 322.1556, 323.7546, 323.9186, 324.2191, 324.9989, 
    325.6559, 324.3144, 325.8208, 320.201, 323.1342, 318.5499, 319.9239, 
    320.8819, 320.4612, 322.6514, 323.1698, 325.2844, 324.1895, 330.7165, 
    327.8376, 335.7901, 333.5638, 318.5646, 319.2605, 321.6937, 320.5338, 
    323.8615, 324.6858, 325.3573, 326.2178, 326.3107, 326.8217, 325.9848, 
    326.7885, 323.758, 325.1089, 321.4146, 322.3101, 321.8978, 321.4462, 
    322.8419, 324.3355, 324.3673, 324.8477, 326.2055, 323.8751, 331.0832, 
    326.6353, 320.0209, 321.3686, 321.5613, 321.0384, 324.6031, 323.3071, 
    326.8092, 325.8591, 327.4172, 326.6421, 326.5282, 325.5355, 324.919, 
    323.3665, 322.1084, 321.1141, 321.3451, 322.4382, 324.427, 326.3192, 
    325.9038, 327.2985, 323.6191, 325.1572, 324.562, 326.1162, 322.7198, 
    325.6104, 321.985, 322.3012, 323.2814, 325.2619, 325.7014, 326.1715, 
    325.8813, 324.4776, 324.2481, 323.2575, 322.9846, 322.2323, 321.6109, 
    322.1787, 322.7761, 324.4781, 326.0195, 327.708, 328.1225, 330.0868, 
    328.4913, 331.1076, 328.8909, 332.7236, 325.7784, 328.8239, 323.326, 
    323.914, 324.9803, 327.4382, 326.1089, 327.664, 324.2391, 322.4761, 
    322.0212, 321.1745, 322.0406, 321.97, 322.8007, 322.5335, 324.5348, 
    323.4583, 326.5254, 327.6516, 330.8053, 332.7162, 334.6725, 335.54, 
    335.8045, 335.9151,
  523.2206, 526.4933, 525.8551, 528.5091, 527.0347, 528.7756, 523.882, 
    526.6239, 524.8715, 523.514, 533.7067, 528.6279, 539.0443, 535.7587, 
    544.0591, 538.5316, 545.1821, 543.8983, 547.7728, 546.6593, 551.6535, 
    548.2877, 554.2643, 550.8472, 551.3801, 548.1772, 529.6448, 533.0712, 
    529.4427, 529.9295, 529.7109, 527.0652, 525.7383, 522.9713, 523.4723, 
    525.5051, 530.1485, 528.5665, 532.564, 532.4733, 536.9666, 534.9349, 
    542.5568, 540.3768, 546.7057, 545.1055, 546.6305, 546.1675, 546.6365, 
    544.292, 545.295, 543.2374, 535.3148, 537.6284, 530.7642, 526.6887, 
    524.002, 522.1057, 522.3732, 522.8839, 525.517, 528.007, 529.9143, 
    531.1948, 532.4603, 536.314, 538.3668, 542.9991, 542.1591, 543.5827, 
    544.9467, 547.2465, 546.8671, 547.8834, 543.5449, 546.4236, 541.6815, 
    542.9734, 532.8061, 528.9927, 527.3828, 525.9778, 522.5791, 524.9234, 
    523.9977, 526.2028, 527.61, 526.9134, 531.2299, 529.5468, 538.4888, 
    534.6146, 544.7874, 542.3314, 545.378, 543.8207, 546.4926, 544.0872, 
    548.2621, 549.1767, 548.5515, 550.9574, 543.9542, 546.6306, 526.894, 
    527.0075, 527.5367, 525.2154, 525.0737, 522.9576, 524.8399, 525.644, 
    527.6916, 528.9075, 530.0664, 532.6254, 535.5015, 539.5549, 542.4902, 
    544.4689, 543.2544, 544.3265, 543.1283, 542.5677, 548.8339, 545.3044, 
    550.6105, 550.3152, 547.9077, 550.3484, 527.0872, 526.4342, 524.175, 
    525.942, 522.7278, 524.5242, 525.5605, 529.5821, 530.4704, 531.2961, 
    532.9311, 535.0387, 538.7607, 542.0249, 545.0261, 544.8054, 544.8831, 
    545.5563, 543.8909, 545.8303, 546.1567, 545.3039, 550.2757, 548.8495, 
    550.3089, 549.3797, 526.6464, 527.7462, 527.1516, 528.2704, 527.4819, 
    530.9993, 532.0594, 537.0543, 534.9971, 538.2753, 535.3289, 535.8496, 
    538.3832, 535.4875, 541.8445, 537.5251, 545.5825, 541.2326, 545.8565, 
    545.0131, 546.4103, 547.6656, 549.2498, 552.1884, 551.5061, 553.9747, 
    529.3908, 530.827, 530.7001, 532.2076, 533.3259, 535.7594, 539.6912, 
    538.2084, 540.9341, 541.4835, 537.3438, 539.881, 531.7907, 533.0879, 
    532.3149, 529.5041, 538.5499, 533.8843, 542.5389, 539.9819, 547.4865, 
    543.7385, 551.131, 554.3303, 557.2732, 560.724, 531.6126, 530.6345, 
    532.3872, 534.8243, 537.0971, 540.1375, 540.4496, 541.0221, 542.5081, 
    543.7615, 541.2035, 544.0762, 533.3898, 538.9572, 530.2654, 532.8649, 
    534.6801, 533.8827, 538.0392, 539.0247, 543.0526, 540.9657, 553.5388, 
    547.9316, 563.3696, 559.064, 530.2933, 531.6091, 536.2202, 534.0201, 
    540.3411, 541.9113, 543.1916, 544.8342, 545.0117, 545.9882, 544.3892, 
    545.9248, 540.144, 542.7179, 535.6904, 537.3906, 536.6075, 535.7504, 
    538.4013, 541.2437, 541.3043, 542.2198, 544.8107, 540.3669, 554.2684, 
    545.6319, 533.0485, 535.6032, 535.9689, 534.9767, 541.7536, 539.2859, 
    545.9643, 544.1492, 547.127, 545.6448, 545.4272, 543.5317, 542.3558, 
    539.3989, 537.0076, 535.1205, 535.5585, 537.634, 541.4181, 545.028, 
    544.2347, 546.9, 539.8797, 542.8099, 541.6752, 544.6401, 538.1691, 
    543.6746, 536.7731, 537.3738, 539.2371, 543.0096, 543.8481, 544.7459, 
    544.1917, 541.5145, 541.0773, 539.1917, 538.6727, 537.2429, 536.0629, 
    537.141, 538.2761, 541.5154, 544.4556, 547.6836, 548.4771, 552.2869, 
    549.1835, 554.3171, 549.9496, 557.4429, 543.9952, 549.821, 539.322, 
    540.441, 542.4726, 547.1673, 544.6262, 547.5993, 541.0601, 537.706, 
    536.8419, 535.235, 536.8787, 536.7448, 538.3229, 537.8151, 541.6234, 
    539.5737, 545.4218, 547.5757, 553.7155, 557.4286, 561.2064, 562.8851, 
    563.3974, 563.6118,
  947.1248, 953.9976, 952.6545, 958.2484, 955.1379, 958.8113, 948.5109, 
    954.2725, 950.5872, 947.7395, 969.1224, 958.4991, 980.1622, 973.3553, 
    990.6236, 979.0976, 992.9783, 990.2868, 998.4278, 996.0826, 1006.636, 
    999.5137, 1012.19, 1004.926, 1006.056, 999.2805, 960.6494, 967.8145, 
    960.2218, 961.2517, 960.7892, 955.2023, 952.4089, 946.6025, 947.6519, 
    951.9185, 961.7155, 958.3695, 966.7713, 966.5849, 975.8534, 971.6542, 
    987.4803, 982.9336, 996.1803, 992.8176, 996.022, 995.0482, 996.0347, 
    991.1115, 993.2153, 988.9034, 972.4383, 977.2244, 963.0198, 954.4091, 
    948.7624, 944.7913, 945.3509, 946.4196, 951.9435, 957.1883, 961.2195, 
    963.933, 966.5581, 974.5031, 978.7556, 988.4049, 986.6498, 989.626, 
    992.4842, 997.3187, 996.5198, 998.6609, 989.5468, 995.5867, 985.6528, 
    988.3514, 967.2691, 959.27, 955.8716, 952.9125, 945.7817, 950.6962, 
    948.7536, 953.3861, 956.3506, 954.8823, 964.0074, 960.4417, 979.0087, 
    970.9935, 992.15, 987.0095, 993.3895, 990.1241, 995.7318, 990.6823, 
    999.4597, 1001.391, 1000.07, 1005.16, 990.4038, 996.0222, 954.8413, 
    955.0805, 956.196, 951.3096, 951.012, 946.5739, 950.5209, 952.2106, 
    956.5228, 959.0901, 961.5416, 966.8977, 972.8239, 981.2234, 987.3412, 
    991.4822, 988.939, 991.1837, 988.6751, 987.5033, 1000.667, 993.235, 
    1004.425, 1003.799, 998.712, 1003.87, 955.2485, 953.8731, 949.1253, 
    952.8373, 946.0928, 949.858, 952.0351, 960.5165, 962.3972, 964.1478, 
    967.5262, 971.8683, 979.5732, 986.3696, 992.6508, 992.188, 992.3509, 
    993.7639, 990.2712, 994.3394, 995.0256, 993.2339, 1003.715, 1000.7, 
    1003.786, 1001.82, 954.3198, 956.6379, 955.384, 957.7443, 956.0806, 
    963.5183, 965.7346, 976.035, 971.7827, 978.5659, 972.4675, 973.5432, 
    978.7897, 972.7952, 985.993, 977.0103, 993.8188, 984.7166, 994.3945, 
    992.6235, 995.5588, 998.2018, 1001.545, 1007.772, 1006.323, 1011.572, 
    960.1119, 963.153, 962.8842, 966.0391, 968.3386, 973.3566, 981.5068, 
    978.427, 984.0943, 985.2396, 976.6346, 981.9017, 965.1827, 967.8488, 
    966.2595, 960.3514, 979.1357, 969.4882, 987.443, 982.1116, 997.8243, 
    989.9521, 1005.528, 1012.33, 1018.811, 1026.49, 964.8172, 962.7449, 
    966.408, 971.426, 976.1237, 982.4354, 983.0851, 984.2776, 987.3785, 
    990.0002, 984.6558, 990.6594, 968.4699, 979.9814, 961.9631, 967.39, 
    971.1287, 969.4849, 978.076, 980.1216, 988.5169, 984.1601, 1010.644, 
    998.7625, 1032.29, 1022.79, 962.0221, 964.8101, 974.3091, 969.7681, 
    982.8592, 986.1322, 988.8076, 992.2482, 992.6207, 994.6713, 991.3152, 
    994.5381, 982.4489, 987.817, 973.2141, 976.7316, 975.1104, 973.3381, 
    978.8272, 984.7396, 984.8658, 986.7764, 992.1991, 982.9128, 1012.198, 
    993.9227, 967.7677, 973.034, 973.7896, 971.7406, 985.8032, 980.6644, 
    994.6211, 990.8124, 997.0671, 993.9498, 993.4928, 989.5191, 987.0604, 
    980.8991, 975.9384, 972.0372, 972.9417, 977.236, 985.1032, 992.6548, 
    990.9914, 996.5891, 981.899, 988.0095, 985.6396, 991.8413, 978.3456, 
    989.8184, 975.4529, 976.6968, 980.5629, 988.4271, 990.1817, 992.0631, 
    990.9012, 985.3043, 984.3926, 980.4684, 979.3905, 976.4257, 973.984, 
    976.2146, 978.5675, 985.3063, 991.4543, 998.2397, 999.9133, 1007.981, 
    1001.405, 1012.302, 1003.025, 1019.188, 990.4897, 1002.753, 980.7393, 
    983.067, 987.3044, 997.152, 991.812, 998.0621, 984.3569, 977.3852, 
    975.5953, 972.2737, 975.6715, 975.3943, 978.6646, 977.6115, 985.5316, 
    981.2624, 993.4815, 998.0122, 1011.02, 1019.156, 1027.567, 1031.239, 
    1032.35, 1032.816,
  1829.886, 1849.348, 1845.52, 1861.544, 1852.608, 1863.169, 1833.786, 
    1850.133, 1839.651, 1831.614, 1893.766, 1862.268, 1928.089, 1906.809, 
    1960.685, 1924.735, 1968.115, 1959.626, 1985.501, 1977.986, 2012.206, 
    1988.998, 2030.642, 2006.59, 2010.298, 1988.246, 1868.489, 1889.765, 
    1867.249, 1870.237, 1868.894, 1852.792, 1844.821, 1828.42, 1831.368, 
    1843.427, 1871.585, 1861.894, 1886.584, 1886.016, 1914.574, 1901.55, 
    1950.842, 1936.753, 1978.298, 1967.606, 1977.792, 1974.687, 1977.833, 
    1962.22, 1968.865, 1955.288, 1903.971, 1918.857, 1875.385, 1850.523, 
    1834.495, 1823.349, 1824.913, 1827.906, 1843.498, 1858.491, 1870.144, 
    1878.052, 1885.935, 1910.37, 1923.66, 1953.728, 1948.255, 1957.552, 
    1966.552, 1981.941, 1979.383, 1986.251, 1957.303, 1976.403, 1945.158, 
    1953.561, 1888.101, 1864.494, 1854.71, 1846.254, 1826.119, 1839.96, 
    1834.47, 1847.603, 1856.084, 1851.876, 1878.27, 1867.887, 1924.456, 
    1899.514, 1965.496, 1949.375, 1969.418, 1959.115, 1976.866, 1960.869, 
    1988.824, 1995.068, 1990.795, 2007.356, 1959.994, 1977.793, 1851.759, 
    1852.443, 1855.64, 1841.699, 1840.855, 1828.339, 1839.463, 1844.257, 
    1856.578, 1863.974, 1871.08, 1886.969, 1905.163, 1931.442, 1950.408, 
    1963.389, 1955.399, 1962.448, 1954.573, 1950.913, 1992.722, 1968.928, 
    2004.949, 2002.904, 1986.415, 2003.134, 1852.924, 1848.992, 1835.518, 
    1846.04, 1826.99, 1837.588, 1843.758, 1868.104, 1873.57, 1878.68, 
    1888.885, 1902.211, 1926.232, 1947.384, 1967.079, 1965.616, 1966.13, 
    1970.605, 1959.577, 1972.432, 1974.615, 1968.924, 2002.631, 1992.829, 
    2002.861, 1996.46, 1850.268, 1856.909, 1853.312, 1860.092, 1855.309, 
    1876.84, 1883.43, 1915.141, 1901.946, 1923.064, 1904.062, 1907.391, 
    1923.767, 1905.075, 1946.214, 1918.187, 1970.779, 1942.257, 1972.608, 
    1966.992, 1976.314, 1984.775, 1995.569, 2015.952, 2011.177, 2028.578, 
    1866.931, 1875.773, 1874.989, 1884.356, 1891.367, 1906.813, 1932.338, 
    1922.628, 1940.333, 1943.877, 1917.013, 1933.58, 1881.755, 1889.87, 
    1885.026, 1867.625, 1924.855, 1894.888, 1950.725, 1934.225, 1983.562, 
    1958.575, 2008.563, 2031.113, 2053.029, 2079.234, 1880.647, 1874.583, 
    1885.478, 1900.846, 1915.417, 1935.22, 1937.22, 1940.9, 1950.524, 
    1958.726, 1942.069, 1960.797, 1891.769, 1927.519, 1872.306, 1888.469, 
    1899.93, 1894.878, 1921.526, 1927.961, 1954.078, 1940.536, 2025.48, 
    1986.578, 2099.502, 2066.699, 1872.477, 1880.625, 1909.768, 1895.747, 
    1936.524, 1946.646, 1954.988, 1965.806, 1966.983, 1973.488, 1962.862, 
    1973.064, 1935.261, 1951.892, 1906.371, 1917.316, 1912.259, 1906.755, 
    1923.885, 1942.328, 1942.719, 1948.649, 1965.651, 1936.689, 2030.672, 
    1971.109, 1889.623, 1905.814, 1908.155, 1901.817, 1945.625, 1929.674, 
    1973.328, 1961.279, 1981.135, 1971.195, 1969.745, 1957.216, 1949.533, 
    1930.416, 1914.839, 1902.732, 1905.528, 1918.894, 1943.454, 1967.091, 
    1961.842, 1979.605, 1933.571, 1952.493, 1945.117, 1964.521, 1922.372, 
    1958.155, 1913.326, 1917.207, 1929.354, 1953.797, 1959.296, 1965.221, 
    1961.558, 1944.077, 1941.255, 1929.055, 1925.657, 1916.36, 1908.758, 
    1915.701, 1923.069, 1944.083, 1963.301, 1984.896, 1990.287, 2016.644, 
    1995.115, 2031.019, 2000.38, 2054.315, 1960.264, 1999.495, 1929.911, 
    1937.164, 1950.293, 1981.406, 1964.429, 1984.326, 1941.145, 1919.361, 
    1913.769, 1903.462, 1914.007, 1913.143, 1923.374, 1920.069, 1944.782, 
    1931.565, 1969.709, 1984.166, 2026.734, 2054.207, 2082.894, 2095.755, 
    2099.718, 2101.382,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.547428, 4.565945, 4.562341, 4.577308, 4.569, 4.578807, 4.551177, 
    4.566682, 4.556779, 4.549091, 4.606452, 4.577976, 4.63615, 4.617896, 
    4.66384, 4.633307, 4.670012, 4.662955, 4.684212, 4.678115, 4.705379, 
    4.687027, 4.71955, 4.700991, 4.703892, 4.686423, 4.583694, 4.602901, 
    4.582559, 4.585294, 4.584066, 4.569172, 4.561681, 4.546013, 4.548854, 
    4.560363, 4.586524, 4.57763, 4.600062, 4.599555, 4.624617, 4.613306, 
    4.655566, 4.643528, 4.67837, 4.669591, 4.677958, 4.675419, 4.67799, 
    4.66512, 4.670632, 4.659317, 4.615423, 4.628294, 4.589979, 4.567049, 
    4.551857, 4.541099, 4.542619, 4.545517, 4.56043, 4.57448, 4.585208, 
    4.592394, 4.599482, 4.620988, 4.632393, 4.658004, 4.653373, 4.661218, 
    4.668718, 4.681332, 4.679254, 4.684817, 4.66101, 4.676824, 4.650737, 
    4.657862, 4.601418, 4.580028, 4.570964, 4.563034, 4.543788, 4.557073, 
    4.551833, 4.564305, 4.572243, 4.568316, 4.592591, 4.583143, 4.63307, 
    4.611519, 4.667843, 4.654323, 4.671087, 4.662528, 4.677202, 4.663993, 
    4.686888, 4.691884, 4.688469, 4.701591, 4.663262, 4.677958, 4.568206, 
    4.568846, 4.57183, 4.558725, 4.557923, 4.545936, 4.556601, 4.561148, 
    4.572703, 4.579549, 4.586062, 4.600407, 4.616464, 4.638978, 4.655199, 
    4.666093, 4.65941, 4.66531, 4.658715, 4.655626, 4.690012, 4.670684, 
    4.699702, 4.698093, 4.684949, 4.698274, 4.569296, 4.565611, 4.552837, 
    4.562832, 4.544631, 4.554814, 4.560677, 4.583342, 4.58833, 4.592962, 
    4.602116, 4.613884, 4.634578, 4.652633, 4.669155, 4.667943, 4.668369, 
    4.672066, 4.662914, 4.67357, 4.67536, 4.670681, 4.697877, 4.690097, 
    4.698059, 4.692991, 4.566809, 4.57301, 4.569659, 4.575963, 4.571522, 
    4.591298, 4.597239, 4.625105, 4.613653, 4.631886, 4.615502, 4.618402, 
    4.632485, 4.616386, 4.651638, 4.627721, 4.67221, 4.648259, 4.673714, 
    4.669083, 4.676751, 4.683626, 4.692283, 4.708287, 4.704577, 4.71798, 
    4.582267, 4.590332, 4.58962, 4.598068, 4.604323, 4.6179, 4.639733, 
    4.631514, 4.646609, 4.649643, 4.626713, 4.640784, 4.595733, 4.602993, 
    4.598669, 4.582903, 4.63341, 4.607443, 4.655468, 4.641343, 4.682645, 
    4.662076, 4.702536, 4.719908, 4.736288, 4.755486, 4.594736, 4.589251, 
    4.599073, 4.612689, 4.625342, 4.642204, 4.64393, 4.647095, 4.655297, 
    4.662201, 4.648098, 4.663933, 4.604681, 4.635667, 4.58718, 4.601746, 
    4.611885, 4.607434, 4.630575, 4.636041, 4.658299, 4.646783, 4.715618, 
    4.685081, 4.770131, 4.746264, 4.587337, 4.594716, 4.620466, 4.608202, 
    4.64333, 4.652005, 4.659064, 4.668101, 4.669076, 4.674436, 4.665655, 
    4.674088, 4.64224, 4.656454, 4.617516, 4.626973, 4.62262, 4.61785, 
    4.632584, 4.64832, 4.648654, 4.653708, 4.667973, 4.643473, 4.719573, 
    4.672482, 4.602773, 4.617031, 4.619067, 4.613539, 4.651135, 4.637489, 
    4.674305, 4.664335, 4.680677, 4.672552, 4.671358, 4.660937, 4.654458, 
    4.638114, 4.624845, 4.61434, 4.616781, 4.628325, 4.649282, 4.669165, 
    4.664805, 4.679434, 4.640777, 4.656961, 4.650702, 4.667034, 4.631296, 
    4.661725, 4.623541, 4.62688, 4.637218, 4.658062, 4.662679, 4.667616, 
    4.664568, 4.649815, 4.6474, 4.636966, 4.634089, 4.626153, 4.61959, 
    4.625587, 4.63189, 4.64982, 4.66602, 4.683724, 4.688062, 4.708823, 
    4.691922, 4.719837, 4.696102, 4.737236, 4.663489, 4.6954, 4.637688, 
    4.643882, 4.655102, 4.680898, 4.666957, 4.683263, 4.647305, 4.628726, 
    4.623924, 4.614978, 4.624128, 4.623384, 4.63215, 4.629331, 4.650416, 
    4.639082, 4.671328, 4.683133, 4.716576, 4.737155, 4.75816, 4.767454, 
    4.770285, 4.771469,
  5.633276, 5.65656, 5.652027, 5.670849, 5.660401, 5.672735, 5.63799, 
    5.657486, 5.645034, 5.635367, 5.707512, 5.67169, 5.744887, 5.721914, 
    5.779748, 5.74131, 5.787521, 5.778634, 5.805405, 5.797727, 5.832071, 
    5.808951, 5.849926, 5.826542, 5.830197, 5.80819, 5.678883, 5.703044, 
    5.677454, 5.680894, 5.67935, 5.660618, 5.651197, 5.631497, 5.63507, 
    5.649539, 5.682442, 5.671255, 5.699474, 5.698835, 5.730371, 5.716137, 
    5.769331, 5.754175, 5.798047, 5.786991, 5.797527, 5.794331, 5.797569, 
    5.781361, 5.788301, 5.774053, 5.718801, 5.735, 5.686788, 5.657947, 
    5.638844, 5.625319, 5.62723, 5.630874, 5.649624, 5.667294, 5.680787, 
    5.689826, 5.698743, 5.725804, 5.740159, 5.7724, 5.766569, 5.776447, 
    5.785892, 5.801777, 5.79916, 5.806167, 5.776185, 5.796099, 5.763251, 
    5.772222, 5.701179, 5.674271, 5.66287, 5.652898, 5.6287, 5.645403, 
    5.638814, 5.654497, 5.66448, 5.659541, 5.690074, 5.678189, 5.741011, 
    5.713889, 5.78479, 5.767766, 5.788876, 5.778096, 5.796576, 5.779942, 
    5.808775, 5.815069, 5.810768, 5.827298, 5.779021, 5.797528, 5.659403, 
    5.660208, 5.66396, 5.64748, 5.646472, 5.6314, 5.644809, 5.650527, 
    5.665059, 5.673669, 5.681862, 5.699906, 5.720111, 5.748448, 5.768868, 
    5.782586, 5.774171, 5.7816, 5.773296, 5.769406, 5.812711, 5.788367, 
    5.824918, 5.822891, 5.806334, 5.82312, 5.660774, 5.65614, 5.640076, 
    5.652645, 5.62976, 5.642562, 5.649934, 5.67844, 5.684714, 5.69054, 
    5.702058, 5.716865, 5.742908, 5.765637, 5.786441, 5.784915, 5.785452, 
    5.790108, 5.778583, 5.792001, 5.794257, 5.788363, 5.82262, 5.812818, 
    5.822848, 5.816464, 5.657646, 5.665445, 5.66123, 5.669159, 5.663573, 
    5.688447, 5.695921, 5.730985, 5.716573, 5.73952, 5.718901, 5.722551, 
    5.740273, 5.720013, 5.764384, 5.734278, 5.790289, 5.76013, 5.792183, 
    5.786351, 5.796008, 5.804667, 5.815571, 5.835734, 5.83106, 5.847949, 
    5.677087, 5.687232, 5.686337, 5.696965, 5.704835, 5.721918, 5.749398, 
    5.739052, 5.758053, 5.761874, 5.73301, 5.750721, 5.694027, 5.703161, 
    5.697721, 5.677888, 5.741437, 5.70876, 5.769207, 5.751424, 5.803432, 
    5.777527, 5.828489, 5.850378, 5.871023, 5.895224, 5.692772, 5.685873, 
    5.698229, 5.715361, 5.731285, 5.752508, 5.754682, 5.758666, 5.768992, 
    5.777686, 5.759927, 5.779866, 5.705284, 5.74428, 5.683268, 5.701591, 
    5.714349, 5.708748, 5.737871, 5.74475, 5.772771, 5.758273, 5.844971, 
    5.806499, 5.913692, 5.883598, 5.683464, 5.692748, 5.725147, 5.709714, 
    5.753926, 5.764847, 5.773735, 5.785114, 5.786342, 5.793092, 5.782034, 
    5.792655, 5.752553, 5.770449, 5.721435, 5.733337, 5.727859, 5.721855, 
    5.740399, 5.760207, 5.760628, 5.766991, 5.784953, 5.754106, 5.849956, 
    5.790631, 5.702884, 5.720824, 5.723386, 5.71643, 5.763752, 5.746573, 
    5.792927, 5.780372, 5.800953, 5.79072, 5.789216, 5.776093, 5.767935, 
    5.74736, 5.730659, 5.717438, 5.72051, 5.735039, 5.76142, 5.786455, 
    5.780964, 5.799387, 5.750712, 5.771088, 5.763207, 5.783771, 5.738779, 
    5.777085, 5.729018, 5.73322, 5.746233, 5.772474, 5.778286, 5.784503, 
    5.780666, 5.76209, 5.759049, 5.745915, 5.742294, 5.732305, 5.724045, 
    5.731592, 5.739525, 5.762096, 5.782494, 5.80479, 5.810255, 5.836409, 
    5.815116, 5.850287, 5.820382, 5.872217, 5.779306, 5.819498, 5.746824, 
    5.754621, 5.768746, 5.801231, 5.783674, 5.80421, 5.75893, 5.735542, 
    5.729499, 5.718242, 5.729757, 5.728819, 5.739852, 5.736305, 5.762847, 
    5.748579, 5.789178, 5.804047, 5.846179, 5.872116, 5.898597, 5.910316, 
    5.913886, 5.915379,
  8.097939, 8.132139, 8.125481, 8.153135, 8.137784, 8.155907, 8.104861, 
    8.133501, 8.115208, 8.10101, 8.207026, 8.15437, 8.261999, 8.228205, 
    8.313304, 8.256735, 8.324747, 8.311664, 8.351082, 8.339774, 8.390363, 
    8.356305, 8.416677, 8.382217, 8.387602, 8.355184, 8.164942, 8.200458, 
    8.162842, 8.167897, 8.165628, 8.138102, 8.124262, 8.095326, 8.100573, 
    8.121826, 8.170172, 8.153732, 8.195209, 8.19427, 8.240644, 8.219709, 
    8.297969, 8.275664, 8.340245, 8.323967, 8.33948, 8.334774, 8.339542, 
    8.315678, 8.325896, 8.30492, 8.223627, 8.247453, 8.17656, 8.134177, 
    8.106116, 8.086254, 8.08906, 8.094411, 8.121951, 8.14791, 8.16774, 
    8.181026, 8.194135, 8.233927, 8.255042, 8.302486, 8.293904, 8.308444, 
    8.322349, 8.345739, 8.341885, 8.352203, 8.308058, 8.337378, 8.289021, 
    8.302225, 8.197715, 8.158164, 8.141411, 8.12676, 8.091218, 8.11575, 
    8.106072, 8.129109, 8.143777, 8.136519, 8.18139, 8.163922, 8.256295, 
    8.216404, 8.320725, 8.295665, 8.326741, 8.310871, 8.338078, 8.313589, 
    8.356046, 8.365314, 8.35898, 8.383331, 8.312234, 8.339482, 8.136316, 
    8.1375, 8.143013, 8.118801, 8.117321, 8.095183, 8.114878, 8.123277, 
    8.144627, 8.157278, 8.169319, 8.195845, 8.225554, 8.267238, 8.297288, 
    8.317481, 8.305094, 8.31603, 8.303805, 8.29808, 8.361841, 8.325992, 
    8.379825, 8.376839, 8.352449, 8.377175, 8.13833, 8.131522, 8.107926, 
    8.126388, 8.092775, 8.111578, 8.122406, 8.164289, 8.173512, 8.182076, 
    8.199007, 8.220779, 8.259088, 8.292533, 8.323157, 8.32091, 8.321701, 
    8.328555, 8.311587, 8.331344, 8.334664, 8.325986, 8.376439, 8.362, 
    8.376775, 8.367371, 8.133735, 8.145195, 8.139001, 8.150652, 8.142443, 
    8.178999, 8.189985, 8.241548, 8.220351, 8.254103, 8.223774, 8.229142, 
    8.255211, 8.22541, 8.290689, 8.246391, 8.328822, 8.284428, 8.331611, 
    8.323025, 8.337242, 8.349994, 8.366055, 8.395761, 8.388874, 8.413762, 
    8.162302, 8.177213, 8.175897, 8.19152, 8.203091, 8.228211, 8.268635, 
    8.253415, 8.281372, 8.286994, 8.244526, 8.270582, 8.187201, 8.200629, 
    8.192631, 8.163479, 8.256924, 8.208861, 8.297786, 8.271617, 8.348175, 
    8.310034, 8.385086, 8.41734, 8.447775, 8.483466, 8.185356, 8.175215, 
    8.193378, 8.218568, 8.241988, 8.273211, 8.27641, 8.282272, 8.297471, 
    8.310267, 8.284129, 8.313478, 8.203751, 8.261105, 8.171386, 8.198322, 
    8.21708, 8.208844, 8.251676, 8.261798, 8.303033, 8.281695, 8.409373, 
    8.352693, 8.510712, 8.466318, 8.171675, 8.185321, 8.23296, 8.210265, 
    8.275298, 8.29137, 8.304452, 8.321203, 8.323011, 8.33295, 8.316669, 
    8.332306, 8.273278, 8.299614, 8.227501, 8.245008, 8.236949, 8.228119, 
    8.255396, 8.284541, 8.285161, 8.294525, 8.320965, 8.275562, 8.416718, 
    8.329326, 8.200222, 8.226602, 8.230371, 8.22014, 8.289758, 8.264479, 
    8.332707, 8.314222, 8.344525, 8.329456, 8.327242, 8.307923, 8.295915, 
    8.265637, 8.241067, 8.221623, 8.226141, 8.247511, 8.286325, 8.323176, 
    8.315094, 8.342219, 8.270569, 8.300555, 8.288957, 8.319226, 8.253012, 
    8.309382, 8.238653, 8.244835, 8.263978, 8.302595, 8.311152, 8.320304, 
    8.314654, 8.287312, 8.282838, 8.263511, 8.258183, 8.243488, 8.231339, 
    8.242439, 8.25411, 8.287322, 8.317346, 8.350177, 8.358225, 8.396755, 
    8.365385, 8.417208, 8.373141, 8.449534, 8.312653, 8.37184, 8.264849, 
    8.27632, 8.297109, 8.344934, 8.319083, 8.349321, 8.282662, 8.248251, 
    8.239362, 8.222805, 8.23974, 8.238361, 8.254591, 8.249372, 8.288426, 
    8.26743, 8.327187, 8.349081, 8.411152, 8.449387, 8.488441, 8.505731, 
    8.510998, 8.513201,
  12.66455, 12.72001, 12.70921, 12.75408, 12.72917, 12.75858, 12.67577, 
    12.72222, 12.69255, 12.66953, 12.84158, 12.75608, 12.93093, 12.87599, 
    13.01441, 12.92237, 13.03304, 13.01174, 13.07593, 13.05751, 13.13995, 
    13.08444, 13.18286, 13.12667, 13.13545, 13.08261, 12.77324, 12.83091, 
    12.76983, 12.77804, 12.77436, 12.72969, 12.70724, 12.66032, 12.66882, 
    12.70329, 12.78173, 12.75505, 12.82239, 12.82086, 12.89621, 12.86219, 
    12.98945, 12.95316, 13.05828, 13.03177, 13.05703, 13.04937, 13.05713, 
    13.01827, 13.03491, 13.00076, 12.86856, 12.90728, 12.7921, 12.72332, 
    12.67781, 12.64561, 12.65016, 12.65883, 12.70349, 12.7456, 12.77778, 
    12.79936, 12.82064, 12.88529, 12.91962, 12.9968, 12.98284, 13.0065, 
    13.02913, 13.06723, 13.06095, 13.07776, 13.00587, 13.05361, 12.97489, 
    12.99638, 12.82646, 12.76224, 12.73505, 12.71129, 12.65366, 12.69343, 
    12.67774, 12.7151, 12.73889, 12.72712, 12.79995, 12.77159, 12.92166, 
    12.85682, 13.02649, 12.9857, 13.03629, 13.01045, 13.05475, 13.01487, 
    13.08402, 13.09912, 13.0888, 13.12849, 13.01267, 13.05704, 12.72679, 
    12.72871, 12.73765, 12.69838, 12.69598, 12.66008, 12.69202, 12.70564, 
    12.74027, 12.7608, 12.78035, 12.82342, 12.87168, 12.93945, 12.98834, 
    13.02121, 13.00105, 13.01885, 12.99895, 12.98963, 13.09346, 13.03507, 
    13.12277, 13.1179, 13.07816, 13.11845, 12.73006, 12.71901, 12.68074, 
    12.71068, 12.65618, 12.68666, 12.70423, 12.77218, 12.78716, 12.80106, 
    12.82856, 12.86393, 12.9262, 12.9806, 13.03045, 13.02679, 13.02808, 
    13.03924, 13.01162, 13.04378, 13.04919, 13.03506, 13.11725, 13.09372, 
    13.1178, 13.10247, 12.7226, 12.74119, 12.73114, 12.75005, 12.73673, 
    12.79606, 12.8139, 12.89768, 12.86323, 12.91809, 12.86879, 12.87752, 
    12.91989, 12.87145, 12.9776, 12.90555, 13.03968, 12.96742, 13.04422, 
    13.03024, 13.05339, 13.07416, 13.10033, 13.14875, 13.13752, 13.17811, 
    12.76896, 12.79316, 12.79103, 12.81639, 12.83519, 12.87601, 12.94173, 
    12.91697, 12.96244, 12.97159, 12.90252, 12.94489, 12.80938, 12.83119, 
    12.8182, 12.77087, 12.92268, 12.84456, 12.98915, 12.94658, 13.0712, 
    13.00909, 13.13135, 13.18395, 13.23361, 13.29189, 12.80639, 12.78992, 
    12.81941, 12.86033, 12.8984, 12.94917, 12.95437, 12.96391, 12.98864, 
    13.00947, 12.96693, 13.01469, 12.83626, 12.92948, 12.7837, 12.82744, 
    12.85792, 12.84454, 12.91415, 12.93061, 12.99769, 12.96297, 13.17095, 
    13.07856, 13.33641, 13.26388, 12.78417, 12.80633, 12.88372, 12.84684, 
    12.95256, 12.97871, 13, 13.02727, 13.03021, 13.0464, 13.01989, 13.04535, 
    12.94928, 12.99213, 12.87485, 12.90331, 12.89021, 12.87585, 12.9202, 
    12.9676, 12.96861, 12.98384, 13.02688, 12.95299, 13.18293, 13.0405, 
    12.83053, 12.87339, 12.87951, 12.86289, 12.97609, 12.93497, 13.046, 
    13.0159, 13.06525, 13.04071, 13.0371, 13.00565, 12.98611, 12.93685, 
    12.8969, 12.8653, 12.87264, 12.90738, 12.9705, 13.03048, 13.01732, 
    13.06149, 12.94487, 12.99366, 12.97478, 13.02405, 12.91632, 13.00803, 
    12.89298, 12.90302, 12.93415, 12.99698, 13.01091, 13.02581, 13.01661, 
    12.97211, 12.96483, 12.93339, 12.92473, 12.90084, 12.88109, 12.89913, 
    12.91811, 12.97213, 13.02099, 13.07446, 13.08757, 13.15037, 13.09924, 
    13.18373, 13.11187, 13.23648, 13.01335, 13.10975, 12.93557, 12.95423, 
    12.98805, 13.06592, 13.02382, 13.07306, 12.96454, 12.90858, 12.89413, 
    12.86722, 12.89474, 12.8925, 12.91889, 12.9104, 12.97392, 12.93977, 
    13.03701, 13.07267, 13.17385, 13.23624, 13.30002, 13.32827, 13.33687, 
    13.34047,
  20.59553, 20.69158, 20.67287, 20.75063, 20.70745, 20.75843, 20.61496, 
    20.69541, 20.64401, 20.60415, 20.90251, 20.75411, 21.05789, 20.96232, 
    21.20334, 21.04299, 21.23583, 21.19868, 21.3107, 21.27854, 21.42258, 
    21.32556, 21.49767, 21.39936, 21.41471, 21.32237, 20.78387, 20.88397, 
    20.77796, 20.79219, 20.7858, 20.70834, 20.66944, 20.5882, 20.60292, 
    20.6626, 20.7986, 20.75231, 20.86917, 20.86652, 20.99748, 20.93832, 
    21.15982, 21.09659, 21.27988, 21.23362, 21.27771, 21.26433, 21.27788, 
    21.21008, 21.2391, 21.17954, 20.94938, 21.01673, 20.8166, 20.69731, 
    20.61848, 20.56276, 20.57063, 20.58563, 20.66295, 20.73593, 20.79175, 
    20.82918, 20.86614, 20.97849, 21.0382, 21.17264, 21.14829, 21.18954, 
    21.22902, 21.2955, 21.28454, 21.31389, 21.18845, 21.27173, 21.13445, 
    21.17189, 20.87623, 20.76479, 20.71765, 20.67646, 20.57668, 20.64553, 
    20.61836, 20.68306, 20.7243, 20.70389, 20.83021, 20.781, 21.04175, 
    20.92898, 21.22441, 21.15329, 21.2415, 21.19643, 21.27372, 21.20415, 
    21.32483, 21.35121, 21.33318, 21.40253, 21.2003, 21.27771, 20.70332, 
    20.70665, 20.72216, 20.6541, 20.64994, 20.5878, 20.64308, 20.66668, 
    20.72669, 20.76229, 20.7962, 20.87096, 20.95482, 21.07273, 21.15789, 
    21.2152, 21.18003, 21.21107, 21.17638, 21.16014, 21.34132, 21.23937, 
    21.39254, 21.38403, 21.31459, 21.38499, 20.70899, 20.68985, 20.62356, 
    20.67542, 20.58105, 20.63381, 20.66423, 20.78203, 20.80801, 20.83214, 
    20.87988, 20.94134, 21.04965, 21.1444, 21.23132, 21.22494, 21.22718, 
    21.24665, 21.19847, 21.25458, 21.26401, 21.23936, 21.38289, 21.34177, 
    21.38385, 21.35707, 20.69607, 20.72829, 20.71087, 20.74364, 20.72055, 
    20.82347, 20.85443, 21.00003, 20.94013, 21.03554, 20.9498, 20.96496, 
    21.03868, 20.95442, 21.13917, 21.01373, 21.24741, 21.12143, 21.25533, 
    21.23094, 21.27134, 21.30761, 21.35332, 21.43797, 21.41833, 21.48935, 
    20.77644, 20.81843, 20.81472, 20.85876, 20.8914, 20.96234, 21.07668, 
    21.0336, 21.11276, 21.1287, 21.00845, 21.0822, 20.84659, 20.88446, 
    20.86189, 20.77975, 21.04353, 20.90769, 21.1593, 21.08513, 21.30243, 
    21.19405, 21.40754, 21.49956, 21.58656, 21.68877, 20.84138, 20.81281, 
    20.86401, 20.93509, 21.00128, 21.08964, 21.09871, 21.11532, 21.15841, 
    21.19472, 21.12058, 21.20383, 20.89326, 21.05536, 20.80202, 20.87795, 
    20.93089, 20.90764, 21.02868, 21.05732, 21.17419, 21.11368, 21.47681, 
    21.31528, 21.76694, 21.63964, 20.80283, 20.84128, 20.97575, 20.91165, 
    21.09555, 21.14111, 21.17821, 21.22577, 21.2309, 21.25914, 21.21289, 
    21.25731, 21.08983, 21.16449, 20.96033, 21.00982, 20.98703, 20.96207, 
    21.03921, 21.12175, 21.1235, 21.15005, 21.22509, 21.0963, 21.49779, 
    21.24884, 20.88331, 20.95779, 20.96844, 20.93954, 21.13654, 21.06491, 
    21.25845, 21.20594, 21.29205, 21.24921, 21.24292, 21.18806, 21.15399, 
    21.06819, 20.99867, 20.94372, 20.95648, 21.0169, 21.1268, 21.23137, 
    21.20842, 21.28549, 21.08216, 21.16716, 21.13426, 21.22015, 21.03246, 
    21.1922, 20.99185, 21.00933, 21.0635, 21.17294, 21.19723, 21.22321, 
    21.20717, 21.1296, 21.11692, 21.06217, 21.04709, 21.00552, 20.97117, 
    21.00255, 21.03557, 21.12963, 21.21481, 21.30812, 21.33103, 21.44081, 
    21.35141, 21.49918, 21.3735, 21.59159, 21.20149, 21.36979, 21.06596, 
    21.09845, 21.15738, 21.29321, 21.21975, 21.30569, 21.11642, 21.01899, 
    20.99385, 20.94706, 20.99492, 20.99102, 21.03693, 21.02216, 21.13276, 
    21.07327, 21.24277, 21.30501, 21.48189, 21.59117, 21.70304, 21.75264, 
    21.76776, 21.77409,
  34.63897, 34.81973, 34.78447, 34.93106, 34.84963, 34.94578, 34.6755, 
    34.82694, 34.73015, 34.65517, 35.21813, 34.93762, 35.51293, 35.33146, 
    35.78991, 35.48461, 35.85193, 35.78102, 35.99502, 35.93352, 36.20935, 
    36.02346, 36.35355, 36.16482, 36.19426, 36.01735, 34.99379, 35.18303, 
    34.98262, 35.00951, 34.99744, 34.85131, 34.77802, 34.6252, 34.65287, 
    34.76514, 35.02161, 34.93423, 35.15501, 35.15001, 35.39817, 35.28596, 
    35.70693, 35.58653, 35.93608, 35.8477, 35.93193, 35.90635, 35.93226, 
    35.80277, 35.85817, 35.74452, 35.30694, 35.43473, 35.05561, 34.83052, 
    34.68213, 34.57739, 34.59217, 34.62037, 34.7658, 34.90333, 35.00867, 
    35.0794, 35.14928, 35.36213, 35.47551, 35.73136, 35.68497, 35.7636, 
    35.83892, 35.96595, 35.945, 36.00113, 35.76151, 35.9205, 35.65859, 
    35.72994, 35.16838, 34.95776, 34.86885, 34.79125, 34.60354, 34.73301, 
    34.68189, 34.80368, 34.8814, 34.84293, 35.08133, 34.98837, 35.48225, 
    35.26827, 35.83013, 35.69448, 35.86275, 35.77674, 35.92431, 35.79145, 
    36.02205, 36.07256, 36.03803, 36.17091, 35.78411, 35.93193, 34.84185, 
    34.84812, 34.87735, 34.74914, 34.74132, 34.62444, 34.7284, 34.77282, 
    34.88591, 34.95306, 35.01707, 35.15841, 35.31726, 35.54113, 35.70325, 
    35.81254, 35.74546, 35.80467, 35.73849, 35.70753, 36.05362, 35.85868, 
    36.15175, 36.13544, 36.00246, 36.13728, 34.85253, 34.81646, 34.69168, 
    34.78928, 34.61175, 34.71097, 34.76821, 34.99032, 35.03938, 35.08499, 
    35.17529, 35.29169, 35.49726, 35.67756, 35.84331, 35.83113, 35.83541, 
    35.8726, 35.78061, 35.88773, 35.90576, 35.85865, 36.13326, 36.05449, 
    36.13509, 36.08377, 34.82817, 34.88892, 34.85608, 34.91788, 34.87433, 
    35.0686, 35.12715, 35.40302, 35.2894, 35.47046, 35.30773, 35.33649, 
    35.47642, 35.31649, 35.66759, 35.42902, 35.87404, 35.6338, 35.88918, 
    35.84259, 35.91977, 35.9891, 36.0766, 36.2389, 36.20121, 36.33756, 
    34.97976, 35.05908, 35.05207, 35.13533, 35.1971, 35.3315, 35.54866, 
    35.46676, 35.61731, 35.64765, 35.41901, 35.55915, 35.1123, 35.18395, 
    35.14126, 34.98601, 35.48563, 35.22794, 35.70594, 35.56472, 35.97921, 
    35.7722, 36.1805, 36.3572, 36.52462, 36.72183, 35.10247, 35.04845, 
    35.14525, 35.27985, 35.40538, 35.57331, 35.59055, 35.62217, 35.70424, 
    35.77346, 35.63218, 35.79085, 35.20062, 35.50812, 35.02806, 35.17163, 
    35.27189, 35.22785, 35.45742, 35.51185, 35.73432, 35.61905, 36.31348, 
    36.00379, 36.87302, 36.62696, 35.0296, 35.10228, 35.35695, 35.23544, 
    35.58456, 35.67128, 35.74199, 35.83271, 35.84252, 35.89645, 35.80814, 
    35.89295, 35.57367, 35.71583, 35.32769, 35.42159, 35.37835, 35.33101, 
    35.47742, 35.63441, 35.63775, 35.68832, 35.83142, 35.58598, 36.35378, 
    35.87677, 35.18178, 35.32288, 35.34307, 35.28827, 35.66257, 35.52628, 
    35.89513, 35.79488, 35.95935, 35.87749, 35.86547, 35.76077, 35.69583, 
    35.53252, 35.40044, 35.29621, 35.32041, 35.43504, 35.64404, 35.84341, 
    35.7996, 35.94681, 35.55907, 35.72091, 35.65824, 35.822, 35.4646, 
    35.76867, 35.38749, 35.42067, 35.52358, 35.73195, 35.77826, 35.82784, 
    35.79723, 35.64936, 35.62521, 35.52107, 35.4924, 35.41344, 35.34827, 
    35.40781, 35.4705, 35.64942, 35.8118, 35.99009, 36.03392, 36.24434, 
    36.07294, 36.35647, 36.11525, 36.53432, 35.78638, 36.10815, 35.52827, 
    35.59007, 35.70228, 35.96158, 35.82122, 35.98544, 35.62427, 35.43901, 
    35.39129, 35.30254, 35.39332, 35.38593, 35.47309, 35.44504, 35.65538, 
    35.54217, 35.86517, 35.98413, 36.32324, 36.53351, 36.7494, 36.84533, 
    36.87461, 36.88686,
  60.67812, 61.07083, 60.99409, 61.31372, 61.13599, 61.34588, 60.75732, 
    61.08654, 60.87596, 60.71325, 61.9436, 61.32805, 62.59597, 62.19373, 
    63.21417, 62.53306, 63.35332, 63.19427, 63.67535, 63.53676, 64.1604, 
    63.73951, 64.48857, 64.05934, 64.12612, 63.72573, 61.45091, 61.86631, 
    61.42648, 61.48533, 61.4589, 61.13966, 60.98005, 60.64828, 60.70824, 
    60.95203, 61.51183, 61.32064, 61.80466, 61.79365, 62.34135, 62.09321, 
    63.02843, 62.75974, 63.54253, 63.34382, 63.53318, 63.47563, 63.53393, 
    63.243, 63.36732, 63.11252, 62.13954, 62.42237, 61.58636, 61.09434, 
    60.77169, 60.54478, 60.57676, 60.63782, 60.95346, 61.25314, 61.48349, 
    61.63854, 61.79206, 62.26156, 62.51286, 63.08306, 62.97934, 63.15522, 
    63.32412, 63.60981, 63.5626, 63.68912, 63.15054, 63.50746, 62.92043, 
    63.0799, 61.83408, 61.3721, 61.17791, 61.00883, 60.60137, 60.88219, 
    60.77119, 61.03589, 61.20528, 61.12138, 61.64279, 61.43905, 62.52781, 
    62.05416, 63.30437, 63.0006, 63.37762, 63.18466, 63.51603, 63.21764, 
    63.73632, 63.85044, 63.77242, 64.07315, 63.20118, 63.53319, 61.11904, 
    61.13271, 61.19645, 60.91724, 60.90023, 60.64664, 60.87217, 60.96872, 
    61.21512, 61.36181, 61.5019, 61.81213, 62.16233, 62.65868, 63.0202, 
    63.26491, 63.11462, 63.24727, 63.09903, 63.02978, 63.80764, 63.36849, 
    64.02972, 63.99275, 63.69214, 63.99691, 61.14231, 61.06372, 60.79243, 
    61.00453, 60.61915, 60.8343, 60.95869, 61.44332, 61.55079, 61.65081, 
    61.84927, 62.10587, 62.56117, 62.96279, 63.33397, 63.30662, 63.31624, 
    63.39974, 63.19334, 63.43375, 63.4743, 63.36842, 63.98781, 63.80959, 
    63.99197, 63.8758, 61.08924, 61.22169, 61.15005, 61.28492, 61.18985, 
    61.61485, 61.7434, 62.35209, 62.1008, 62.50164, 62.14127, 62.20483, 
    62.51487, 62.16063, 62.94054, 62.40971, 63.40299, 62.8651, 63.43701, 
    63.33235, 63.50581, 63.66199, 63.85958, 64.22751, 64.14191, 64.4521, 
    61.4202, 61.59397, 61.57861, 61.76139, 61.89728, 62.19381, 62.67543, 
    62.49343, 62.82833, 62.89601, 62.38752, 62.69877, 61.71079, 61.86833, 
    61.77442, 61.43389, 62.53532, 61.96521, 63.02622, 62.71117, 63.63968, 
    63.17449, 64.0949, 64.49689, 64.87986, 65.33361, 61.68919, 61.57065, 
    61.7832, 62.07972, 62.35733, 62.7303, 62.7687, 62.83917, 63.02241, 
    63.17733, 62.86151, 63.21629, 61.90504, 62.58529, 61.52598, 61.84122, 
    62.06215, 61.96502, 62.4727, 62.59358, 63.08968, 62.83222, 64.39722, 
    63.69513, 65.68346, 65.11497, 61.52935, 61.68877, 62.2501, 61.98175, 
    62.75534, 62.94876, 63.10686, 63.31018, 63.33218, 63.45336, 63.25504, 
    63.44549, 62.7311, 63.04832, 62.18539, 62.39325, 62.29744, 62.19271, 
    62.51709, 62.86647, 62.87393, 62.98683, 63.30727, 62.75852, 64.48909, 
    63.40913, 61.86354, 62.17475, 62.2194, 62.09831, 62.92932, 62.62565, 
    63.45039, 63.22533, 63.59494, 63.41073, 63.38372, 63.14891, 63.00361, 
    62.63952, 62.34637, 62.11584, 62.16929, 62.42305, 62.88795, 63.3342, 
    63.23591, 63.56669, 62.6986, 63.0597, 62.91965, 63.28613, 62.48862, 
    63.16659, 62.31769, 62.39119, 62.61966, 63.08437, 63.18806, 63.29924, 
    63.23058, 62.89984, 62.84597, 62.61407, 62.55037, 62.37517, 62.23088, 
    62.3627, 62.50174, 62.89996, 63.26326, 63.66423, 63.76313, 64.23988, 
    63.8513, 64.49522, 63.94703, 64.90211, 63.20626, 63.93095, 62.63008, 
    62.76763, 63.01803, 63.59995, 63.2844, 63.65373, 62.84385, 62.43187, 
    62.3261, 62.12981, 62.3306, 62.31422, 62.50748, 62.44524, 62.91327, 
    62.66099, 63.38305, 63.65079, 64.41946, 64.90024, 65.39728, 65.61927, 
    65.68715, 65.71558,
  116.3177, 117.5456, 117.3041, 118.3151, 117.7513, 118.4176, 116.5637, 
    117.5951, 116.9338, 116.4267, 120.3481, 118.3608, 122.5137, 121.171, 
    124.6257, 122.3021, 125.1096, 124.5568, 126.2417, 125.7524, 127.9808, 
    126.4694, 129.1813, 127.615, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9486, 118.3372, 119.895, 119.8591, 121.6609, 120.8392, 
    123.9848, 123.0673, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7257, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9052, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3957, 122.2342, 124.1727, 123.8163, 124.4217, 
    125.0078, 126.0099, 125.8434, 126.2906, 124.4055, 125.6493, 123.6146, 
    124.1618, 119.9907, 118.5013, 117.8839, 117.3504, 116.08, 116.9533, 
    116.6069, 117.4356, 117.9706, 117.7051, 119.3704, 118.7153, 122.2844, 
    120.7108, 124.939, 123.8892, 125.1944, 124.5235, 125.6795, 124.6378, 
    126.4581, 126.8647, 126.5865, 127.6649, 124.5807, 125.7398, 117.6977, 
    117.7409, 117.9426, 117.063, 117.0098, 116.2201, 116.922, 117.2244, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9565, 
    124.8018, 124.2815, 124.7405, 124.2277, 123.9894, 126.712, 125.1625, 
    127.5082, 127.375, 126.3013, 127.39, 117.7713, 117.5232, 116.6731, 
    117.3369, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.8809, 122.3965, 123.7596, 125.0421, 124.9468, 124.9804, 
    125.2717, 124.5536, 125.3907, 125.5329, 125.1623, 127.3572, 126.7189, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9217, 
    119.2802, 119.696, 121.6967, 120.8642, 122.1966, 120.9977, 121.2077, 
    122.241, 121.0616, 123.6834, 121.8889, 125.2831, 123.4257, 125.4021, 
    125.0365, 125.6435, 126.1945, 126.8974, 128.2247, 127.9137, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1967, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8148, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3096, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4883, 127.7435, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7948, 121.7141, 122.9675, 123.0977, 123.3373, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.0139, 
    120.737, 120.4182, 122.0996, 122.5056, 124.1955, 123.3137, 128.8451, 
    126.3119, 133.7281, 131.5293, 119.0049, 119.519, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2547, 124.9592, 125.0359, 125.4594, 124.7675, 
    125.4319, 122.9702, 124.0532, 121.1434, 121.8339, 121.5149, 121.1676, 
    122.2484, 123.4304, 123.4558, 123.842, 124.9491, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1082, 121.256, 120.856, 123.645, 122.6137, 
    125.4491, 124.6644, 125.9574, 125.3102, 125.2157, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.0429, 
    124.7011, 125.8578, 122.8601, 124.0923, 123.612, 124.8756, 122.153, 
    124.461, 121.5822, 121.8271, 122.5935, 124.1772, 124.5353, 124.9212, 
    124.6826, 123.5443, 123.3605, 122.5746, 122.3602, 121.7736, 121.294, 
    121.7321, 122.1969, 123.5447, 124.7961, 126.2024, 126.5534, 128.2697, 
    126.8678, 129.2058, 127.2107, 130.7228, 124.5983, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9751, 124.8695, 126.1652, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5901, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6128, 133.4764, 
    133.7426, 133.8543,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02010275, -0.01977501, -0.01983828, -0.0195772, -0.01972158, 
    -0.01955128, -0.02003586, -0.0197621, -0.0199364, -0.02007303, 
    -0.01908098, -0.01956564, -0.01859137, -0.01889043, -0.01814891, 
    -0.01863755, -0.01805208, -0.01816285, -0.01783174, -0.01792593, 
    -0.01750948, -0.01778846, -0.0172978, -0.01757569, -0.01753189, 
    -0.01779774, -0.01946709, -0.0191406, -0.01948661, -0.01943964, 
    -0.01946071, -0.01971857, -0.01984988, -0.02012807, -0.02007726, 
    -0.01987311, -0.01941856, -0.01957162, -0.01918842, -0.01919698, 
    -0.01877963, -0.01896658, -0.01827973, -0.01847218, -0.01792199, 
    -0.01805866, -0.01792838, -0.01796778, -0.01792786, -0.01812877, 
    -0.01804239, -0.01822028, -0.01893141, -0.01871934, -0.0193595, 
    -0.01975569, -0.02002376, -0.02021632, -0.02018898, -0.02013695, 
    -0.01987192, -0.01962619, -0.01944111, -0.01931835, -0.01919821, 
    -0.01883935, -0.01865243, -0.01824106, -0.0183146, -0.01819023, 
    -0.01807232, -0.01787616, -0.0179083, -0.01782243, -0.01819353, 
    -0.01794596, -0.01835663, -0.0182433, -0.01916556, -0.01953021, 
    -0.01968734, -0.01982609, -0.02016798, -0.0199312, -0.02002418, 
    -0.01980377, -0.01966506, -0.01973354, -0.019315, -0.01947657, 
    -0.01864142, -0.01899631, -0.01808603, -0.01829949, -0.01803527, 
    -0.01816958, -0.0179401, -0.01814649, -0.0177906, -0.0177141, 
    -0.01776634, -0.01756662, -0.018158, -0.01792836, -0.01973545, 
    -0.01972426, -0.01967225, -0.01990201, -0.01991616, -0.02012946, 
    -0.01993956, -0.01985927, -0.01965706, -0.01953847, -0.01942646, 
    -0.01918261, -0.01891415, -0.01854556, -0.01828557, -0.01811349, 
    -0.0182188, -0.01812579, -0.0182298, -0.01827877, -0.01774271, 
    -0.01804158, -0.0175952, -0.01761959, -0.01782039, -0.01761683, 
    -0.01971641, -0.01978086, -0.02000633, -0.01982964, -0.02015284, 
    -0.01997122, -0.01986758, -0.01947314, -0.01938765, -0.0193087, 
    -0.0191538, -0.01895696, -0.0186169, -0.01832639, -0.01806549, 
    -0.01808447, -0.01807779, -0.01802, -0.01816349, -0.01799656, 
    -0.01796869, -0.01804163, -0.01762285, -0.01774141, -0.0176201, 
    -0.01769719, -0.01975989, -0.01965171, -0.01971008, -0.01960046, 
    -0.01967761, -0.01933701, -0.01923613, -0.01877162, -0.01896081, 
    -0.0186607, -0.0189301, -0.01888205, -0.01865095, -0.01891544, 
    -0.01834226, -0.01872873, -0.01801776, -0.01839625, -0.01799432, 
    -0.01806661, -0.0179471, -0.01784077, -0.017708, -0.01746579, 
    -0.01752156, -0.01732109, -0.01949164, -0.01935348, -0.01936563, 
    -0.0192221, -0.01911669, -0.01889037, -0.01853337, -0.01866676, 
    -0.01842269, -0.0183741, -0.01874523, -0.01851639, -0.01926163, 
    -0.01913904, -0.01921195, -0.01948069, -0.0186359, -0.01906439, 
    -0.0182813, -0.01850738, -0.01785589, -0.01817671, -0.01755234, 
    -0.01729249, -0.01705186, -0.01677512, -0.01927856, -0.01937192, 
    -0.01920512, -0.01897684, -0.01876771, -0.0184935, -0.0184657, 
    -0.01841489, -0.018284, -0.01817472, -0.01839883, -0.01814744, 
    -0.01911068, -0.01859921, -0.01940732, -0.01916004, -0.01899022, 
    -0.01906454, -0.01868208, -0.01859314, -0.01823639, -0.01841989, 
    -0.01735622, -0.01781837, -0.01656775, -0.01690734, -0.01940465, 
    -0.01927889, -0.01884797, -0.0190517, -0.01847536, -0.01833639, 
    -0.01822428, -0.018082, -0.01806672, -0.01798307, -0.01812037, 
    -0.01798848, -0.01849292, -0.01826563, -0.01889673, -0.01874097, 
    -0.01881246, -0.0188912, -0.01864932, -0.01839527, -0.01838993, 
    -0.01830928, -0.01808399, -0.01847307, -0.01729745, -0.0180135, 
    -0.01914275, -0.01890476, -0.01887107, -0.0189627, -0.01835027, 
    -0.01856967, -0.01798511, -0.01814112, -0.01788627, -0.01801242, 
    -0.01803106, -0.01819468, -0.01829735, -0.01855954, -0.01877588, 
    -0.01894939, -0.01890889, -0.01871883, -0.01837987, -0.01806533, 
    -0.01813372, -0.01790551, -0.01851651, -0.01825758, -0.01835718, 
    -0.01809871, -0.01867031, -0.01818224, -0.01879731, -0.0187425, 
    -0.01857406, -0.01824014, -0.0181672, -0.0180896, -0.01813745, 
    -0.01837135, -0.01841, -0.01857814, -0.01862483, -0.01875442, 
    -0.01886243, -0.01876371, -0.01866063, -0.01837127, -0.01811464, 
    -0.01783926, -0.01777258, -0.01745775, -0.01771352, -0.01729354, 
    -0.01764982, -0.01703806, -0.01815444, -0.0176605, -0.01856644, 
    -0.01846648, -0.0182871, -0.01788286, -0.01809992, -0.01784636, 
    -0.01841152, -0.01871229, -0.01879102, -0.01893878, -0.01878766, 
    -0.0187999, -0.0186564, -0.01870239, -0.01836175, -0.01854389, 
    -0.01803152, -0.01784836, -0.01734197, -0.01703923, -0.016737, 
    -0.01660542, -0.0165656, -0.01654898,
  -0.05392943, -0.05288667, -0.05308774, -0.05225881, -0.05271698, 
    -0.05217662, -0.05371634, -0.05284567, -0.05339978, -0.05383474, 
    -0.05068873, -0.05222216, -0.04914657, -0.05008766, -0.04775909, 
    -0.04929172, -0.04745623, -0.04780269, -0.04676819, -0.04706212, 
    -0.04576458, -0.04663319, -0.04510711, -0.0459705, -0.04583425, 
    -0.04666212, -0.05190979, -0.05087699, -0.05197164, -0.05182284, 
    -0.05188958, -0.05270743, -0.05312464, -0.0540101, -0.05384822, 
    -0.05319848, -0.05175608, -0.05224111, -0.05102803, -0.0510551, 
    -0.04973868, -0.05032773, -0.0481687, -0.04877222, -0.04704981, 
    -0.04747681, -0.04706976, -0.04719281, -0.04706816, -0.04769607, 
    -0.04742596, -0.0479825, -0.05021683, -0.04954894, -0.0515691, 
    -0.05282532, -0.05367781, -0.05429145, -0.05420425, -0.05403841, 
    -0.0531947, -0.0524142, -0.05182748, -0.05143887, -0.05105899, 
    -0.04992677, -0.04933851, -0.04804758, -0.04827797, -0.04788843, 
    -0.04751952, -0.04690678, -0.04700707, -0.04673915, -0.04789873, 
    -0.04712469, -0.04840971, -0.04805459, -0.05095584, -0.0521098, 
    -0.05260827, -0.05304901, -0.0541373, -0.05338324, -0.05367916, 
    -0.05297806, -0.05253753, -0.05275494, -0.05142828, -0.05193981, 
    -0.04930387, -0.05042151, -0.04756239, -0.0482306, -0.0474037, 
    -0.04782378, -0.04710637, -0.04775151, -0.04663988, -0.04640144, 
    -0.04656423, -0.04594228, -0.04778754, -0.04706973, -0.05276103, 
    -0.0527255, -0.05256036, -0.05329038, -0.05333541, -0.05401452, 
    -0.05340984, -0.05315448, -0.05251215, -0.052136, -0.05178109, 
    -0.05100969, -0.05016243, -0.04900263, -0.04818698, -0.04764827, 
    -0.04797786, -0.04768675, -0.04801229, -0.04816569, -0.0464906, 
    -0.04742342, -0.04603119, -0.04610709, -0.04673278, -0.04609854, 
    -0.05270058, -0.05290526, -0.05362232, -0.05306029, -0.05408903, 
    -0.05351058, -0.0531809, -0.05192898, -0.0516582, -0.05140833, 
    -0.05091866, -0.05029739, -0.04922679, -0.04831493, -0.04749816, 
    -0.04755751, -0.04753661, -0.04735596, -0.04780472, -0.04728272, 
    -0.04719567, -0.04742358, -0.04611727, -0.04648654, -0.04610871, 
    -0.04634875, -0.05283865, -0.05249519, -0.05268048, -0.05233259, 
    -0.05257739, -0.05149793, -0.05117886, -0.04971346, -0.05030953, 
    -0.0493645, -0.05021269, -0.05006126, -0.04933384, -0.05016649, 
    -0.04836467, -0.04957848, -0.04734895, -0.04853397, -0.04727572, 
    -0.04750166, -0.04712822, -0.04679636, -0.04638244, -0.04562875, 
    -0.04580213, -0.04517936, -0.05198757, -0.05155006, -0.05158849, 
    -0.05113449, -0.05080143, -0.05008747, -0.04896433, -0.04938354, 
    -0.04861689, -0.04846449, -0.04963041, -0.04891101, -0.05125948, 
    -0.05087205, -0.05110241, -0.05195287, -0.04928651, -0.05063631, 
    -0.04817361, -0.04888273, -0.04684352, -0.04784608, -0.04589786, 
    -0.04509065, -0.04434501, -0.04348984, -0.051313, -0.05160841, 
    -0.0510808, -0.05036008, -0.04970117, -0.04883914, -0.04875188, 
    -0.04859244, -0.04818207, -0.04783985, -0.04854207, -0.04775448, 
    -0.0507825, -0.04917118, -0.05172049, -0.05093837, -0.0504023, 
    -0.05063679, -0.04943172, -0.04915211, -0.04803294, -0.04860812, 
    -0.04528841, -0.04672649, -0.04285068, -0.04389814, -0.05171202, 
    -0.05131405, -0.0499539, -0.05059626, -0.0487822, -0.04834628, -0.047995, 
    -0.04754978, -0.04750203, -0.04724059, -0.04766979, -0.04725749, 
    -0.04883733, -0.04812454, -0.05010751, -0.049617, -0.04984204, 
    -0.05009008, -0.04932872, -0.04853091, -0.04851413, -0.04826128, 
    -0.04755606, -0.04877499, -0.04510605, -0.0473357, -0.05088376, 
    -0.05013283, -0.05002668, -0.0503155, -0.04838979, -0.04907837, 
    -0.04724696, -0.0477347, -0.04693833, -0.04733228, -0.04739052, 
    -0.04790233, -0.04822389, -0.04904655, -0.04972688, -0.05027351, 
    -0.05014585, -0.04954734, -0.04848258, -0.04749765, -0.04771156, 
    -0.04699836, -0.04891139, -0.04809931, -0.04841144, -0.04760206, 
    -0.04939471, -0.04786341, -0.04979433, -0.04962181, -0.04909214, 
    -0.04804467, -0.04781631, -0.04757355, -0.04772322, -0.04845589, 
    -0.04857711, -0.04910497, -0.04925172, -0.04965933, -0.04999943, 
    -0.04968857, -0.04936428, -0.04845563, -0.04765186, -0.04679164, 
    -0.04658368, -0.04560377, -0.04639963, -0.04509393, -0.04620127, 
    -0.04430235, -0.0477764, -0.04623449, -0.04906822, -0.04875431, 
    -0.0481918, -0.04692768, -0.04760583, -0.0468138, -0.04858187, 
    -0.04952677, -0.04977454, -0.05024008, -0.04976394, -0.0498025, 
    -0.04935098, -0.04949561, -0.04842576, -0.04899736, -0.04739196, 
    -0.04682003, -0.04524416, -0.04430595, -0.04337225, -0.04296667, 
    -0.04284403, -0.04279287,
  -0.07870924, -0.07705818, -0.07737636, -0.07606516, -0.07678971, 
    -0.07593523, -0.07837165, -0.07699331, -0.07787032, -0.07855922, 
    -0.07358571, -0.07600722, -0.0711557, -0.07263794, -0.06897408, 
    -0.07138418, -0.06849848, -0.06904257, -0.06741881, -0.0678799, 
    -0.06584604, -0.06720711, -0.06481704, -0.06616854, -0.06595513, 
    -0.06725248, -0.07551352, -0.07388272, -0.07561126, -0.07537615, 
    -0.07548159, -0.0767746, -0.07743477, -0.07883705, -0.07858057, 
    -0.07755164, -0.07527067, -0.07603717, -0.07412106, -0.07416377, 
    -0.07208805, -0.07301638, -0.06961767, -0.07056662, -0.0678606, 
    -0.06853079, -0.0678919, -0.06808499, -0.06788938, -0.0688751, 
    -0.06845095, -0.06932504, -0.07284154, -0.0717892, -0.07497531, 
    -0.07696112, -0.07831063, -0.07928298, -0.07914475, -0.07888192, 
    -0.07754566, -0.07631084, -0.07538347, -0.07476964, -0.07416992, 
    -0.07238439, -0.07145784, -0.06942732, -0.06978942, -0.06917726, 
    -0.06859785, -0.0676362, -0.06779353, -0.06737328, -0.06919344, 
    -0.06797808, -0.06999652, -0.06943832, -0.07400715, -0.07582962, 
    -0.07661777, -0.07731507, -0.07903864, -0.07784414, -0.07831276, 
    -0.07720278, -0.07650588, -0.07684977, -0.07475293, -0.07556096, 
    -0.07140331, -0.07316426, -0.06866516, -0.06971495, -0.06841601, 
    -0.06907568, -0.06794934, -0.06896217, -0.0672176, -0.06684379, 
    -0.06709899, -0.06612432, -0.06901876, -0.06789184, -0.07685939, 
    -0.07680319, -0.07654198, -0.07769712, -0.07776841, -0.07884407, 
    -0.07788625, -0.07748199, -0.07646573, -0.07587102, -0.07531017, 
    -0.07409212, -0.07275581, -0.07092916, -0.06964639, -0.06880002, 
    -0.06931777, -0.06886046, -0.06937186, -0.06961294, -0.06698356, 
    -0.06844697, -0.0662636, -0.06638252, -0.06736329, -0.06636911, 
    -0.07676376, -0.07708759, -0.07822274, -0.07733292, -0.07896215, 
    -0.07804577, -0.07752381, -0.07554385, -0.07511605, -0.07472142, 
    -0.07394847, -0.07296856, -0.07128196, -0.06984752, -0.06856431, 
    -0.06865751, -0.06862468, -0.06834107, -0.06904575, -0.0682261, 
    -0.06808948, -0.06844721, -0.06639846, -0.06697719, -0.06638505, 
    -0.0667612, -0.07698219, -0.07643891, -0.07673196, -0.07618181, 
    -0.07656892, -0.07486291, -0.07435914, -0.07204833, -0.07298768, 
    -0.07149876, -0.07283503, -0.07259634, -0.07145049, -0.07276219, 
    -0.06992572, -0.07183573, -0.06833007, -0.07019191, -0.06821511, 
    -0.06856981, -0.06798363, -0.067463, -0.06681401, -0.06563336, 
    -0.06590483, -0.06493006, -0.07563642, -0.07494523, -0.07500593, 
    -0.0742891, -0.0737635, -0.07263763, -0.07086889, -0.07152874, 
    -0.07032232, -0.07008265, -0.0719175, -0.07078499, -0.0744864, 
    -0.07387493, -0.07423845, -0.0755816, -0.07137597, -0.07350302, 
    -0.06962537, -0.07074048, -0.06753697, -0.06911073, -0.06605475, 
    -0.06479131, -0.06362566, -0.06229055, -0.0745709, -0.07503739, 
    -0.07420436, -0.0730674, -0.07202896, -0.07067192, -0.07053464, 
    -0.07028385, -0.06963868, -0.06910094, -0.07020465, -0.06896683, 
    -0.07373364, -0.07119443, -0.07521444, -0.07397957, -0.07313397, 
    -0.07350378, -0.07160459, -0.0711644, -0.06940432, -0.07030851, 
    -0.06510069, -0.06735342, -0.06129391, -0.06292776, -0.07520106, 
    -0.07457256, -0.07242714, -0.07343984, -0.07058234, -0.06989679, 
    -0.06934469, -0.06864536, -0.06857038, -0.06815997, -0.06883382, 
    -0.06818649, -0.07066905, -0.06954825, -0.07266922, -0.07189638, 
    -0.07225089, -0.07264175, -0.07144242, -0.07018711, -0.0701607, 
    -0.06976318, -0.06865524, -0.070571, -0.06481541, -0.06830927, 
    -0.0738934, -0.07270915, -0.07254183, -0.07299709, -0.06996521, 
    -0.07104834, -0.06816997, -0.06893576, -0.06768569, -0.06830388, 
    -0.06839532, -0.06919909, -0.06970441, -0.07099827, -0.07206946, 
    -0.0729309, -0.07272966, -0.07178667, -0.0701111, -0.06856351, 
    -0.06889943, -0.06777987, -0.07078558, -0.06950861, -0.06999925, 
    -0.06872745, -0.07154632, -0.06913798, -0.07217573, -0.07190396, 
    -0.07107002, -0.06942276, -0.06906396, -0.06868269, -0.06891773, 
    -0.07006913, -0.07025974, -0.07109021, -0.07132121, -0.07196305, 
    -0.0724989, -0.07200911, -0.07149841, -0.07006872, -0.06880566, 
    -0.0674556, -0.06712949, -0.06559426, -0.06684097, -0.06479645, 
    -0.06653011, -0.06355903, -0.06900127, -0.06658214, -0.07103237, 
    -0.07053846, -0.06965398, -0.06766899, -0.06873337, -0.06749036, 
    -0.07026724, -0.07175428, -0.07214453, -0.07287819, -0.07212785, 
    -0.07218859, -0.07147747, -0.07170519, -0.07002176, -0.07092087, 
    -0.06839757, -0.06750013, -0.06503145, -0.06356463, -0.06210711, 
    -0.06147469, -0.06128355, -0.06120382,
  -0.08618427, -0.08427422, -0.08464219, -0.08312611, -0.08396376, 
    -0.08297592, -0.0857936, -0.0841992, -0.08521358, -0.08601065, 
    -0.08026168, -0.08305913, -0.07745761, -0.07916761, -0.07494303, 
    -0.07772112, -0.07439522, -0.07502193, -0.07315211, -0.0736829, 
    -0.07134254, -0.07290844, -0.07015945, -0.07171346, -0.07146801, 
    -0.07296066, -0.08248852, -0.08060464, -0.08260148, -0.08232977, 
    -0.08245162, -0.0839463, -0.08470976, -0.08633218, -0.08603535, 
    -0.08484493, -0.0822079, -0.08309374, -0.08087985, -0.08092919, 
    -0.07853308, -0.07960439, -0.07568455, -0.07677835, -0.07366068, 
    -0.07443242, -0.07369672, -0.07391904, -0.07369382, -0.074829, 
    -0.07434046, -0.07534736, -0.0794026, -0.07818829, -0.08186662, 
    -0.08416198, -0.085723, -0.08684832, -0.08668832, -0.08638411, 
    -0.08483801, -0.0834101, -0.08233823, -0.08162901, -0.08093628, 
    -0.07887504, -0.07780607, -0.07546521, -0.07588247, -0.07517709, 
    -0.07450965, -0.07340235, -0.07358347, -0.07309969, -0.07519573, 
    -0.07379595, -0.07612116, -0.07547789, -0.08074833, -0.08285384, 
    -0.08376496, -0.08457131, -0.0865655, -0.08518329, -0.08572546, 
    -0.08444144, -0.08363559, -0.0840332, -0.0816097, -0.08254334, 
    -0.07774318, -0.07977511, -0.07458719, -0.07579666, -0.07430023, 
    -0.07506007, -0.07376286, -0.0749293, -0.07292051, -0.07249032, 
    -0.07278401, -0.0716626, -0.0749945, -0.07369666, -0.08404434, 
    -0.08397935, -0.08367731, -0.08501322, -0.08509567, -0.0863403, 
    -0.085232, -0.08476437, -0.08358917, -0.0829017, -0.08225354, 
    -0.08084644, -0.07930364, -0.07719637, -0.07571765, -0.07474252, 
    -0.07533897, -0.07481213, -0.07540131, -0.07567909, -0.07265117, 
    -0.07433589, -0.07182281, -0.07195961, -0.0730882, -0.07194418, 
    -0.08393376, -0.08430821, -0.0856213, -0.08459195, -0.08647696, 
    -0.08541656, -0.08481275, -0.08252358, -0.08202922, -0.08157331, 
    -0.08068054, -0.0795492, -0.07760322, -0.07594944, -0.07447103, 
    -0.07457837, -0.07454056, -0.07421392, -0.07502559, -0.07408153, 
    -0.07392421, -0.07433616, -0.07197795, -0.07264383, -0.07196252, 
    -0.07239529, -0.08418632, -0.08355816, -0.08389699, -0.08326095, 
    -0.08370848, -0.08173677, -0.08115483, -0.07848725, -0.07957128, 
    -0.07785328, -0.07939508, -0.07911961, -0.0777976, -0.07931101, 
    -0.07603956, -0.07824198, -0.07420126, -0.07634639, -0.07406887, 
    -0.07447736, -0.07380233, -0.07320297, -0.07245606, -0.07109796, 
    -0.07141015, -0.07028935, -0.08263056, -0.08183188, -0.081902, 
    -0.08107393, -0.08046695, -0.07916726, -0.07712685, -0.07788785, 
    -0.07649671, -0.07622044, -0.07833631, -0.07703013, -0.08130183, 
    -0.08059563, -0.08101544, -0.08256719, -0.07771165, -0.08016621, 
    -0.07569343, -0.0769788, -0.07328811, -0.07510045, -0.07158258, 
    -0.07012987, -0.0687905, -0.06725754, -0.08139943, -0.08193834, 
    -0.08097605, -0.0796633, -0.0784649, -0.07689974, -0.07674147, 
    -0.07645236, -0.07570876, -0.07508917, -0.07636107, -0.07493467, 
    -0.08043249, -0.07750227, -0.08214291, -0.08071647, -0.07974014, 
    -0.08016707, -0.07797533, -0.07746763, -0.07543871, -0.07648079, 
    -0.07048551, -0.07307684, -0.06611397, -0.06798903, -0.08212746, 
    -0.08140134, -0.07892435, -0.08009325, -0.07679646, -0.07600623, 
    -0.07537, -0.07456437, -0.07447801, -0.07400538, -0.07478146, 
    -0.07403592, -0.07689645, -0.07560456, -0.07920371, -0.07831194, 
    -0.07872096, -0.07917201, -0.07778828, -0.07634084, -0.07631041, 
    -0.07585224, -0.07457577, -0.0767834, -0.07015759, -0.07417732, 
    -0.08061695, -0.07924981, -0.0790567, -0.07958214, -0.07608507, 
    -0.07733379, -0.07401689, -0.07489888, -0.07345932, -0.0741711, 
    -0.0742764, -0.07520224, -0.0757845, -0.07727605, -0.07851163, 
    -0.07950573, -0.07927346, -0.07818538, -0.07625324, -0.07447011, 
    -0.07485703, -0.07356773, -0.07703081, -0.07555888, -0.07612431, 
    -0.07465893, -0.07790813, -0.07513185, -0.07863424, -0.07832069, 
    -0.0773588, -0.07545996, -0.07504657, -0.07460736, -0.0748781, 
    -0.07620486, -0.07642458, -0.07738208, -0.07764848, -0.07838886, 
    -0.07900714, -0.078442, -0.07785287, -0.07620437, -0.07474902, 
    -0.07319444, -0.0728191, -0.071053, -0.07248709, -0.07013579, 
    -0.07212943, -0.06871399, -0.07497436, -0.07218929, -0.07731538, 
    -0.07674588, -0.0757264, -0.0734401, -0.07466576, -0.07323447, 
    -0.07643321, -0.07814801, -0.07859825, -0.0794449, -0.078579, 
    -0.07864907, -0.07782871, -0.07809139, -0.07615025, -0.07718679, 
    -0.074279, -0.07324571, -0.07040591, -0.06872041, -0.067047, -0.06632135, 
    -0.06610209, -0.06601063,
  -0.06732004, -0.06577259, -0.06607071, -0.0648424, -0.06552105, 
    -0.06472071, -0.06700354, -0.06571181, -0.06653363, -0.06717939, 
    -0.06252158, -0.06478814, -0.06024957, -0.06163511, -0.05821211, 
    -0.06046309, -0.05776823, -0.05827603, -0.05676099, -0.05719108, 
    -0.0552948, -0.05656356, -0.05433623, -0.05559534, -0.05539646, 
    -0.05660587, -0.06432582, -0.06279946, -0.06441734, -0.06419721, 
    -0.06429593, -0.06550691, -0.06612546, -0.06743987, -0.06719939, 
    -0.06623497, -0.06409846, -0.06481618, -0.06302244, -0.06306241, 
    -0.06112098, -0.06198902, -0.05881293, -0.0596992, -0.05717307, 
    -0.05779837, -0.05720226, -0.0573824, -0.05719992, -0.05811971, 
    -0.05772387, -0.05853972, -0.06182551, -0.06084162, -0.06382195, 
    -0.06568167, -0.06694634, -0.06785801, -0.06772839, -0.06748194, 
    -0.06622937, -0.06507248, -0.06420405, -0.06362943, -0.06306816, 
    -0.06139806, -0.06053192, -0.05863521, -0.0589733, -0.05840176, 
    -0.05786095, -0.05696375, -0.05711051, -0.05671852, -0.05841686, 
    -0.05728268, -0.0591667, -0.05864548, -0.06291588, -0.06462181, 
    -0.06535999, -0.06601328, -0.06762889, -0.0665091, -0.06694835, 
    -0.06590807, -0.06525518, -0.06557732, -0.06361379, -0.06437024, 
    -0.06048096, -0.06212734, -0.05792378, -0.05890376, -0.05769127, 
    -0.05830694, -0.05725586, -0.05820099, -0.05657335, -0.05622479, 
    -0.05646274, -0.05555413, -0.05825381, -0.05720222, -0.06558634, 
    -0.06553368, -0.06528898, -0.06637131, -0.06643812, -0.06744645, 
    -0.06654856, -0.0661697, -0.06521757, -0.06466058, -0.06413543, 
    -0.06299536, -0.06174533, -0.0600379, -0.05883975, -0.05804964, 
    -0.05853292, -0.05810604, -0.05858343, -0.05880851, -0.05635511, 
    -0.05772016, -0.05568394, -0.05579478, -0.05670922, -0.05578228, 
    -0.06549675, -0.06580013, -0.06686395, -0.06603, -0.06755716, 
    -0.06669807, -0.0662089, -0.06435422, -0.06395369, -0.0635843, 
    -0.06286095, -0.06194429, -0.06036755, -0.05902756, -0.05782966, 
    -0.05791663, -0.05788599, -0.05762134, -0.058279, -0.05751406, 
    -0.0573866, -0.05772039, -0.05580964, -0.05634916, -0.05579714, 
    -0.05614779, -0.06570138, -0.06519245, -0.06546696, -0.06495164, 
    -0.06531423, -0.06371674, -0.06324524, -0.06108385, -0.06196218, 
    -0.06057017, -0.06181942, -0.06159621, -0.06052506, -0.0617513, 
    -0.05910059, -0.06088512, -0.05761107, -0.0593492, -0.05750381, 
    -0.05783479, -0.05728784, -0.05680221, -0.05619702, -0.05509663, 
    -0.05534958, -0.05444149, -0.0644409, -0.0637938, -0.06385062, 
    -0.06317969, -0.06268789, -0.06163483, -0.05998158, -0.06059818, 
    -0.05947099, -0.05924714, -0.06096154, -0.0599032, -0.06336434, 
    -0.06279215, -0.06313229, -0.06438956, -0.06045541, -0.06244422, 
    -0.05882012, -0.05986162, -0.05687119, -0.05833966, -0.05548929, 
    -0.05431227, -0.0532271, -0.05198515, -0.06344341, -0.06388006, 
    -0.06310038, -0.06203675, -0.06106574, -0.05979756, -0.05966932, 
    -0.05943506, -0.05883255, -0.05833052, -0.05936109, -0.05820533, 
    -0.06265997, -0.06028576, -0.0640458, -0.06289006, -0.062099, 
    -0.06244491, -0.06066906, -0.06025769, -0.05861374, -0.0594581, 
    -0.05460042, -0.05670001, -0.05105871, -0.05257777, -0.06403328, 
    -0.06344496, -0.06143801, -0.0623851, -0.05971387, -0.05907357, 
    -0.05855806, -0.0579053, -0.05783532, -0.05745236, -0.05808119, 
    -0.05747711, -0.05979489, -0.05874811, -0.06166436, -0.0609418, 
    -0.06127321, -0.06163868, -0.0605175, -0.0593447, -0.05932004, 
    -0.0589488, -0.05791454, -0.05970328, -0.05433473, -0.05759169, 
    -0.06280942, -0.06170171, -0.06154524, -0.06197098, -0.05913746, 
    -0.06014925, -0.05746169, -0.05817633, -0.05700991, -0.05758664, 
    -0.05767196, -0.05842213, -0.05889392, -0.06010246, -0.0611036, 
    -0.06190907, -0.06172088, -0.06083925, -0.05927372, -0.05782891, 
    -0.05814242, -0.05709776, -0.05990375, -0.0587111, -0.05916925, 
    -0.05798191, -0.06061461, -0.05836511, -0.06120294, -0.06094889, 
    -0.06016951, -0.05863095, -0.05829599, -0.05794013, -0.0581595, 
    -0.05923452, -0.05941254, -0.06018837, -0.06040423, -0.06100413, 
    -0.06150509, -0.06104718, -0.06056983, -0.05923413, -0.0580549, 
    -0.0567953, -0.05649117, -0.05506022, -0.05622217, -0.05431708, 
    -0.05593238, -0.05316512, -0.05823749, -0.05598088, -0.06013433, 
    -0.05967289, -0.05884684, -0.05699434, -0.05798744, -0.05682773, 
    -0.05941954, -0.06080898, -0.06117378, -0.06185978, -0.06115818, 
    -0.06121496, -0.06055025, -0.0607631, -0.05919028, -0.06003014, 
    -0.05767407, -0.05683684, -0.05453592, -0.05317032, -0.05181458, 
    -0.05122671, -0.05104908, -0.05097499,
  -0.06391456, -0.06222175, -0.06254764, -0.06120573, -0.0619469, -0.0610729, 
    -0.06356808, -0.06215534, -0.06305389, -0.06376056, -0.05867596, 
    -0.0611465, -0.05620686, -0.05771168, -0.05399928, -0.05643857, 
    -0.05351921, -0.05406844, -0.05243101, -0.05289546, -0.05084996, 
    -0.05221789, -0.04981826, -0.05117374, -0.05095946, -0.05226356, 
    -0.06064199, -0.05897845, -0.06074184, -0.06050169, -0.06060938, 
    -0.06193145, -0.0626075, -0.06404577, -0.06378247, -0.06272724, 
    -0.06039399, -0.0611771, -0.05922126, -0.0592648, -0.05715295, 
    -0.05809651, -0.0546496, -0.0556099, -0.052876, -0.0535518, -0.05290755, 
    -0.05310217, -0.05290501, -0.05389932, -0.05347124, -0.05435381, 
    -0.05791869, -0.05684952, -0.06009248, -0.06212239, -0.06350547, 
    -0.06450379, -0.06436179, -0.06409185, -0.0627211, -0.06145694, 
    -0.06050916, -0.0598826, -0.05927106, -0.05745401, -0.05651328, 
    -0.05445718, -0.05482327, -0.05420449, -0.05361946, -0.05264993, 
    -0.05280843, -0.05238516, -0.05422083, -0.05299442, -0.05503277, 
    -0.05446829, -0.05910522, -0.06096495, -0.06177095, -0.06248485, 
    -0.06425279, -0.06302705, -0.06350766, -0.06236983, -0.06165646, 
    -0.06200837, -0.05986555, -0.06069045, -0.05645797, -0.05824696, 
    -0.0536874, -0.05474796, -0.053436, -0.05410188, -0.05296544, 
    -0.05398725, -0.05222845, -0.05185237, -0.0521091, -0.05112933, 
    -0.0540444, -0.0529075, -0.06201823, -0.0619607, -0.06169338, 
    -0.06287634, -0.0629494, -0.06405298, -0.06307022, -0.06265587, 
    -0.06161538, -0.06100727, -0.06043431, -0.05919177, -0.05783151, 
    -0.05597721, -0.05467863, -0.05382352, -0.05434645, -0.05388454, 
    -0.05440112, -0.05464481, -0.05199296, -0.05346724, -0.05126922, 
    -0.05138869, -0.05237511, -0.05137521, -0.06192034, -0.06225186, 
    -0.0634153, -0.06250314, -0.06417423, -0.06323379, -0.06269873, 
    -0.06067298, -0.06023612, -0.05983341, -0.0590454, -0.05804787, 
    -0.05633489, -0.05488204, -0.05358562, -0.05367967, -0.05364654, 
    -0.0533604, -0.05407165, -0.05324445, -0.0531067, -0.05346747, 
    -0.05140471, -0.05198655, -0.05139123, -0.05176932, -0.06214393, 
    -0.06158794, -0.0618878, -0.06132499, -0.06172096, -0.05997778, 
    -0.05946396, -0.05711262, -0.05806733, -0.0565548, -0.05791207, 
    -0.0576694, -0.05650584, -0.057838, -0.05496115, -0.05689676, 
    -0.05334931, -0.05523052, -0.05323337, -0.05359117, -0.053, -0.0524755, 
    -0.05182242, -0.05063653, -0.05090896, -0.04993146, -0.06076755, 
    -0.06006179, -0.06012373, -0.05939254, -0.05885698, -0.05771137, 
    -0.05591612, -0.0565852, -0.05536251, -0.05511992, -0.05697977, 
    -0.05583112, -0.05959371, -0.05897049, -0.05934092, -0.06071153, 
    -0.05643024, -0.05859175, -0.05465738, -0.05578601, -0.05254998, 
    -0.05413729, -0.05105947, -0.04979249, -0.04862653, -0.04729471, 
    -0.05967988, -0.06015583, -0.05930616, -0.05814842, -0.05709295, 
    -0.05571655, -0.0555775, -0.05532357, -0.05467084, -0.0541274, 
    -0.0552434, -0.05399195, -0.05882659, -0.05624613, -0.06033656, 
    -0.0590771, -0.05821614, -0.05859251, -0.05666216, -0.05621567, 
    -0.05443393, -0.05534853, -0.05010244, -0.05236518, -0.04630309, 
    -0.04792986, -0.06032291, -0.05968157, -0.05749743, -0.05852742, 
    -0.05562581, -0.05493188, -0.05437366, -0.05366741, -0.05359174, 
    -0.05317777, -0.05385765, -0.05320451, -0.05571366, -0.05457941, 
    -0.05774348, -0.05695833, -0.05731835, -0.05771555, -0.05649763, 
    -0.05522564, -0.05519892, -0.05479674, -0.05367741, -0.05561433, 
    -0.04981665, -0.05332836, -0.0589893, -0.05778408, -0.05761399, 
    -0.05807689, -0.05500109, -0.05609801, -0.05318785, -0.05396057, 
    -0.05269978, -0.0533229, -0.05341513, -0.05422654, -0.0547373, 
    -0.05604725, -0.05713407, -0.05800956, -0.05780492, -0.05684696, 
    -0.05514873, -0.05358482, -0.05392389, -0.05279465, -0.05583171, 
    -0.05453934, -0.05503554, -0.05375027, -0.05660304, -0.05416483, 
    -0.057242, -0.05696603, -0.05611999, -0.05445257, -0.05409004, 
    -0.05370509, -0.05394236, -0.05510625, -0.05529917, -0.05614045, 
    -0.05637469, -0.05702602, -0.05757035, -0.05707279, -0.05655444, 
    -0.05510582, -0.05382922, -0.05246804, -0.05213978, -0.05059732, 
    -0.05184955, -0.04979766, -0.05153703, -0.04855999, -0.05402675, 
    -0.05158933, -0.05608182, -0.05558137, -0.05468631, -0.05268296, 
    -0.05375625, -0.05250306, -0.05530675, -0.05681408, -0.05721032, 
    -0.05795596, -0.05719337, -0.05725506, -0.05653318, -0.05676426, 
    -0.05505832, -0.0559688, -0.05341741, -0.05251289, -0.05003305, 
    -0.04856558, -0.04711202, -0.04648279, -0.0462928, -0.04621357,
  -0.04035198, -0.0390736, -0.03931955, -0.03830725, -0.03886621, 
    -0.03820712, -0.04009017, -0.03902348, -0.03970178, -0.04023561, 
    -0.03640242, -0.0382626, -0.03454812, -0.03567765, -0.03289467, 
    -0.03472192, -0.03253571, -0.03294641, -0.03172284, -0.03206963, 
    -0.03054396, -0.03156378, -0.02977613, -0.03078517, -0.03062552, 
    -0.03159786, -0.03788237, -0.03662993, -0.0379576, -0.03777666, 
    -0.03785779, -0.03885456, -0.03936474, -0.04045115, -0.04025216, 
    -0.03945513, -0.03769552, -0.03828567, -0.03681261, -0.03684536, 
    -0.03525804, -0.03596681, -0.03338129, -0.03410058, -0.0320551, 
    -0.03256007, -0.03207866, -0.03222405, -0.03207677, -0.03281992, 
    -0.03249985, -0.03315992, -0.03583318, -0.03503028, -0.03746842, 
    -0.03899862, -0.04004287, -0.0407974, -0.04069004, -0.04048597, 
    -0.0394505, -0.03849667, -0.03778229, -0.03731038, -0.03685008, 
    -0.03548411, -0.03477797, -0.03323727, -0.03351132, -0.03304819, 
    -0.03261065, -0.03188627, -0.03200463, -0.03168861, -0.03306042, 
    -0.03214355, -0.0336682, -0.03324559, -0.0367253, -0.03812575, 
    -0.03873349, -0.03927216, -0.04060763, -0.03968151, -0.04004452, 
    -0.03918535, -0.03864713, -0.03891259, -0.03729755, -0.03791888, 
    -0.03473647, -0.03607989, -0.03266145, -0.03345493, -0.03247351, 
    -0.03297143, -0.0321219, -0.03288567, -0.03157166, -0.03129109, 
    -0.0314826, -0.03075208, -0.03292842, -0.03207862, -0.03892003, 
    -0.03887663, -0.03867498, -0.03956771, -0.03962288, -0.0404566, 
    -0.03971411, -0.03940125, -0.03861615, -0.03815765, -0.0377259, 
    -0.03679042, -0.03576768, -0.03437592, -0.03340304, -0.03276323, 
    -0.03315441, -0.03280886, -0.03319532, -0.03337771, -0.03139596, 
    -0.03249686, -0.03085632, -0.03094536, -0.03168111, -0.03093532, 
    -0.03884618, -0.03909632, -0.03997475, -0.03928596, -0.04054825, 
    -0.03983765, -0.03943361, -0.03790571, -0.0375766, -0.03727335, 
    -0.0366803, -0.03593025, -0.03464415, -0.03355532, -0.03258536, 
    -0.03265567, -0.0326309, -0.03241701, -0.03294881, -0.03233036, 
    -0.03222743, -0.03249704, -0.0309573, -0.03139117, -0.03094725, 
    -0.03122915, -0.03901488, -0.03859545, -0.03882163, -0.03839717, 
    -0.03869578, -0.03738205, -0.03699524, -0.03522776, -0.03594487, 
    -0.03480912, -0.0358282, -0.03564588, -0.03477238, -0.03577255, 
    -0.03361456, -0.03506573, -0.03240872, -0.03381632, -0.03232208, 
    -0.0325895, -0.03214772, -0.03175605, -0.03126875, -0.03038502, 
    -0.0305879, -0.02986032, -0.03797698, -0.03744531, -0.03749195, 
    -0.03694149, -0.03653856, -0.03567742, -0.03433011, -0.03483193, 
    -0.0339152, -0.03373348, -0.03512803, -0.03426639, -0.03709291, 
    -0.03662394, -0.03690264, -0.03793477, -0.03471567, -0.0363391, 
    -0.03338712, -0.03423258, -0.03181165, -0.03299792, -0.03070002, 
    -0.02975697, -0.0288907, -0.02790317, -0.03715777, -0.03751613, 
    -0.03687649, -0.03600582, -0.035213, -0.03418051, -0.0340763, 
    -0.03388602, -0.0333972, -0.03299051, -0.03382597, -0.03288919, 
    -0.03651571, -0.03457757, -0.03765227, -0.03670414, -0.03605672, 
    -0.03633967, -0.03488967, -0.03455473, -0.03321987, -0.03390473, 
    -0.02998751, -0.0316737, -0.02716935, -0.02837386, -0.03764197, 
    -0.03715903, -0.03551672, -0.03629073, -0.0341125, -0.03359265, 
    -0.03317477, -0.0326465, -0.03258993, -0.03228053, -0.03278875, 
    -0.03230052, -0.03417834, -0.03332876, -0.03570154, -0.03511194, 
    -0.03538223, -0.03568056, -0.03476623, -0.03381266, -0.03379264, 
    -0.03349146, -0.03265398, -0.0341039, -0.02977493, -0.03239306, 
    -0.03663809, -0.03573205, -0.03560426, -0.03595206, -0.03364448, 
    -0.03446649, -0.03228806, -0.03286573, -0.0319235, -0.03238898, 
    -0.03245791, -0.03306469, -0.03344695, -0.03442843, -0.03524387, 
    -0.03590146, -0.0357477, -0.03502835, -0.03375505, -0.03258475, 
    -0.03283829, -0.03199435, -0.03426683, -0.03329877, -0.03367027, 
    -0.03270845, -0.03484531, -0.03301852, -0.0353249, -0.03511772, 
    -0.03448297, -0.03323382, -0.03296257, -0.03267467, -0.03285211, 
    -0.03372324, -0.03386774, -0.03449832, -0.034674, -0.03516275, 
    -0.03557148, -0.03519786, -0.03480885, -0.03372291, -0.03276749, 
    -0.03175048, -0.0315055, -0.03035583, -0.03128899, -0.02976081, 
    -0.03105594, -0.02884131, -0.03291522, -0.03109493, -0.03445435, 
    -0.0340792, -0.03340878, -0.03191094, -0.03271293, -0.03177662, 
    -0.03387342, -0.03500368, -0.03530111, -0.03586118, -0.03528839, 
    -0.03533471, -0.0347929, -0.03496629, -0.03368733, -0.03436961, 
    -0.03245961, -0.03178396, -0.02993589, -0.02884545, -0.02776788, 
    -0.02730224, -0.02716173, -0.02710316,
  -0.01970498, -0.01870054, -0.01889315, -0.01810236, -0.01853836, 
    -0.01802443, -0.01949861, -0.01866132, -0.0191931, -0.01961321, 
    -0.01662923, -0.0180676, -0.01521544, -0.01607415, -0.01397336, 
    -0.01534705, -0.01370618, -0.01401194, -0.01310463, -0.01336067, 
    -0.01224115, -0.0129875, -0.01168477, -0.01241693, -0.01230054, 
    -0.01301258, -0.01777204, -0.01680411, -0.01783047, -0.01769001, 
    -0.01775297, -0.01852925, -0.01892857, -0.01978323, -0.01962626, 
    -0.01899946, -0.01762709, -0.01808556, -0.01694474, -0.01696998, 
    -0.01575423, -0.01629523, -0.01433699, -0.01487744, -0.01334993, 
    -0.01372429, -0.01336735, -0.01347497, -0.01336595, -0.01391764, 
    -0.01367955, -0.01417136, -0.016193, -0.01558102, -0.01745117, 
    -0.01864188, -0.01946137, -0.02005681, -0.01997192, -0.01981072, 
    -0.01899583, -0.01824993, -0.01769438, -0.01732891, -0.01697361, 
    -0.01592645, -0.01538954, -0.0142292, -0.01443443, -0.0140879, 
    -0.01376189, -0.01322518, -0.01331261, -0.01307941, -0.01409703, 
    -0.01341536, -0.01455215, -0.01423542, -0.01687751, -0.01796114, 
    -0.01843468, -0.01885602, -0.0199068, -0.01917717, -0.01946267, 
    -0.01878802, -0.01836728, -0.01857461, -0.01731899, -0.01780039, 
    -0.01535808, -0.01638183, -0.01379967, -0.01439216, -0.01365998, 
    -0.0140306, -0.01339934, -0.01396665, -0.0129933, -0.01278713, 
    -0.01292779, -0.01239279, -0.01399853, -0.01336732, -0.01858043, 
    -0.0185465, -0.01838901, -0.0190878, -0.01913112, -0.01978753, 
    -0.01920278, -0.01895721, -0.01834311, -0.01798595, -0.01765065, 
    -0.01692765, -0.01614293, -0.01508524, -0.01435328, -0.01387542, 
    -0.01416725, -0.0139094, -0.01419783, -0.01433431, -0.01286412, 
    -0.01367732, -0.01246887, -0.01253393, -0.01307388, -0.01252659, 
    -0.01852271, -0.01871832, -0.01940775, -0.01886683, -0.01985989, 
    -0.01929989, -0.01898258, -0.01779017, -0.01753494, -0.01730028, 
    -0.01684286, -0.01626726, -0.01528814, -0.01446743, -0.01374308, 
    -0.01379537, -0.01377694, -0.01361804, -0.01401373, -0.01355376, 
    -0.01347748, -0.01367746, -0.01254266, -0.0128606, -0.01253532, 
    -0.0127417, -0.01865459, -0.01832696, -0.01850353, -0.01817239, 
    -0.01840525, -0.01738434, -0.01708553, -0.01573118, -0.01627845, 
    -0.01541315, -0.0161892, -0.01604989, -0.0153853, -0.01614666, 
    -0.01451188, -0.01560796, -0.01361189, -0.01466344, -0.01354762, 
    -0.01374616, -0.01341845, -0.01312911, -0.01277075, -0.01212558, 
    -0.01227314, -0.01174553, -0.01784551, -0.01743328, -0.01746939, 
    -0.01704408, -0.01673384, -0.01607397, -0.01505064, -0.01543046, 
    -0.01473782, -0.01460118, -0.01565532, -0.01500252, -0.0171609, 
    -0.01679951, -0.01701413, -0.01781273, -0.01534232, -0.01658061, 
    -0.01434136, -0.014977, -0.01317011, -0.01405037, -0.01235483, 
    -0.01167095, -0.01104943, -0.01034922, -0.01721098, -0.0174881, 
    -0.01699397, -0.0163251, -0.01571995, -0.01493772, -0.01485914, 
    -0.01471587, -0.0143489, -0.01404485, -0.0146707, -0.01396927, 
    -0.01671627, -0.01523773, -0.01759356, -0.01686122, -0.01636408, 
    -0.01658105, -0.01547426, -0.01522044, -0.01421619, -0.01472995, 
    -0.01183745, -0.01306842, -0.009834968, -0.01068182, -0.01758559, 
    -0.01721196, -0.01595132, -0.01654349, -0.01488643, -0.01449544, 
    -0.01418246, -0.01378855, -0.01374648, -0.01351682, -0.01389443, 
    -0.01353163, -0.01493608, -0.01429766, -0.0160924, -0.01564309, 
    -0.0158488, -0.01607637, -0.01538063, -0.0146607, -0.01464565, 
    -0.01441954, -0.01379411, -0.01487995, -0.0116839, -0.01360027, 
    -0.01681039, -0.0161157, -0.01601812, -0.01628395, -0.01453434, 
    -0.0151537, -0.0135224, -0.01395178, -0.01325267, -0.01359724, 
    -0.0136484, -0.01410022, -0.01438618, -0.01512493, -0.01574344, 
    -0.01624523, -0.01612766, -0.01557956, -0.01461739, -0.01374263, 
    -0.01393133, -0.01330501, -0.01500286, -0.01427521, -0.01455371, 
    -0.01383464, -0.01544061, -0.01406575, -0.01580513, -0.01564748, 
    -0.01516616, -0.01422662, -0.014024, -0.0138095, -0.01394163, 
    -0.01459349, -0.01470212, -0.01517777, -0.01531075, -0.01568172, 
    -0.0159931, -0.01570843, -0.01541295, -0.01459324, -0.01387859, 
    -0.01312501, -0.01294462, -0.01210438, -0.01278559, -0.01167372, 
    -0.01261482, -0.01101419, -0.01398868, -0.01264336, -0.01514452, 
    -0.01486133, -0.01435758, -0.0132434, -0.01383797, -0.01314428, 
    -0.01470639, -0.01556082, -0.01578701, -0.01621442, -0.01577733, 
    -0.0158126, -0.01540086, -0.01553242, -0.01456652, -0.01508047, 
    -0.01364966, -0.01314969, -0.01180012, -0.01101715, -0.01025401, 
    -0.009927696, -0.009829662, -0.009788851,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  297.9075, 299.1678, 298.9225, 299.9397, 299.3759, 300.0412, 298.1628, 
    299.2177, 298.544, 298.0209, 301.9109, 299.985, 303.923, 302.687, 
    305.7948, 303.7302, 306.206, 305.7363, 307.1524, 306.7462, 308.5623, 
    307.34, 309.5076, 308.2702, 308.4634, 307.2997, 300.3721, 301.6705, 
    300.2952, 300.4801, 300.3972, 299.3875, 298.8771, 297.8115, 298.0048, 
    298.7877, 300.5632, 299.9619, 301.4799, 301.4455, 303.1422, 302.3763, 
    305.2393, 304.4235, 306.7632, 306.1783, 306.7356, 306.5666, 306.7378, 
    305.8805, 306.2476, 305.4933, 302.5195, 303.3911, 300.7971, 299.2422, 
    298.2089, 297.4771, 297.5805, 297.7776, 298.7923, 299.7488, 300.4746, 
    300.9608, 301.4406, 302.8955, 303.6685, 305.4043, 305.0908, 305.6201, 
    306.1202, 306.9603, 306.822, 307.1925, 305.6064, 306.6599, 304.9122, 
    305.3951, 301.57, 300.1241, 299.5089, 298.9696, 297.66, 298.5638, 
    298.2072, 299.0563, 299.5967, 299.3294, 300.9742, 300.3348, 303.7144, 
    302.2551, 306.0619, 305.1552, 306.278, 305.7079, 306.6851, 305.8056, 
    307.3306, 307.6633, 307.4359, 308.3105, 305.7569, 306.7355, 299.3219, 
    299.3654, 299.5686, 298.6762, 298.6217, 297.8062, 298.5319, 298.8412, 
    299.6281, 300.0916, 300.5323, 301.503, 302.5898, 304.1149, 305.2145, 
    305.9454, 305.4997, 305.8933, 305.453, 305.2436, 307.5385, 306.2509, 
    308.1846, 308.0774, 307.2013, 308.0895, 299.3961, 299.1453, 298.2757, 
    298.9561, 297.7175, 298.4102, 298.809, 300.3479, 300.6859, 300.9991, 
    301.6188, 302.4154, 303.8168, 305.0404, 306.1494, 306.0687, 306.097, 
    306.3432, 305.7337, 306.4433, 306.5624, 306.2509, 308.063, 307.5445, 
    308.0751, 307.7374, 299.2268, 299.649, 299.4208, 299.8491, 299.5475, 
    300.8862, 301.2881, 303.1748, 302.3997, 303.6343, 302.525, 302.7213, 
    303.6742, 302.5849, 304.9726, 303.3518, 306.3527, 304.7433, 306.4529, 
    306.1446, 306.6553, 307.1132, 307.6901, 308.7566, 308.5095, 309.4032, 
    300.2755, 300.821, 300.7731, 301.3448, 301.7681, 302.6874, 304.1662, 
    303.6096, 304.6324, 304.838, 303.2844, 304.2373, 301.1866, 301.6776, 
    301.3853, 300.3185, 303.7375, 301.9789, 305.2326, 304.2754, 307.0478, 
    305.6773, 308.3734, 309.531, 310.6245, 311.9051, 301.1192, 300.7482, 
    301.4129, 302.3341, 303.1914, 304.3336, 304.4508, 304.6652, 305.2213, 
    305.6862, 304.7328, 305.8016, 301.7912, 303.8906, 300.6078, 301.5931, 
    302.2798, 301.9786, 303.546, 303.9163, 305.4244, 304.6442, 309.2448, 
    307.2097, 312.8836, 311.2897, 300.6186, 301.118, 302.8609, 302.0307, 
    304.4102, 304.998, 305.4766, 306.0789, 306.1441, 306.5009, 305.9163, 
    306.4779, 304.3361, 305.2996, 302.6615, 303.3018, 303.0072, 302.6841, 
    303.6821, 304.7478, 304.7709, 305.1133, 306.0687, 304.4198, 309.5076, 
    306.3693, 301.6633, 302.628, 302.7664, 302.3922, 304.939, 304.0142, 
    306.4923, 305.8284, 306.9169, 306.3756, 306.296, 305.6016, 305.1642, 
    304.0565, 303.1576, 302.4465, 302.6117, 303.3933, 304.8132, 306.1498, 
    305.8593, 306.834, 304.2371, 305.3338, 304.9095, 306.0081, 303.5947, 
    305.6527, 303.0696, 303.2957, 303.9959, 305.4081, 305.718, 306.0466, 
    305.8439, 304.8493, 304.6858, 303.9789, 303.7838, 303.2465, 302.802, 
    303.208, 303.6348, 304.8499, 305.9403, 307.1196, 307.4089, 308.7915, 
    307.6652, 309.5251, 307.9426, 310.6863, 305.7711, 307.8968, 304.0279, 
    304.4476, 305.2075, 306.9309, 306.0029, 307.0886, 304.6794, 303.4202, 
    303.0954, 302.4896, 303.1093, 303.0589, 303.6527, 303.4618, 304.8903, 
    304.1223, 306.2939, 307.0801, 309.3093, 310.6819, 312.0844, 312.705, 
    312.8941, 312.9731 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.359073e-08, 6.38703e-08, 6.381595e-08, 6.404144e-08, 6.391635e-08, 
    6.406401e-08, 6.364741e-08, 6.38814e-08, 6.373202e-08, 6.361589e-08, 
    6.447906e-08, 6.405151e-08, 6.492314e-08, 6.465046e-08, 6.533541e-08, 
    6.488071e-08, 6.542709e-08, 6.532228e-08, 6.563771e-08, 6.554734e-08, 
    6.595081e-08, 6.567942e-08, 6.615994e-08, 6.588599e-08, 6.592885e-08, 
    6.567046e-08, 6.413754e-08, 6.442583e-08, 6.412046e-08, 6.416157e-08, 
    6.414312e-08, 6.391894e-08, 6.380597e-08, 6.356935e-08, 6.36123e-08, 
    6.37861e-08, 6.418006e-08, 6.404632e-08, 6.438335e-08, 6.437574e-08, 
    6.475095e-08, 6.458178e-08, 6.521241e-08, 6.503318e-08, 6.555111e-08, 
    6.542086e-08, 6.5545e-08, 6.550735e-08, 6.554549e-08, 6.535446e-08, 
    6.54363e-08, 6.52682e-08, 6.461346e-08, 6.480589e-08, 6.423198e-08, 
    6.388689e-08, 6.365767e-08, 6.349501e-08, 6.3518e-08, 6.356184e-08, 
    6.378711e-08, 6.39989e-08, 6.41603e-08, 6.426826e-08, 6.437465e-08, 
    6.469666e-08, 6.486707e-08, 6.524866e-08, 6.517979e-08, 6.529645e-08, 
    6.54079e-08, 6.559502e-08, 6.556422e-08, 6.564666e-08, 6.529337e-08, 
    6.552817e-08, 6.514056e-08, 6.524657e-08, 6.440359e-08, 6.408239e-08, 
    6.39459e-08, 6.38264e-08, 6.353569e-08, 6.373644e-08, 6.36573e-08, 
    6.384558e-08, 6.396522e-08, 6.390604e-08, 6.427122e-08, 6.412925e-08, 
    6.487718e-08, 6.455502e-08, 6.53949e-08, 6.519392e-08, 6.544307e-08, 
    6.531594e-08, 6.553378e-08, 6.533772e-08, 6.567733e-08, 6.575129e-08, 
    6.570075e-08, 6.589487e-08, 6.532685e-08, 6.5545e-08, 6.390439e-08, 
    6.391404e-08, 6.395899e-08, 6.376138e-08, 6.374928e-08, 6.356817e-08, 
    6.372932e-08, 6.379795e-08, 6.397214e-08, 6.407519e-08, 6.417314e-08, 
    6.43885e-08, 6.462902e-08, 6.496534e-08, 6.520695e-08, 6.536891e-08, 
    6.52696e-08, 6.535728e-08, 6.525926e-08, 6.521332e-08, 6.572358e-08, 
    6.543706e-08, 6.586696e-08, 6.584317e-08, 6.564862e-08, 6.584585e-08, 
    6.392082e-08, 6.386528e-08, 6.367247e-08, 6.382336e-08, 6.354846e-08, 
    6.370234e-08, 6.379082e-08, 6.413222e-08, 6.420723e-08, 6.427678e-08, 
    6.441415e-08, 6.459044e-08, 6.489969e-08, 6.516876e-08, 6.541438e-08, 
    6.539639e-08, 6.540272e-08, 6.54576e-08, 6.532167e-08, 6.547991e-08, 
    6.550647e-08, 6.543703e-08, 6.583998e-08, 6.572486e-08, 6.584266e-08, 
    6.57677e-08, 6.388333e-08, 6.397677e-08, 6.392628e-08, 6.402123e-08, 
    6.395434e-08, 6.425178e-08, 6.434096e-08, 6.475822e-08, 6.458697e-08, 
    6.485951e-08, 6.461465e-08, 6.465804e-08, 6.486842e-08, 6.462788e-08, 
    6.515393e-08, 6.47973e-08, 6.545973e-08, 6.510361e-08, 6.548205e-08, 
    6.541332e-08, 6.55271e-08, 6.562901e-08, 6.575721e-08, 6.599377e-08, 
    6.593899e-08, 6.613681e-08, 6.411607e-08, 6.423728e-08, 6.42266e-08, 
    6.435343e-08, 6.444724e-08, 6.465053e-08, 6.49766e-08, 6.485399e-08, 
    6.507909e-08, 6.512427e-08, 6.478229e-08, 6.499227e-08, 6.431839e-08, 
    6.442727e-08, 6.436243e-08, 6.412564e-08, 6.488224e-08, 6.449396e-08, 
    6.521095e-08, 6.500061e-08, 6.561448e-08, 6.530919e-08, 6.590884e-08, 
    6.616519e-08, 6.640643e-08, 6.668839e-08, 6.430341e-08, 6.422106e-08, 
    6.436851e-08, 6.457253e-08, 6.47618e-08, 6.501344e-08, 6.503917e-08, 
    6.508632e-08, 6.520843e-08, 6.531109e-08, 6.510123e-08, 6.533683e-08, 
    6.445253e-08, 6.491594e-08, 6.418993e-08, 6.440856e-08, 6.45605e-08, 
    6.449384e-08, 6.483997e-08, 6.492154e-08, 6.525305e-08, 6.508168e-08, 
    6.610193e-08, 6.565055e-08, 6.690304e-08, 6.655304e-08, 6.419229e-08, 
    6.430313e-08, 6.468889e-08, 6.450534e-08, 6.503023e-08, 6.515943e-08, 
    6.526445e-08, 6.539872e-08, 6.541321e-08, 6.549276e-08, 6.53624e-08, 
    6.54876e-08, 6.501397e-08, 6.522563e-08, 6.464479e-08, 6.478616e-08, 
    6.472112e-08, 6.464978e-08, 6.486996e-08, 6.510454e-08, 6.510954e-08, 
    6.518476e-08, 6.539673e-08, 6.503235e-08, 6.61602e-08, 6.546369e-08, 
    6.442399e-08, 6.46375e-08, 6.466798e-08, 6.458527e-08, 6.514647e-08, 
    6.494314e-08, 6.549082e-08, 6.53428e-08, 6.558533e-08, 6.546481e-08, 
    6.544708e-08, 6.529229e-08, 6.519593e-08, 6.495246e-08, 6.475436e-08, 
    6.459727e-08, 6.46338e-08, 6.480636e-08, 6.511888e-08, 6.541453e-08, 
    6.534977e-08, 6.556689e-08, 6.499217e-08, 6.523317e-08, 6.514002e-08, 
    6.538289e-08, 6.485072e-08, 6.530392e-08, 6.473489e-08, 6.478478e-08, 
    6.49391e-08, 6.524952e-08, 6.531818e-08, 6.539152e-08, 6.534626e-08, 
    6.512681e-08, 6.509086e-08, 6.493535e-08, 6.489241e-08, 6.477391e-08, 
    6.467581e-08, 6.476544e-08, 6.485958e-08, 6.51269e-08, 6.536781e-08, 
    6.563047e-08, 6.569473e-08, 6.600164e-08, 6.575182e-08, 6.616408e-08, 
    6.58136e-08, 6.642029e-08, 6.533017e-08, 6.580328e-08, 6.494612e-08, 
    6.503846e-08, 6.520549e-08, 6.558857e-08, 6.538175e-08, 6.562362e-08, 
    6.508945e-08, 6.481232e-08, 6.47406e-08, 6.460682e-08, 6.474366e-08, 
    6.473253e-08, 6.486347e-08, 6.482139e-08, 6.513578e-08, 6.49669e-08, 
    6.544663e-08, 6.562171e-08, 6.611609e-08, 6.641916e-08, 6.672765e-08, 
    6.686385e-08, 6.690531e-08, 6.692264e-08 ;

 SOM_C_LEACHED =
  -2.580915e-20, 5.488722e-21, 2.163574e-20, 4.52675e-20, -2.863905e-20, 
    1.497707e-20, 3.979948e-20, 5.936901e-20, -4.64529e-21, 1.430571e-20, 
    1.07572e-21, -9.29276e-20, 3.652199e-20, -9.097889e-21, -1.874964e-20, 
    -1.849422e-21, -7.956211e-21, -2.371593e-21, 2.583996e-20, 1.409271e-20, 
    -2.409642e-20, -1.040429e-20, 1.42148e-20, 6.039679e-20, 4.096204e-20, 
    -4.649275e-20, 4.076069e-20, 1.361194e-20, -1.049523e-19, 5.166292e-20, 
    5.112202e-20, 4.576502e-20, -2.049144e-20, -4.889231e-21, -2.916979e-20, 
    5.422341e-20, 5.274296e-20, 3.488688e-21, 2.181559e-20, -1.552187e-20, 
    -3.867689e-20, 9.752535e-20, 2.125859e-20, -4.564014e-20, -1.142837e-19, 
    -1.618532e-20, 4.975575e-21, 5.886318e-20, -4.13997e-20, -4.206056e-20, 
    1.269409e-20, -2.396206e-20, 1.251604e-20, 2.82445e-20, 7.768741e-21, 
    1.296333e-19, 6.602652e-20, 2.144505e-20, -8.431332e-20, 5.192204e-21, 
    -3.049297e-20, 2.111274e-20, -3.013636e-20, -2.11216e-20, -6.797484e-20, 
    -4.52306e-20, 2.33276e-20, 2.314317e-20, -4.732538e-20, -1.261311e-20, 
    1.695546e-20, 1.379817e-20, -4.311946e-20, 2.846877e-20, -4.552828e-20, 
    4.18286e-20, 1.070687e-20, 5.106348e-20, 5.79658e-21, -8.225666e-20, 
    3.519009e-20, 1.664342e-20, -5.942192e-20, -2.374379e-20, -3.255773e-21, 
    -2.903132e-21, 1.141106e-21, 3.999945e-20, 5.866729e-20, 4.366009e-20, 
    -4.710246e-21, 2.06427e-20, -2.536508e-20, -1.540324e-20, -9.878145e-21, 
    -1.012701e-19, -7.012542e-21, 4.446194e-20, -2.231333e-20, 3.705577e-20, 
    -1.393824e-22, -1.639307e-20, -2.178692e-20, -6.040975e-20, 2.900924e-20, 
    1.830389e-20, -9.007997e-21, 7.201179e-20, 3.38241e-20, 3.320803e-20, 
    -1.131611e-20, -2.683806e-20, 3.958965e-20, -2.444104e-20, -6.089109e-20, 
    5.014783e-20, -2.738569e-20, -1.241563e-20, 8.024015e-21, -2.4682e-20, 
    -9.451748e-20, -1.319528e-20, -2.585071e-20, -4.703325e-20, 
    -7.796463e-20, -2.748322e-20, 5.227693e-21, -3.486548e-20, -3.866734e-20, 
    1.182518e-21, -1.266809e-21, -3.578021e-20, 1.342963e-20, -8.746621e-21, 
    1.501018e-20, -1.061466e-20, 2.803959e-20, -2.639792e-20, 2.372041e-20, 
    -3.35621e-20, -8.976037e-20, -5.431003e-20, 5.628559e-21, -5.47368e-20, 
    -7.275087e-20, -7.348548e-20, 1.004615e-20, -1.85586e-20, 1.691867e-20, 
    -3.989524e-22, -3.808963e-21, -2.023128e-21, -3.701898e-20, 
    -2.878824e-20, -3.554437e-20, -1.583556e-20, 2.64037e-20, 2.050013e-20, 
    3.303368e-20, -1.582955e-20, -4.364187e-20, -9.35831e-20, -1.017542e-20, 
    8.719139e-20, -4.876127e-20, -1.800497e-20, -6.80586e-20, -5.280279e-20, 
    1.626254e-20, -5.995927e-20, -5.291962e-20, -7.088234e-20, 3.177427e-20, 
    6.071789e-21, -1.011789e-19, 1.717502e-21, 1.906755e-20, -2.128743e-20, 
    -5.411761e-20, -2.018782e-20, -3.687745e-20, 3.228847e-21, 1.753824e-20, 
    8.482334e-22, -3.155767e-20, -8.588705e-20, -2.863254e-20, 2.093249e-20, 
    5.891629e-20, -4.080638e-21, 5.592527e-20, -4.649321e-20, -4.835335e-20, 
    -3.702215e-21, 2.757981e-20, -2.397592e-20, -2.097523e-21, 1.849629e-21, 
    -3.633164e-20, 7.150261e-20, 1.058005e-20, -3.728663e-20, 2.28916e-20, 
    -1.210755e-20, 7.452384e-20, 6.89005e-22, 4.330013e-21, 5.923648e-20, 
    -5.295411e-20, 6.67191e-20, 4.561269e-20, -5.991856e-20, -9.289759e-23, 
    4.184986e-20, 7.519213e-20, 7.891959e-20, -4.885033e-20, -2.341142e-20, 
    3.636769e-20, 7.917817e-21, -9.413319e-20, 1.734892e-20, -4.335985e-20, 
    5.958988e-20, -3.036344e-20, -9.653483e-20, -3.264351e-20, 3.157911e-20, 
    2.40107e-20, 5.873171e-20, 7.04366e-21, 5.823991e-20, 1.51136e-21, 
    2.340235e-22, 2.923403e-20, 1.813896e-20, 1.01311e-20, -9.259736e-20, 
    4.014413e-20, -3.602547e-21, 9.625271e-21, -1.805763e-20, -2.239885e-20, 
    9.120939e-21, -3.045746e-20, 6.158878e-20, 1.764901e-20, 2.733533e-20, 
    2.545497e-20, -1.098022e-20, 1.19751e-20, 3.181844e-20, 4.588969e-21, 
    -5.371735e-20, -3.162706e-20, -3.796944e-20, 2.208542e-21, -4.695412e-21, 
    -3.411539e-20, 3.260274e-20, 2.794853e-20, -9.447879e-21, 2.83923e-20, 
    6.145263e-20, 4.888457e-20, 3.270822e-20, 4.863431e-20, -3.845568e-20, 
    8.844938e-21, 1.049979e-20, 3.056839e-20, 9.754027e-20, -1.150911e-21, 
    1.722967e-20, -1.560409e-20, 5.282847e-20, -5.827559e-20, 4.721832e-22, 
    2.735147e-21, 6.919253e-20, 2.834708e-20, 4.088215e-20, 1.996237e-20, 
    -6.554297e-21, -5.954928e-20, 1.640046e-20, 9.26701e-21, -3.770105e-20, 
    -5.715841e-20, 1.773359e-20, -1.118399e-20, -7.960145e-20, -1.286328e-20, 
    -3.71269e-20, 2.876586e-20, -5.161031e-20, -2.542049e-20, -8.080565e-20, 
    -2.827145e-22, -2.502624e-20, -2.162675e-20, -5.470216e-21, 4.600025e-22, 
    -1.458517e-20, 3.36148e-20, -4.557132e-20, 3.319852e-20, 1.261215e-20, 
    -3.342714e-20, 5.014685e-20, -2.88194e-21, 8.724449e-20, -3.247801e-21, 
    8.750476e-21, 4.456843e-22, -2.805908e-20, -8.397285e-21, -1.000506e-20, 
    -1.27163e-22, 5.274863e-20, 1.280756e-20, -4.538496e-20, 9.185736e-21, 
    -5.602072e-20, 6.778697e-21, 1.251619e-20, -4.331454e-20, -3.844122e-20, 
    8.588146e-21, -8.662836e-21, -2.986373e-20, -7.120203e-20, -2.581071e-20, 
    1.399998e-20, 3.498347e-21, -6.87128e-21, 3.653643e-21, 4.162553e-20 ;

 SR =
  6.359163e-08, 6.387121e-08, 6.381686e-08, 6.404235e-08, 6.391726e-08, 
    6.406492e-08, 6.364831e-08, 6.388231e-08, 6.373293e-08, 6.36168e-08, 
    6.447997e-08, 6.405241e-08, 6.492405e-08, 6.465138e-08, 6.533632e-08, 
    6.488163e-08, 6.542801e-08, 6.53232e-08, 6.563863e-08, 6.554826e-08, 
    6.595173e-08, 6.568033e-08, 6.616087e-08, 6.588692e-08, 6.592978e-08, 
    6.567138e-08, 6.413845e-08, 6.442674e-08, 6.412137e-08, 6.416248e-08, 
    6.414403e-08, 6.391985e-08, 6.380688e-08, 6.357025e-08, 6.361321e-08, 
    6.3787e-08, 6.418097e-08, 6.404723e-08, 6.438426e-08, 6.437665e-08, 
    6.475187e-08, 6.458269e-08, 6.521333e-08, 6.503409e-08, 6.555204e-08, 
    6.542178e-08, 6.554592e-08, 6.550827e-08, 6.554641e-08, 6.535537e-08, 
    6.543722e-08, 6.526912e-08, 6.461438e-08, 6.480681e-08, 6.423289e-08, 
    6.38878e-08, 6.365858e-08, 6.349591e-08, 6.351891e-08, 6.356274e-08, 
    6.378801e-08, 6.399981e-08, 6.416121e-08, 6.426918e-08, 6.437556e-08, 
    6.469757e-08, 6.486799e-08, 6.524958e-08, 6.518071e-08, 6.529738e-08, 
    6.540882e-08, 6.559594e-08, 6.556514e-08, 6.564758e-08, 6.529429e-08, 
    6.552909e-08, 6.514148e-08, 6.52475e-08, 6.44045e-08, 6.40833e-08, 
    6.394681e-08, 6.38273e-08, 6.353659e-08, 6.373735e-08, 6.365821e-08, 
    6.384649e-08, 6.396612e-08, 6.390695e-08, 6.427213e-08, 6.413016e-08, 
    6.487809e-08, 6.455593e-08, 6.539582e-08, 6.519484e-08, 6.544399e-08, 
    6.531685e-08, 6.55347e-08, 6.533864e-08, 6.567826e-08, 6.575221e-08, 
    6.570168e-08, 6.58958e-08, 6.532778e-08, 6.554592e-08, 6.39053e-08, 
    6.391495e-08, 6.39599e-08, 6.376228e-08, 6.375019e-08, 6.356908e-08, 
    6.373023e-08, 6.379886e-08, 6.397305e-08, 6.40761e-08, 6.417405e-08, 
    6.438941e-08, 6.462994e-08, 6.496626e-08, 6.520787e-08, 6.536983e-08, 
    6.527052e-08, 6.53582e-08, 6.526018e-08, 6.521424e-08, 6.572451e-08, 
    6.543799e-08, 6.586788e-08, 6.584409e-08, 6.564954e-08, 6.584677e-08, 
    6.392172e-08, 6.386619e-08, 6.367338e-08, 6.382427e-08, 6.354936e-08, 
    6.370324e-08, 6.379173e-08, 6.413313e-08, 6.420814e-08, 6.427769e-08, 
    6.441505e-08, 6.459135e-08, 6.49006e-08, 6.516968e-08, 6.54153e-08, 
    6.539731e-08, 6.540364e-08, 6.545852e-08, 6.53226e-08, 6.548083e-08, 
    6.550739e-08, 6.543795e-08, 6.58409e-08, 6.572579e-08, 6.584358e-08, 
    6.576862e-08, 6.388424e-08, 6.397768e-08, 6.392719e-08, 6.402214e-08, 
    6.395525e-08, 6.425269e-08, 6.434187e-08, 6.475913e-08, 6.458788e-08, 
    6.486043e-08, 6.461556e-08, 6.465896e-08, 6.486933e-08, 6.462879e-08, 
    6.515485e-08, 6.479821e-08, 6.546065e-08, 6.510453e-08, 6.548296e-08, 
    6.541424e-08, 6.552803e-08, 6.562993e-08, 6.575814e-08, 6.59947e-08, 
    6.593991e-08, 6.613774e-08, 6.411698e-08, 6.423819e-08, 6.422751e-08, 
    6.435434e-08, 6.444814e-08, 6.465145e-08, 6.497752e-08, 6.485489e-08, 
    6.508e-08, 6.512519e-08, 6.47832e-08, 6.499319e-08, 6.431929e-08, 
    6.442818e-08, 6.436335e-08, 6.412655e-08, 6.488316e-08, 6.449487e-08, 
    6.521186e-08, 6.500152e-08, 6.56154e-08, 6.531011e-08, 6.590976e-08, 
    6.616612e-08, 6.640736e-08, 6.668932e-08, 6.430432e-08, 6.422197e-08, 
    6.436942e-08, 6.457343e-08, 6.476271e-08, 6.501435e-08, 6.504009e-08, 
    6.508724e-08, 6.520934e-08, 6.531201e-08, 6.510215e-08, 6.533775e-08, 
    6.445345e-08, 6.491686e-08, 6.419084e-08, 6.440948e-08, 6.456141e-08, 
    6.449476e-08, 6.484088e-08, 6.492246e-08, 6.525397e-08, 6.50826e-08, 
    6.610285e-08, 6.565147e-08, 6.690398e-08, 6.655396e-08, 6.41932e-08, 
    6.430404e-08, 6.46898e-08, 6.450625e-08, 6.503114e-08, 6.516034e-08, 
    6.526538e-08, 6.539964e-08, 6.541413e-08, 6.549368e-08, 6.536332e-08, 
    6.548853e-08, 6.501489e-08, 6.522654e-08, 6.46457e-08, 6.478708e-08, 
    6.472204e-08, 6.46507e-08, 6.487087e-08, 6.510545e-08, 6.511046e-08, 
    6.518567e-08, 6.539766e-08, 6.503327e-08, 6.616113e-08, 6.546461e-08, 
    6.44249e-08, 6.463841e-08, 6.466889e-08, 6.458619e-08, 6.514739e-08, 
    6.494405e-08, 6.549174e-08, 6.534372e-08, 6.558625e-08, 6.546573e-08, 
    6.5448e-08, 6.529321e-08, 6.519684e-08, 6.495338e-08, 6.475528e-08, 
    6.459818e-08, 6.463471e-08, 6.480727e-08, 6.51198e-08, 6.541545e-08, 
    6.535068e-08, 6.556781e-08, 6.499309e-08, 6.523408e-08, 6.514095e-08, 
    6.538381e-08, 6.485164e-08, 6.530484e-08, 6.47358e-08, 6.47857e-08, 
    6.494002e-08, 6.525044e-08, 6.53191e-08, 6.539243e-08, 6.534718e-08, 
    6.512773e-08, 6.509178e-08, 6.493626e-08, 6.489333e-08, 6.477483e-08, 
    6.467673e-08, 6.476636e-08, 6.486049e-08, 6.512782e-08, 6.536873e-08, 
    6.563138e-08, 6.569566e-08, 6.600256e-08, 6.575274e-08, 6.616501e-08, 
    6.581453e-08, 6.642122e-08, 6.533109e-08, 6.58042e-08, 6.494704e-08, 
    6.503938e-08, 6.520641e-08, 6.558949e-08, 6.538266e-08, 6.562454e-08, 
    6.509037e-08, 6.481324e-08, 6.474151e-08, 6.460773e-08, 6.474458e-08, 
    6.473344e-08, 6.486439e-08, 6.482231e-08, 6.51367e-08, 6.496782e-08, 
    6.544756e-08, 6.562262e-08, 6.611701e-08, 6.642009e-08, 6.672858e-08, 
    6.686479e-08, 6.690624e-08, 6.692357e-08 ;

 STORVEGC =
  0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537 ;

 STORVEGN =
  0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999944, 0.9999943, 
    0.9999943, 0.9999943, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999943, 0.9999942, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999943, 0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999943, 0.9999942, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999944, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999943, 0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999944, 0.9999944, 0.9999944, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999942, 0.9999943, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999944, 0.9999943, 0.9999945, 0.9999944, 
    0.9999942, 0.9999942, 0.9999943, 0.9999942, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999944, 0.9999943, 0.9999942, 0.9999943, 0.9999943, 0.9999942, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999944, 0.9999943, 0.9999944, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999944, 0.9999944, 0.9999944, 0.9999945, 
    0.9999945, 0.9999945 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.1478047, -0.1478197, -0.1478169, -0.1478285, -0.1478223, -0.1478297, 
    -0.1478079, -0.1478202, -0.1478124, -0.1478062, -0.1478488, -0.147829, 
    -0.1478635, -0.147855, -0.1478875, -0.1478622, -0.1478903, -0.1478872, 
    -0.1478969, -0.1478941, -0.1479062, -0.1478982, -0.1479127, -0.1479044, 
    -0.1479056, -0.1478979, -0.1478335, -0.1478469, -0.1478326, -0.1478346, 
    -0.1478337, -0.1478223, -0.1478161, -0.1478038, -0.147806, -0.1478152, 
    -0.1478355, -0.147829, -0.1478458, -0.1478455, -0.1478583, -0.1478529, 
    -0.1478838, -0.147867, -0.1478943, -0.1478903, -0.147894, -0.1478929, 
    -0.1478941, -0.1478882, -0.1478907, -0.1478856, -0.1478538, -0.14786, 
    -0.1478381, -0.1478202, -0.1478084, -0.1477997, -0.147801, -0.1478032, 
    -0.1478152, -0.1478266, -0.1478347, -0.1478401, -0.1478454, -0.1478562, 
    -0.1478619, -0.1478849, -0.1478829, -0.1478864, -0.1478899, -0.1478956, 
    -0.1478946, -0.1478971, -0.1478864, -0.1478935, -0.1478817, -0.1478849, 
    -0.147846, -0.1478308, -0.1478235, -0.1478174, -0.1478019, -0.1478126, 
    -0.1478083, -0.1478186, -0.1478249, -0.1478218, -0.1478402, -0.1478331, 
    -0.1478622, -0.1478519, -0.1478895, -0.1478833, -0.1478909, -0.1478871, 
    -0.1478937, -0.1478877, -0.1478981, -0.1479003, -0.1478988, -0.1479047, 
    -0.1478874, -0.147894, -0.1478217, -0.1478222, -0.1478246, -0.1478139, 
    -0.1478133, -0.1478037, -0.1478123, -0.1478159, -0.1478253, -0.1478304, 
    -0.1478353, -0.147846, -0.1478543, -0.1478648, -0.1478837, -0.1478887, 
    -0.1478857, -0.1478883, -0.1478853, -0.147884, -0.1478994, -0.1478907, 
    -0.1479039, -0.1479032, -0.1478971, -0.1479032, -0.1478225, -0.1478196, 
    -0.1478092, -0.1478174, -0.1478026, -0.1478108, -0.1478154, -0.1478331, 
    -0.147837, -0.1478404, -0.147847, -0.1478531, -0.1478629, -0.1478825, 
    -0.1478901, -0.1478895, -0.1478897, -0.1478914, -0.1478872, -0.1478921, 
    -0.1478928, -0.1478907, -0.1479031, -0.1478996, -0.1479032, -0.1479009, 
    -0.1478206, -0.1478255, -0.1478229, -0.1478276, -0.1478243, -0.147839, 
    -0.1478434, -0.1478584, -0.147853, -0.1478617, -0.1478539, -0.1478553, 
    -0.1478617, -0.1478544, -0.1478819, -0.1478596, -0.1478914, -0.1478688, 
    -0.1478921, -0.14789, -0.1478935, -0.1478966, -0.1479005, -0.1479077, 
    -0.147906, -0.1479121, -0.1478325, -0.1478384, -0.147838, -0.1478443, 
    -0.1478482, -0.1478551, -0.1478652, -0.1478617, -0.1478684, -0.1478812, 
    -0.1478594, -0.1478657, -0.1478425, -0.1478473, -0.1478447, -0.1478328, 
    -0.1478623, -0.1478497, -0.1478838, -0.147866, -0.1478961, -0.1478867, 
    -0.1479051, -0.1479127, -0.1479203, -0.1479287, -0.1478418, -0.1478377, 
    -0.1478451, -0.1478524, -0.1478586, -0.1478663, -0.1478672, -0.1478686, 
    -0.1478838, -0.1478869, -0.1478689, -0.1478877, -0.1478479, -0.1478634, 
    -0.1478361, -0.1478466, -0.1478521, -0.1478499, -0.1478613, -0.1478637, 
    -0.147885, -0.1478685, -0.1479107, -0.1478971, -0.1479354, -0.1479246, 
    -0.1478363, -0.1478418, -0.1478562, -0.1478503, -0.1478669, -0.1478822, 
    -0.1478855, -0.1478895, -0.14789, -0.1478924, -0.1478885, -0.1478923, 
    -0.1478663, -0.1478843, -0.1478549, -0.1478594, -0.1478574, -0.1478551, 
    -0.1478622, -0.1478804, -0.1478807, -0.147883, -0.1478889, -0.1478669, 
    -0.1479122, -0.147891, -0.1478474, -0.1478545, -0.1478556, -0.147853, 
    -0.1478818, -0.1478643, -0.1478924, -0.1478879, -0.1478953, -0.1478916, 
    -0.1478911, -0.1478863, -0.1478834, -0.1478645, -0.1478584, -0.1478534, 
    -0.1478546, -0.1478601, -0.1478809, -0.14789, -0.147888, -0.1478947, 
    -0.1478657, -0.1478844, -0.1478816, -0.1478891, -0.1478615, -0.1478862, 
    -0.1478579, -0.1478595, -0.1478641, -0.1478848, -0.1478871, -0.1478893, 
    -0.147888, -0.1478812, -0.1478687, -0.1478641, -0.1478627, -0.1478591, 
    -0.1478559, -0.1478588, -0.1478617, -0.1478812, -0.1478886, -0.1478966, 
    -0.1478986, -0.1479076, -0.1479001, -0.1479123, -0.1479015, -0.1479203, 
    -0.1478872, -0.1479016, -0.1478644, -0.1478672, -0.1478835, -0.1478952, 
    -0.147889, -0.1478963, -0.1478686, -0.1478602, -0.147858, -0.1478537, 
    -0.1478581, -0.1478578, -0.147862, -0.1478607, -0.1478815, -0.147865, 
    -0.147891, -0.1478963, -0.1479114, -0.1479205, -0.1479302, -0.1479343, 
    -0.1479356, -0.1479361 ;

 TAUY =
  -0.1478047, -0.1478197, -0.1478169, -0.1478285, -0.1478223, -0.1478297, 
    -0.1478079, -0.1478202, -0.1478124, -0.1478062, -0.1478488, -0.147829, 
    -0.1478635, -0.147855, -0.1478875, -0.1478622, -0.1478903, -0.1478872, 
    -0.1478969, -0.1478941, -0.1479062, -0.1478982, -0.1479127, -0.1479044, 
    -0.1479056, -0.1478979, -0.1478335, -0.1478469, -0.1478326, -0.1478346, 
    -0.1478337, -0.1478223, -0.1478161, -0.1478038, -0.147806, -0.1478152, 
    -0.1478355, -0.147829, -0.1478458, -0.1478455, -0.1478583, -0.1478529, 
    -0.1478838, -0.147867, -0.1478943, -0.1478903, -0.147894, -0.1478929, 
    -0.1478941, -0.1478882, -0.1478907, -0.1478856, -0.1478538, -0.14786, 
    -0.1478381, -0.1478202, -0.1478084, -0.1477997, -0.147801, -0.1478032, 
    -0.1478152, -0.1478266, -0.1478347, -0.1478401, -0.1478454, -0.1478562, 
    -0.1478619, -0.1478849, -0.1478829, -0.1478864, -0.1478899, -0.1478956, 
    -0.1478946, -0.1478971, -0.1478864, -0.1478935, -0.1478817, -0.1478849, 
    -0.147846, -0.1478308, -0.1478235, -0.1478174, -0.1478019, -0.1478126, 
    -0.1478083, -0.1478186, -0.1478249, -0.1478218, -0.1478402, -0.1478331, 
    -0.1478622, -0.1478519, -0.1478895, -0.1478833, -0.1478909, -0.1478871, 
    -0.1478937, -0.1478877, -0.1478981, -0.1479003, -0.1478988, -0.1479047, 
    -0.1478874, -0.147894, -0.1478217, -0.1478222, -0.1478246, -0.1478139, 
    -0.1478133, -0.1478037, -0.1478123, -0.1478159, -0.1478253, -0.1478304, 
    -0.1478353, -0.147846, -0.1478543, -0.1478648, -0.1478837, -0.1478887, 
    -0.1478857, -0.1478883, -0.1478853, -0.147884, -0.1478994, -0.1478907, 
    -0.1479039, -0.1479032, -0.1478971, -0.1479032, -0.1478225, -0.1478196, 
    -0.1478092, -0.1478174, -0.1478026, -0.1478108, -0.1478154, -0.1478331, 
    -0.147837, -0.1478404, -0.147847, -0.1478531, -0.1478629, -0.1478825, 
    -0.1478901, -0.1478895, -0.1478897, -0.1478914, -0.1478872, -0.1478921, 
    -0.1478928, -0.1478907, -0.1479031, -0.1478996, -0.1479032, -0.1479009, 
    -0.1478206, -0.1478255, -0.1478229, -0.1478276, -0.1478243, -0.147839, 
    -0.1478434, -0.1478584, -0.147853, -0.1478617, -0.1478539, -0.1478553, 
    -0.1478617, -0.1478544, -0.1478819, -0.1478596, -0.1478914, -0.1478688, 
    -0.1478921, -0.14789, -0.1478935, -0.1478966, -0.1479005, -0.1479077, 
    -0.147906, -0.1479121, -0.1478325, -0.1478384, -0.147838, -0.1478443, 
    -0.1478482, -0.1478551, -0.1478652, -0.1478617, -0.1478684, -0.1478812, 
    -0.1478594, -0.1478657, -0.1478425, -0.1478473, -0.1478447, -0.1478328, 
    -0.1478623, -0.1478497, -0.1478838, -0.147866, -0.1478961, -0.1478867, 
    -0.1479051, -0.1479127, -0.1479203, -0.1479287, -0.1478418, -0.1478377, 
    -0.1478451, -0.1478524, -0.1478586, -0.1478663, -0.1478672, -0.1478686, 
    -0.1478838, -0.1478869, -0.1478689, -0.1478877, -0.1478479, -0.1478634, 
    -0.1478361, -0.1478466, -0.1478521, -0.1478499, -0.1478613, -0.1478637, 
    -0.147885, -0.1478685, -0.1479107, -0.1478971, -0.1479354, -0.1479246, 
    -0.1478363, -0.1478418, -0.1478562, -0.1478503, -0.1478669, -0.1478822, 
    -0.1478855, -0.1478895, -0.14789, -0.1478924, -0.1478885, -0.1478923, 
    -0.1478663, -0.1478843, -0.1478549, -0.1478594, -0.1478574, -0.1478551, 
    -0.1478622, -0.1478804, -0.1478807, -0.147883, -0.1478889, -0.1478669, 
    -0.1479122, -0.147891, -0.1478474, -0.1478545, -0.1478556, -0.147853, 
    -0.1478818, -0.1478643, -0.1478924, -0.1478879, -0.1478953, -0.1478916, 
    -0.1478911, -0.1478863, -0.1478834, -0.1478645, -0.1478584, -0.1478534, 
    -0.1478546, -0.1478601, -0.1478809, -0.14789, -0.147888, -0.1478947, 
    -0.1478657, -0.1478844, -0.1478816, -0.1478891, -0.1478615, -0.1478862, 
    -0.1478579, -0.1478595, -0.1478641, -0.1478848, -0.1478871, -0.1478893, 
    -0.147888, -0.1478812, -0.1478687, -0.1478641, -0.1478627, -0.1478591, 
    -0.1478559, -0.1478588, -0.1478617, -0.1478812, -0.1478886, -0.1478966, 
    -0.1478986, -0.1479076, -0.1479001, -0.1479123, -0.1479015, -0.1479203, 
    -0.1478872, -0.1479016, -0.1478644, -0.1478672, -0.1478835, -0.1478952, 
    -0.147889, -0.1478963, -0.1478686, -0.1478602, -0.147858, -0.1478537, 
    -0.1478581, -0.1478578, -0.147862, -0.1478607, -0.1478815, -0.147865, 
    -0.147891, -0.1478963, -0.1479114, -0.1479205, -0.1479302, -0.1479343, 
    -0.1479356, -0.1479361 ;

 TBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.6572, 261.6737, 261.6705, 261.6837, 261.6764, 261.6851, 261.6606, 
    261.6743, 261.6655, 261.6587, 261.7094, 261.6843, 261.7357, 261.7196, 
    261.7599, 261.7332, 261.7654, 261.7592, 261.7778, 261.7725, 261.7962, 
    261.7803, 261.8086, 261.7924, 261.795, 261.7798, 261.6894, 261.7063, 
    261.6884, 261.6908, 261.6897, 261.6765, 261.6698, 261.656, 261.6585, 
    261.6687, 261.6919, 261.6841, 261.7039, 261.7035, 261.7256, 261.7156, 
    261.7527, 261.7423, 261.7727, 261.765, 261.7723, 261.7701, 261.7724, 
    261.7611, 261.7659, 261.756, 261.7175, 261.7288, 261.695, 261.6746, 
    261.6612, 261.6516, 261.653, 261.6555, 261.6688, 261.6812, 261.6908, 
    261.6971, 261.7034, 261.7223, 261.7324, 261.7548, 261.7508, 261.7577, 
    261.7643, 261.7753, 261.7735, 261.7784, 261.7575, 261.7713, 261.7485, 
    261.7547, 261.7049, 261.6862, 261.6781, 261.6711, 261.654, 261.6658, 
    261.6611, 261.6722, 261.6793, 261.6758, 261.6973, 261.6889, 261.733, 
    261.714, 261.7635, 261.7516, 261.7663, 261.7589, 261.7717, 261.7601, 
    261.7802, 261.7845, 261.7815, 261.793, 261.7595, 261.7723, 261.6757, 
    261.6763, 261.6789, 261.6672, 261.6665, 261.6559, 261.6654, 261.6694, 
    261.6797, 261.6857, 261.6915, 261.7042, 261.7184, 261.7382, 261.7524, 
    261.762, 261.7561, 261.7613, 261.7555, 261.7528, 261.7829, 261.766, 
    261.7914, 261.7899, 261.7784, 261.7901, 261.6767, 261.6734, 261.662, 
    261.6709, 261.6548, 261.6638, 261.669, 261.6891, 261.6935, 261.6976, 
    261.7057, 261.7161, 261.7343, 261.7501, 261.7646, 261.7636, 261.7639, 
    261.7672, 261.7592, 261.7685, 261.7701, 261.766, 261.7898, 261.783, 
    261.7899, 261.7855, 261.6745, 261.68, 261.677, 261.6826, 261.6786, 
    261.6961, 261.7014, 261.726, 261.7159, 261.732, 261.7175, 261.7201, 
    261.7324, 261.7183, 261.7492, 261.7283, 261.7673, 261.7463, 261.7686, 
    261.7646, 261.7713, 261.7773, 261.7849, 261.7988, 261.7956, 261.8073, 
    261.6882, 261.6953, 261.6947, 261.7021, 261.7076, 261.7197, 261.7389, 
    261.7317, 261.745, 261.7475, 261.7274, 261.7398, 261.7, 261.7064, 
    261.7026, 261.6887, 261.7333, 261.7104, 261.7526, 261.7403, 261.7764, 
    261.7584, 261.7938, 261.8089, 261.8232, 261.8397, 261.6992, 261.6943, 
    261.703, 261.715, 261.7262, 261.7411, 261.7426, 261.7454, 261.7525, 
    261.7585, 261.7462, 261.7601, 261.7079, 261.7353, 261.6925, 261.7053, 
    261.7143, 261.7104, 261.7309, 261.7357, 261.7551, 261.7451, 261.8051, 
    261.7785, 261.8524, 261.8318, 261.6927, 261.6992, 261.7219, 261.7111, 
    261.7421, 261.7496, 261.7558, 261.7637, 261.7646, 261.7693, 261.7616, 
    261.769, 261.7411, 261.7535, 261.7193, 261.7277, 261.7238, 261.7196, 
    261.7326, 261.7463, 261.7466, 261.7511, 261.7634, 261.7422, 261.8085, 
    261.7674, 261.7063, 261.7188, 261.7207, 261.7158, 261.7488, 261.7369, 
    261.7692, 261.7604, 261.7747, 261.7676, 261.7666, 261.7574, 261.7517, 
    261.7375, 261.7258, 261.7165, 261.7187, 261.7289, 261.7472, 261.7646, 
    261.7608, 261.7737, 261.7398, 261.7539, 261.7484, 261.7628, 261.7315, 
    261.758, 261.7247, 261.7276, 261.7367, 261.7549, 261.759, 261.7633, 
    261.7606, 261.7477, 261.7457, 261.7365, 261.7339, 261.727, 261.7212, 
    261.7264, 261.732, 261.7477, 261.7619, 261.7774, 261.7812, 261.7992, 
    261.7845, 261.8087, 261.788, 261.8239, 261.7596, 261.7875, 261.7371, 
    261.7426, 261.7523, 261.7749, 261.7627, 261.7769, 261.7456, 261.7292, 
    261.725, 261.7171, 261.7252, 261.7245, 261.7322, 261.7298, 261.7482, 
    261.7383, 261.7665, 261.7769, 261.806, 261.8239, 261.8421, 261.8501, 
    261.8526, 261.8536 ;

 TG_R =
  261.6572, 261.6737, 261.6705, 261.6837, 261.6764, 261.6851, 261.6606, 
    261.6743, 261.6655, 261.6587, 261.7094, 261.6843, 261.7357, 261.7196, 
    261.7599, 261.7332, 261.7654, 261.7592, 261.7778, 261.7725, 261.7962, 
    261.7803, 261.8086, 261.7924, 261.795, 261.7798, 261.6894, 261.7063, 
    261.6884, 261.6908, 261.6897, 261.6765, 261.6698, 261.656, 261.6585, 
    261.6687, 261.6919, 261.6841, 261.7039, 261.7035, 261.7256, 261.7156, 
    261.7527, 261.7423, 261.7727, 261.765, 261.7723, 261.7701, 261.7724, 
    261.7611, 261.7659, 261.756, 261.7175, 261.7288, 261.695, 261.6746, 
    261.6612, 261.6516, 261.653, 261.6555, 261.6688, 261.6812, 261.6908, 
    261.6971, 261.7034, 261.7223, 261.7324, 261.7548, 261.7508, 261.7577, 
    261.7643, 261.7753, 261.7735, 261.7784, 261.7575, 261.7713, 261.7485, 
    261.7547, 261.7049, 261.6862, 261.6781, 261.6711, 261.654, 261.6658, 
    261.6611, 261.6722, 261.6793, 261.6758, 261.6973, 261.6889, 261.733, 
    261.714, 261.7635, 261.7516, 261.7663, 261.7589, 261.7717, 261.7601, 
    261.7802, 261.7845, 261.7815, 261.793, 261.7595, 261.7723, 261.6757, 
    261.6763, 261.6789, 261.6672, 261.6665, 261.6559, 261.6654, 261.6694, 
    261.6797, 261.6857, 261.6915, 261.7042, 261.7184, 261.7382, 261.7524, 
    261.762, 261.7561, 261.7613, 261.7555, 261.7528, 261.7829, 261.766, 
    261.7914, 261.7899, 261.7784, 261.7901, 261.6767, 261.6734, 261.662, 
    261.6709, 261.6548, 261.6638, 261.669, 261.6891, 261.6935, 261.6976, 
    261.7057, 261.7161, 261.7343, 261.7501, 261.7646, 261.7636, 261.7639, 
    261.7672, 261.7592, 261.7685, 261.7701, 261.766, 261.7898, 261.783, 
    261.7899, 261.7855, 261.6745, 261.68, 261.677, 261.6826, 261.6786, 
    261.6961, 261.7014, 261.726, 261.7159, 261.732, 261.7175, 261.7201, 
    261.7324, 261.7183, 261.7492, 261.7283, 261.7673, 261.7463, 261.7686, 
    261.7646, 261.7713, 261.7773, 261.7849, 261.7988, 261.7956, 261.8073, 
    261.6882, 261.6953, 261.6947, 261.7021, 261.7076, 261.7197, 261.7389, 
    261.7317, 261.745, 261.7475, 261.7274, 261.7398, 261.7, 261.7064, 
    261.7026, 261.6887, 261.7333, 261.7104, 261.7526, 261.7403, 261.7764, 
    261.7584, 261.7938, 261.8089, 261.8232, 261.8397, 261.6992, 261.6943, 
    261.703, 261.715, 261.7262, 261.7411, 261.7426, 261.7454, 261.7525, 
    261.7585, 261.7462, 261.7601, 261.7079, 261.7353, 261.6925, 261.7053, 
    261.7143, 261.7104, 261.7309, 261.7357, 261.7551, 261.7451, 261.8051, 
    261.7785, 261.8524, 261.8318, 261.6927, 261.6992, 261.7219, 261.7111, 
    261.7421, 261.7496, 261.7558, 261.7637, 261.7646, 261.7693, 261.7616, 
    261.769, 261.7411, 261.7535, 261.7193, 261.7277, 261.7238, 261.7196, 
    261.7326, 261.7463, 261.7466, 261.7511, 261.7634, 261.7422, 261.8085, 
    261.7674, 261.7063, 261.7188, 261.7207, 261.7158, 261.7488, 261.7369, 
    261.7692, 261.7604, 261.7747, 261.7676, 261.7666, 261.7574, 261.7517, 
    261.7375, 261.7258, 261.7165, 261.7187, 261.7289, 261.7472, 261.7646, 
    261.7608, 261.7737, 261.7398, 261.7539, 261.7484, 261.7628, 261.7315, 
    261.758, 261.7247, 261.7276, 261.7367, 261.7549, 261.759, 261.7633, 
    261.7606, 261.7477, 261.7457, 261.7365, 261.7339, 261.727, 261.7212, 
    261.7264, 261.732, 261.7477, 261.7619, 261.7774, 261.7812, 261.7992, 
    261.7845, 261.8087, 261.788, 261.8239, 261.7596, 261.7875, 261.7371, 
    261.7426, 261.7523, 261.7749, 261.7627, 261.7769, 261.7456, 261.7292, 
    261.725, 261.7171, 261.7252, 261.7245, 261.7322, 261.7298, 261.7482, 
    261.7383, 261.7665, 261.7769, 261.806, 261.8239, 261.8421, 261.8501, 
    261.8526, 261.8536 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.0227, 254.0245, 254.0242, 254.0256, 254.0248, 254.0258, 254.0231, 
    254.0246, 254.0236, 254.0229, 254.0284, 254.0257, 254.0313, 254.0296, 
    254.034, 254.0311, 254.0346, 254.034, 254.036, 254.0354, 254.038, 
    254.0363, 254.0394, 254.0376, 254.0379, 254.0362, 254.0263, 254.028, 
    254.0262, 254.0264, 254.0263, 254.0248, 254.0241, 254.0226, 254.0229, 
    254.024, 254.0265, 254.0257, 254.0279, 254.0278, 254.0303, 254.0292, 
    254.0332, 254.0321, 254.0355, 254.0346, 254.0354, 254.0352, 254.0354, 
    254.0342, 254.0347, 254.0336, 254.0294, 254.0306, 254.0269, 254.0246, 
    254.0231, 254.0221, 254.0222, 254.0225, 254.024, 254.0254, 254.0264, 
    254.0271, 254.0278, 254.0298, 254.031, 254.0335, 254.0331, 254.0338, 
    254.0345, 254.0357, 254.0355, 254.0361, 254.0338, 254.0353, 254.0328, 
    254.0335, 254.0279, 254.0259, 254.025, 254.0242, 254.0224, 254.0237, 
    254.0231, 254.0244, 254.0252, 254.0248, 254.0271, 254.0262, 254.0311, 
    254.029, 254.0344, 254.0331, 254.0348, 254.0339, 254.0353, 254.0341, 
    254.0363, 254.0367, 254.0364, 254.0377, 254.034, 254.0354, 254.0248, 
    254.0248, 254.0251, 254.0238, 254.0237, 254.0226, 254.0236, 254.0241, 
    254.0252, 254.0259, 254.0265, 254.0279, 254.0294, 254.0316, 254.0332, 
    254.0343, 254.0336, 254.0342, 254.0336, 254.0333, 254.0366, 254.0347, 
    254.0375, 254.0374, 254.0361, 254.0374, 254.0249, 254.0245, 254.0232, 
    254.0242, 254.0224, 254.0234, 254.024, 254.0262, 254.0267, 254.0272, 
    254.0281, 254.0292, 254.0312, 254.033, 254.0346, 254.0345, 254.0345, 
    254.0349, 254.034, 254.035, 254.0352, 254.0347, 254.0373, 254.0366, 
    254.0374, 254.0369, 254.0246, 254.0252, 254.0249, 254.0255, 254.0251, 
    254.027, 254.0276, 254.0303, 254.0292, 254.0309, 254.0294, 254.0296, 
    254.031, 254.0295, 254.0328, 254.0305, 254.0349, 254.0325, 254.035, 
    254.0346, 254.0353, 254.036, 254.0368, 254.0383, 254.038, 254.0393, 
    254.0261, 254.0269, 254.0269, 254.0277, 254.0283, 254.0296, 254.0317, 
    254.0309, 254.0324, 254.0327, 254.0305, 254.0318, 254.0274, 254.0281, 
    254.0277, 254.0262, 254.0311, 254.0286, 254.0332, 254.0319, 254.0359, 
    254.0339, 254.0378, 254.0394, 254.041, 254.0428, 254.0274, 254.0268, 
    254.0278, 254.0291, 254.0303, 254.032, 254.0321, 254.0324, 254.0332, 
    254.0339, 254.0325, 254.0341, 254.0282, 254.0313, 254.0266, 254.028, 
    254.029, 254.0286, 254.0309, 254.0314, 254.0335, 254.0324, 254.039, 
    254.0361, 254.0443, 254.0419, 254.0266, 254.0274, 254.0298, 254.0287, 
    254.0321, 254.0329, 254.0336, 254.0345, 254.0346, 254.0351, 254.0342, 
    254.035, 254.032, 254.0333, 254.0296, 254.0305, 254.0301, 254.0296, 
    254.0311, 254.0325, 254.0326, 254.0331, 254.0343, 254.0321, 254.0393, 
    254.0348, 254.0282, 254.0295, 254.0297, 254.0292, 254.0328, 254.0315, 
    254.0351, 254.0341, 254.0357, 254.0349, 254.0348, 254.0338, 254.0331, 
    254.0316, 254.0303, 254.0293, 254.0295, 254.0306, 254.0326, 254.0346, 
    254.0341, 254.0356, 254.0318, 254.0334, 254.0328, 254.0344, 254.0309, 
    254.0337, 254.0302, 254.0305, 254.0315, 254.0335, 254.034, 254.0344, 
    254.0341, 254.0327, 254.0325, 254.0315, 254.0312, 254.0304, 254.0298, 
    254.0304, 254.031, 254.0327, 254.0343, 254.036, 254.0364, 254.0383, 
    254.0367, 254.0393, 254.037, 254.041, 254.034, 254.037, 254.0315, 
    254.0321, 254.0332, 254.0357, 254.0343, 254.0359, 254.0325, 254.0306, 
    254.0302, 254.0293, 254.0302, 254.0302, 254.031, 254.0307, 254.0327, 
    254.0317, 254.0348, 254.0359, 254.0391, 254.0411, 254.0431, 254.044, 
    254.0443, 254.0444 ;

 THBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23991, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23998, 18.23999, 18.23999, 18.24, 18.23999, 18.23999, 
    18.23997, 18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 
    18.23991, 18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 
    18.23994, 18.23995, 18.23995, 18.23993, 18.23995, 18.23992, 18.23994, 
    18.23991, 18.23992, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 
    18.23988, 18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 
    18.23996, 18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 
    18.23993, 18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 
    18.23992, 18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 
    18.23985, 18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 
    18.23993, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23996, 
    18.23993, 18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 
    18.23992, 18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 
    18.23996, 18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 
    18.23994, 18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23992, 
    18.23991, 18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 
    18.23995, 18.23992, 18.23993, 18.2399, 18.23991, 18.2399, 18.23991, 
    18.23991, 18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 
    18.23994, 18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 
    18.23992, 18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 
    18.23992, 18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 
    18.23993, 18.23994, 18.23994, 18.23994, 18.23994, 18.23992, 18.23991, 
    18.2399, 18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 
    18.23991, 18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 
    18.2399, 18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 
    18.23994, 18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 
    18.23986, 18.23985, 18.23984, 18.23984, 18.23983 ;

 TOTCOLCH4 =
  1.384702e-05, 1.376081e-05, 1.377745e-05, 1.370882e-05, 1.374677e-05, 
    1.370201e-05, 1.382942e-05, 1.375742e-05, 1.380326e-05, 1.383921e-05, 
    1.357851e-05, 1.370578e-05, 1.35267e-05, 1.361748e-05, 1.339417e-05, 
    1.354064e-05, 1.336547e-05, 1.339832e-05, 1.330058e-05, 1.332825e-05, 
    1.320669e-05, 1.32879e-05, 1.314575e-05, 1.322589e-05, 1.321319e-05, 
    1.329062e-05, 1.367989e-05, 1.359415e-05, 1.368502e-05, 1.367268e-05, 
    1.367822e-05, 1.374598e-05, 1.378049e-05, 1.385369e-05, 1.384032e-05, 
    1.378661e-05, 1.366714e-05, 1.370736e-05, 1.360674e-05, 1.360898e-05, 
    1.358374e-05, 1.364075e-05, 1.343314e-05, 1.34908e-05, 1.332709e-05, 
    1.336743e-05, 1.332897e-05, 1.334058e-05, 1.332882e-05, 1.33882e-05, 
    1.336261e-05, 1.341541e-05, 1.363e-05, 1.356543e-05, 1.365164e-05, 
    1.375572e-05, 1.382624e-05, 1.387691e-05, 1.386972e-05, 1.385602e-05, 
    1.37863e-05, 1.37217e-05, 1.367307e-05, 1.364084e-05, 1.360931e-05, 
    1.360189e-05, 1.354515e-05, 1.342159e-05, 1.344355e-05, 1.340646e-05, 
    1.337147e-05, 1.331361e-05, 1.332306e-05, 1.329785e-05, 1.340745e-05, 
    1.333414e-05, 1.345613e-05, 1.342227e-05, 1.360069e-05, 1.369648e-05, 
    1.373775e-05, 1.377425e-05, 1.386419e-05, 1.380189e-05, 1.382635e-05, 
    1.376838e-05, 1.373191e-05, 1.374992e-05, 1.363996e-05, 1.368239e-05, 
    1.354182e-05, 1.364984e-05, 1.337553e-05, 1.343904e-05, 1.336051e-05, 
    1.340033e-05, 1.333242e-05, 1.339347e-05, 1.328852e-05, 1.326616e-05, 
    1.328142e-05, 1.322327e-05, 1.339689e-05, 1.332896e-05, 1.375042e-05, 
    1.374748e-05, 1.373381e-05, 1.379421e-05, 1.379794e-05, 1.385405e-05, 
    1.380409e-05, 1.378297e-05, 1.372982e-05, 1.369865e-05, 1.366922e-05, 
    1.360521e-05, 1.362472e-05, 1.351288e-05, 1.343488e-05, 1.338367e-05, 
    1.341497e-05, 1.338732e-05, 1.341825e-05, 1.343285e-05, 1.327451e-05, 
    1.336237e-05, 1.323156e-05, 1.323864e-05, 1.329725e-05, 1.323784e-05, 
    1.374542e-05, 1.376236e-05, 1.382165e-05, 1.377519e-05, 1.386021e-05, 
    1.381242e-05, 1.378515e-05, 1.368148e-05, 1.365903e-05, 1.36383e-05, 
    1.359765e-05, 1.363781e-05, 1.353442e-05, 1.344707e-05, 1.336945e-05, 
    1.337507e-05, 1.337309e-05, 1.335599e-05, 1.339852e-05, 1.334907e-05, 
    1.334084e-05, 1.336239e-05, 1.323959e-05, 1.327414e-05, 1.323879e-05, 
    1.326124e-05, 1.375685e-05, 1.372841e-05, 1.374375e-05, 1.371494e-05, 
    1.373521e-05, 1.364572e-05, 1.361924e-05, 1.35813e-05, 1.363898e-05, 
    1.354766e-05, 1.36296e-05, 1.361493e-05, 1.354469e-05, 1.362512e-05, 
    1.345181e-05, 1.356827e-05, 1.335533e-05, 1.346797e-05, 1.334841e-05, 
    1.336978e-05, 1.333449e-05, 1.330323e-05, 1.326439e-05, 1.319408e-05, 
    1.321021e-05, 1.315243e-05, 1.368635e-05, 1.365005e-05, 1.365325e-05, 
    1.361557e-05, 1.358791e-05, 1.361747e-05, 1.350921e-05, 1.354951e-05, 
    1.347593e-05, 1.346136e-05, 1.35733e-05, 1.350409e-05, 1.362594e-05, 
    1.359377e-05, 1.361291e-05, 1.368346e-05, 1.354015e-05, 1.357418e-05, 
    1.34336e-05, 1.350138e-05, 1.330766e-05, 1.340243e-05, 1.321912e-05, 
    1.314421e-05, 1.307563e-05, 1.299758e-05, 1.363039e-05, 1.365491e-05, 
    1.361112e-05, 1.364388e-05, 1.358012e-05, 1.34972e-05, 1.348885e-05, 
    1.347359e-05, 1.343442e-05, 1.340186e-05, 1.346876e-05, 1.339375e-05, 
    1.358631e-05, 1.352907e-05, 1.366419e-05, 1.359927e-05, 1.364798e-05, 
    1.357423e-05, 1.355415e-05, 1.352725e-05, 1.34202e-05, 1.347509e-05, 
    1.31625e-05, 1.329664e-05, 1.293972e-05, 1.303475e-05, 1.36635e-05, 
    1.363048e-05, 1.360454e-05, 1.357087e-05, 1.349175e-05, 1.345007e-05, 
    1.34166e-05, 1.337433e-05, 1.336982e-05, 1.334509e-05, 1.338571e-05, 
    1.334669e-05, 1.349703e-05, 1.342893e-05, 1.361941e-05, 1.3572e-05, 
    1.359373e-05, 1.361773e-05, 1.354423e-05, 1.346769e-05, 1.34661e-05, 
    1.344196e-05, 1.337488e-05, 1.349106e-05, 1.31456e-05, 1.335403e-05, 
    1.359476e-05, 1.362185e-05, 1.361158e-05, 1.363957e-05, 1.345422e-05, 
    1.352016e-05, 1.334569e-05, 1.339187e-05, 1.331659e-05, 1.335376e-05, 
    1.335926e-05, 1.340779e-05, 1.34384e-05, 1.35171e-05, 1.35826e-05, 
    1.36355e-05, 1.362313e-05, 1.356528e-05, 1.346308e-05, 1.336939e-05, 
    1.338967e-05, 1.332224e-05, 1.350414e-05, 1.342652e-05, 1.345628e-05, 
    1.337929e-05, 1.355058e-05, 1.340404e-05, 1.358913e-05, 1.357247e-05, 
    1.352148e-05, 1.342131e-05, 1.339962e-05, 1.337658e-05, 1.339078e-05, 
    1.346053e-05, 1.347212e-05, 1.352272e-05, 1.353682e-05, 1.357609e-05, 
    1.360895e-05, 1.357891e-05, 1.354764e-05, 1.346051e-05, 1.338401e-05, 
    1.330278e-05, 1.328325e-05, 1.319173e-05, 1.326597e-05, 1.314448e-05, 
    1.324737e-05, 1.307168e-05, 1.33958e-05, 1.325051e-05, 1.351919e-05, 
    1.348908e-05, 1.343532e-05, 1.331556e-05, 1.337965e-05, 1.330485e-05, 
    1.347258e-05, 1.356329e-05, 1.358721e-05, 1.363225e-05, 1.358619e-05, 
    1.358991e-05, 1.354637e-05, 1.35603e-05, 1.345766e-05, 1.351239e-05, 
    1.335939e-05, 1.330544e-05, 1.315842e-05, 1.307203e-05, 1.298693e-05, 
    1.29502e-05, 1.293913e-05, 1.293451e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23991, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23998, 18.23999, 18.23999, 18.24, 18.23999, 18.23999, 
    18.23997, 18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 
    18.23991, 18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 
    18.23994, 18.23995, 18.23995, 18.23993, 18.23995, 18.23992, 18.23994, 
    18.23991, 18.23992, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 
    18.23988, 18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 
    18.23996, 18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 
    18.23993, 18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 
    18.23992, 18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 
    18.23985, 18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 
    18.23993, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23996, 
    18.23993, 18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 
    18.23992, 18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 
    18.23996, 18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 
    18.23994, 18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23992, 
    18.23991, 18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 
    18.23995, 18.23992, 18.23993, 18.2399, 18.23991, 18.2399, 18.23991, 
    18.23991, 18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 
    18.23994, 18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 
    18.23992, 18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 
    18.23992, 18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 
    18.23993, 18.23994, 18.23994, 18.23994, 18.23994, 18.23992, 18.23991, 
    18.2399, 18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 
    18.23991, 18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 
    18.2399, 18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 
    18.23994, 18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 
    18.23986, 18.23985, 18.23984, 18.23984, 18.23983 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  6.210302e-05, 6.210287e-05, 6.21029e-05, 6.210276e-05, 6.210284e-05, 
    6.210276e-05, 6.210299e-05, 6.210286e-05, 6.210294e-05, 6.2103e-05, 
    6.210252e-05, 6.210276e-05, 6.210227e-05, 6.210242e-05, 6.210204e-05, 
    6.21023e-05, 6.210199e-05, 6.210204e-05, 6.210187e-05, 6.210192e-05, 
    6.21017e-05, 6.210185e-05, 6.210158e-05, 6.210173e-05, 6.210171e-05, 
    6.210186e-05, 6.210271e-05, 6.210255e-05, 6.210272e-05, 6.21027e-05, 
    6.210271e-05, 6.210284e-05, 6.21029e-05, 6.210303e-05, 6.210301e-05, 
    6.210291e-05, 6.210269e-05, 6.210276e-05, 6.210258e-05, 6.210258e-05, 
    6.210237e-05, 6.210247e-05, 6.210211e-05, 6.210221e-05, 6.210192e-05, 
    6.210199e-05, 6.210192e-05, 6.210194e-05, 6.210192e-05, 6.210203e-05, 
    6.210199e-05, 6.210208e-05, 6.210244e-05, 6.210234e-05, 6.210266e-05, 
    6.210285e-05, 6.210298e-05, 6.210308e-05, 6.210306e-05, 6.210304e-05, 
    6.210291e-05, 6.210279e-05, 6.21027e-05, 6.210264e-05, 6.210258e-05, 
    6.21024e-05, 6.210231e-05, 6.210209e-05, 6.210212e-05, 6.210206e-05, 
    6.2102e-05, 6.21019e-05, 6.210191e-05, 6.210187e-05, 6.210207e-05, 
    6.210194e-05, 6.210215e-05, 6.210209e-05, 6.210256e-05, 6.210274e-05, 
    6.210282e-05, 6.210289e-05, 6.210306e-05, 6.210294e-05, 6.210298e-05, 
    6.210288e-05, 6.210281e-05, 6.210284e-05, 6.210264e-05, 6.210272e-05, 
    6.21023e-05, 6.210248e-05, 6.210201e-05, 6.210212e-05, 6.210198e-05, 
    6.210205e-05, 6.210193e-05, 6.210204e-05, 6.210185e-05, 6.21018e-05, 
    6.210183e-05, 6.210172e-05, 6.210204e-05, 6.210192e-05, 6.210284e-05, 
    6.210284e-05, 6.210282e-05, 6.210292e-05, 6.210293e-05, 6.210303e-05, 
    6.210295e-05, 6.21029e-05, 6.210281e-05, 6.210275e-05, 6.210269e-05, 
    6.210258e-05, 6.210244e-05, 6.210225e-05, 6.210211e-05, 6.210202e-05, 
    6.210208e-05, 6.210203e-05, 6.210208e-05, 6.210211e-05, 6.210183e-05, 
    6.210199e-05, 6.210175e-05, 6.210175e-05, 6.210186e-05, 6.210175e-05, 
    6.210284e-05, 6.210287e-05, 6.210298e-05, 6.210289e-05, 6.210305e-05, 
    6.210296e-05, 6.210291e-05, 6.210271e-05, 6.210268e-05, 6.210263e-05, 
    6.210256e-05, 6.210246e-05, 6.210228e-05, 6.210213e-05, 6.210199e-05, 
    6.210201e-05, 6.2102e-05, 6.210197e-05, 6.210205e-05, 6.210196e-05, 
    6.210194e-05, 6.210199e-05, 6.210176e-05, 6.210183e-05, 6.210175e-05, 
    6.21018e-05, 6.210286e-05, 6.21028e-05, 6.210283e-05, 6.210278e-05, 
    6.210282e-05, 6.210265e-05, 6.21026e-05, 6.210236e-05, 6.210246e-05, 
    6.210231e-05, 6.210244e-05, 6.210242e-05, 6.21023e-05, 6.210244e-05, 
    6.210214e-05, 6.210234e-05, 6.210197e-05, 6.210217e-05, 6.210196e-05, 
    6.210199e-05, 6.210194e-05, 6.210188e-05, 6.21018e-05, 6.210167e-05, 
    6.21017e-05, 6.210159e-05, 6.210273e-05, 6.210266e-05, 6.210266e-05, 
    6.210259e-05, 6.210254e-05, 6.210242e-05, 6.210224e-05, 6.210231e-05, 
    6.210218e-05, 6.210216e-05, 6.210235e-05, 6.210223e-05, 6.210261e-05, 
    6.210255e-05, 6.210259e-05, 6.210272e-05, 6.210229e-05, 6.210251e-05, 
    6.210211e-05, 6.210223e-05, 6.210188e-05, 6.210206e-05, 6.210172e-05, 
    6.210158e-05, 6.210144e-05, 6.210129e-05, 6.210262e-05, 6.210266e-05, 
    6.210258e-05, 6.210247e-05, 6.210236e-05, 6.210222e-05, 6.21022e-05, 
    6.210218e-05, 6.210211e-05, 6.210205e-05, 6.210218e-05, 6.210204e-05, 
    6.210254e-05, 6.210228e-05, 6.210268e-05, 6.210256e-05, 6.210247e-05, 
    6.210251e-05, 6.210232e-05, 6.210227e-05, 6.210209e-05, 6.210218e-05, 
    6.210162e-05, 6.210186e-05, 6.210116e-05, 6.210136e-05, 6.210268e-05, 
    6.210262e-05, 6.21024e-05, 6.210251e-05, 6.210221e-05, 6.210214e-05, 
    6.210208e-05, 6.210201e-05, 6.210199e-05, 6.210195e-05, 6.210202e-05, 
    6.210196e-05, 6.210222e-05, 6.21021e-05, 6.210243e-05, 6.210235e-05, 
    6.210239e-05, 6.210242e-05, 6.21023e-05, 6.210217e-05, 6.210217e-05, 
    6.210212e-05, 6.210201e-05, 6.210221e-05, 6.210158e-05, 6.210197e-05, 
    6.210255e-05, 6.210243e-05, 6.210242e-05, 6.210246e-05, 6.210215e-05, 
    6.210226e-05, 6.210196e-05, 6.210204e-05, 6.21019e-05, 6.210197e-05, 
    6.210198e-05, 6.210207e-05, 6.210212e-05, 6.210226e-05, 6.210236e-05, 
    6.210245e-05, 6.210244e-05, 6.210234e-05, 6.210216e-05, 6.210199e-05, 
    6.210203e-05, 6.210191e-05, 6.210223e-05, 6.21021e-05, 6.210215e-05, 
    6.210202e-05, 6.210231e-05, 6.210206e-05, 6.210238e-05, 6.210235e-05, 
    6.210226e-05, 6.210209e-05, 6.210205e-05, 6.210201e-05, 6.210204e-05, 
    6.210216e-05, 6.210218e-05, 6.210226e-05, 6.210229e-05, 6.210236e-05, 
    6.210241e-05, 6.210236e-05, 6.210231e-05, 6.210216e-05, 6.210202e-05, 
    6.210188e-05, 6.210184e-05, 6.210167e-05, 6.21018e-05, 6.210158e-05, 
    6.210178e-05, 6.210143e-05, 6.210204e-05, 6.210178e-05, 6.210226e-05, 
    6.21022e-05, 6.210211e-05, 6.21019e-05, 6.210202e-05, 6.210188e-05, 
    6.210218e-05, 6.210234e-05, 6.210237e-05, 6.210245e-05, 6.210237e-05, 
    6.210238e-05, 6.210231e-05, 6.210233e-05, 6.210215e-05, 6.210225e-05, 
    6.210198e-05, 6.210188e-05, 6.21016e-05, 6.210143e-05, 6.210127e-05, 
    6.210119e-05, 6.210116e-05, 6.210116e-05 ;

 TOTLITC_1m =
  6.210302e-05, 6.210287e-05, 6.21029e-05, 6.210276e-05, 6.210284e-05, 
    6.210276e-05, 6.210299e-05, 6.210286e-05, 6.210294e-05, 6.2103e-05, 
    6.210252e-05, 6.210276e-05, 6.210227e-05, 6.210242e-05, 6.210204e-05, 
    6.21023e-05, 6.210199e-05, 6.210204e-05, 6.210187e-05, 6.210192e-05, 
    6.21017e-05, 6.210185e-05, 6.210158e-05, 6.210173e-05, 6.210171e-05, 
    6.210186e-05, 6.210271e-05, 6.210255e-05, 6.210272e-05, 6.21027e-05, 
    6.210271e-05, 6.210284e-05, 6.21029e-05, 6.210303e-05, 6.210301e-05, 
    6.210291e-05, 6.210269e-05, 6.210276e-05, 6.210258e-05, 6.210258e-05, 
    6.210237e-05, 6.210247e-05, 6.210211e-05, 6.210221e-05, 6.210192e-05, 
    6.210199e-05, 6.210192e-05, 6.210194e-05, 6.210192e-05, 6.210203e-05, 
    6.210199e-05, 6.210208e-05, 6.210244e-05, 6.210234e-05, 6.210266e-05, 
    6.210285e-05, 6.210298e-05, 6.210308e-05, 6.210306e-05, 6.210304e-05, 
    6.210291e-05, 6.210279e-05, 6.21027e-05, 6.210264e-05, 6.210258e-05, 
    6.21024e-05, 6.210231e-05, 6.210209e-05, 6.210212e-05, 6.210206e-05, 
    6.2102e-05, 6.21019e-05, 6.210191e-05, 6.210187e-05, 6.210207e-05, 
    6.210194e-05, 6.210215e-05, 6.210209e-05, 6.210256e-05, 6.210274e-05, 
    6.210282e-05, 6.210289e-05, 6.210306e-05, 6.210294e-05, 6.210298e-05, 
    6.210288e-05, 6.210281e-05, 6.210284e-05, 6.210264e-05, 6.210272e-05, 
    6.21023e-05, 6.210248e-05, 6.210201e-05, 6.210212e-05, 6.210198e-05, 
    6.210205e-05, 6.210193e-05, 6.210204e-05, 6.210185e-05, 6.21018e-05, 
    6.210183e-05, 6.210172e-05, 6.210204e-05, 6.210192e-05, 6.210284e-05, 
    6.210284e-05, 6.210282e-05, 6.210292e-05, 6.210293e-05, 6.210303e-05, 
    6.210295e-05, 6.21029e-05, 6.210281e-05, 6.210275e-05, 6.210269e-05, 
    6.210258e-05, 6.210244e-05, 6.210225e-05, 6.210211e-05, 6.210202e-05, 
    6.210208e-05, 6.210203e-05, 6.210208e-05, 6.210211e-05, 6.210183e-05, 
    6.210199e-05, 6.210175e-05, 6.210175e-05, 6.210186e-05, 6.210175e-05, 
    6.210284e-05, 6.210287e-05, 6.210298e-05, 6.210289e-05, 6.210305e-05, 
    6.210296e-05, 6.210291e-05, 6.210271e-05, 6.210268e-05, 6.210263e-05, 
    6.210256e-05, 6.210246e-05, 6.210228e-05, 6.210213e-05, 6.210199e-05, 
    6.210201e-05, 6.2102e-05, 6.210197e-05, 6.210205e-05, 6.210196e-05, 
    6.210194e-05, 6.210199e-05, 6.210176e-05, 6.210183e-05, 6.210175e-05, 
    6.21018e-05, 6.210286e-05, 6.21028e-05, 6.210283e-05, 6.210278e-05, 
    6.210282e-05, 6.210265e-05, 6.21026e-05, 6.210236e-05, 6.210246e-05, 
    6.210231e-05, 6.210244e-05, 6.210242e-05, 6.21023e-05, 6.210244e-05, 
    6.210214e-05, 6.210234e-05, 6.210197e-05, 6.210217e-05, 6.210196e-05, 
    6.210199e-05, 6.210194e-05, 6.210188e-05, 6.21018e-05, 6.210167e-05, 
    6.21017e-05, 6.210159e-05, 6.210273e-05, 6.210266e-05, 6.210266e-05, 
    6.210259e-05, 6.210254e-05, 6.210242e-05, 6.210224e-05, 6.210231e-05, 
    6.210218e-05, 6.210216e-05, 6.210235e-05, 6.210223e-05, 6.210261e-05, 
    6.210255e-05, 6.210259e-05, 6.210272e-05, 6.210229e-05, 6.210251e-05, 
    6.210211e-05, 6.210223e-05, 6.210188e-05, 6.210206e-05, 6.210172e-05, 
    6.210158e-05, 6.210144e-05, 6.210129e-05, 6.210262e-05, 6.210266e-05, 
    6.210258e-05, 6.210247e-05, 6.210236e-05, 6.210222e-05, 6.21022e-05, 
    6.210218e-05, 6.210211e-05, 6.210205e-05, 6.210218e-05, 6.210204e-05, 
    6.210254e-05, 6.210228e-05, 6.210268e-05, 6.210256e-05, 6.210247e-05, 
    6.210251e-05, 6.210232e-05, 6.210227e-05, 6.210209e-05, 6.210218e-05, 
    6.210162e-05, 6.210186e-05, 6.210116e-05, 6.210136e-05, 6.210268e-05, 
    6.210262e-05, 6.21024e-05, 6.210251e-05, 6.210221e-05, 6.210214e-05, 
    6.210208e-05, 6.210201e-05, 6.210199e-05, 6.210195e-05, 6.210202e-05, 
    6.210196e-05, 6.210222e-05, 6.21021e-05, 6.210243e-05, 6.210235e-05, 
    6.210239e-05, 6.210242e-05, 6.21023e-05, 6.210217e-05, 6.210217e-05, 
    6.210212e-05, 6.210201e-05, 6.210221e-05, 6.210158e-05, 6.210197e-05, 
    6.210255e-05, 6.210243e-05, 6.210242e-05, 6.210246e-05, 6.210215e-05, 
    6.210226e-05, 6.210196e-05, 6.210204e-05, 6.21019e-05, 6.210197e-05, 
    6.210198e-05, 6.210207e-05, 6.210212e-05, 6.210226e-05, 6.210236e-05, 
    6.210245e-05, 6.210244e-05, 6.210234e-05, 6.210216e-05, 6.210199e-05, 
    6.210203e-05, 6.210191e-05, 6.210223e-05, 6.21021e-05, 6.210215e-05, 
    6.210202e-05, 6.210231e-05, 6.210206e-05, 6.210238e-05, 6.210235e-05, 
    6.210226e-05, 6.210209e-05, 6.210205e-05, 6.210201e-05, 6.210204e-05, 
    6.210216e-05, 6.210218e-05, 6.210226e-05, 6.210229e-05, 6.210236e-05, 
    6.210241e-05, 6.210236e-05, 6.210231e-05, 6.210216e-05, 6.210202e-05, 
    6.210188e-05, 6.210184e-05, 6.210167e-05, 6.21018e-05, 6.210158e-05, 
    6.210178e-05, 6.210143e-05, 6.210204e-05, 6.210178e-05, 6.210226e-05, 
    6.21022e-05, 6.210211e-05, 6.21019e-05, 6.210202e-05, 6.210188e-05, 
    6.210218e-05, 6.210234e-05, 6.210237e-05, 6.210245e-05, 6.210237e-05, 
    6.210238e-05, 6.210231e-05, 6.210233e-05, 6.210215e-05, 6.210225e-05, 
    6.210198e-05, 6.210188e-05, 6.21016e-05, 6.210143e-05, 6.210127e-05, 
    6.210119e-05, 6.210116e-05, 6.210116e-05 ;

 TOTLITN =
  1.429816e-06, 1.429811e-06, 1.429812e-06, 1.429808e-06, 1.42981e-06, 
    1.429808e-06, 1.429815e-06, 1.429811e-06, 1.429813e-06, 1.429815e-06, 
    1.429802e-06, 1.429808e-06, 1.429795e-06, 1.429799e-06, 1.429788e-06, 
    1.429795e-06, 1.429787e-06, 1.429788e-06, 1.429783e-06, 1.429785e-06, 
    1.429778e-06, 1.429783e-06, 1.429775e-06, 1.429779e-06, 1.429779e-06, 
    1.429783e-06, 1.429807e-06, 1.429802e-06, 1.429807e-06, 1.429807e-06, 
    1.429807e-06, 1.42981e-06, 1.429812e-06, 1.429816e-06, 1.429815e-06, 
    1.429813e-06, 1.429806e-06, 1.429808e-06, 1.429803e-06, 1.429803e-06, 
    1.429797e-06, 1.4298e-06, 1.42979e-06, 1.429793e-06, 1.429785e-06, 
    1.429787e-06, 1.429785e-06, 1.429785e-06, 1.429785e-06, 1.429788e-06, 
    1.429786e-06, 1.429789e-06, 1.429799e-06, 1.429796e-06, 1.429805e-06, 
    1.429811e-06, 1.429815e-06, 1.429817e-06, 1.429817e-06, 1.429816e-06, 
    1.429813e-06, 1.429809e-06, 1.429807e-06, 1.429805e-06, 1.429803e-06, 
    1.429798e-06, 1.429795e-06, 1.429789e-06, 1.42979e-06, 1.429789e-06, 
    1.429787e-06, 1.429784e-06, 1.429784e-06, 1.429783e-06, 1.429789e-06, 
    1.429785e-06, 1.429791e-06, 1.429789e-06, 1.429803e-06, 1.429808e-06, 
    1.42981e-06, 1.429812e-06, 1.429817e-06, 1.429813e-06, 1.429815e-06, 
    1.429812e-06, 1.42981e-06, 1.429811e-06, 1.429805e-06, 1.429807e-06, 
    1.429795e-06, 1.4298e-06, 1.429787e-06, 1.42979e-06, 1.429786e-06, 
    1.429788e-06, 1.429785e-06, 1.429788e-06, 1.429783e-06, 1.429781e-06, 
    1.429782e-06, 1.429779e-06, 1.429788e-06, 1.429785e-06, 1.429811e-06, 
    1.42981e-06, 1.42981e-06, 1.429813e-06, 1.429813e-06, 1.429816e-06, 
    1.429813e-06, 1.429812e-06, 1.42981e-06, 1.429808e-06, 1.429806e-06, 
    1.429803e-06, 1.429799e-06, 1.429794e-06, 1.42979e-06, 1.429788e-06, 
    1.429789e-06, 1.429788e-06, 1.429789e-06, 1.42979e-06, 1.429782e-06, 
    1.429786e-06, 1.42978e-06, 1.42978e-06, 1.429783e-06, 1.42978e-06, 
    1.42981e-06, 1.429811e-06, 1.429814e-06, 1.429812e-06, 1.429816e-06, 
    1.429814e-06, 1.429812e-06, 1.429807e-06, 1.429806e-06, 1.429805e-06, 
    1.429803e-06, 1.4298e-06, 1.429795e-06, 1.429791e-06, 1.429787e-06, 
    1.429787e-06, 1.429787e-06, 1.429786e-06, 1.429788e-06, 1.429786e-06, 
    1.429785e-06, 1.429786e-06, 1.42978e-06, 1.429782e-06, 1.42978e-06, 
    1.429781e-06, 1.429811e-06, 1.429809e-06, 1.42981e-06, 1.429809e-06, 
    1.42981e-06, 1.429805e-06, 1.429804e-06, 1.429797e-06, 1.4298e-06, 
    1.429795e-06, 1.429799e-06, 1.429799e-06, 1.429795e-06, 1.429799e-06, 
    1.429791e-06, 1.429796e-06, 1.429786e-06, 1.429792e-06, 1.429786e-06, 
    1.429787e-06, 1.429785e-06, 1.429783e-06, 1.429781e-06, 1.429778e-06, 
    1.429779e-06, 1.429775e-06, 1.429807e-06, 1.429805e-06, 1.429805e-06, 
    1.429804e-06, 1.429802e-06, 1.429799e-06, 1.429794e-06, 1.429796e-06, 
    1.429792e-06, 1.429791e-06, 1.429797e-06, 1.429793e-06, 1.429804e-06, 
    1.429802e-06, 1.429803e-06, 1.429807e-06, 1.429795e-06, 1.429801e-06, 
    1.42979e-06, 1.429793e-06, 1.429784e-06, 1.429788e-06, 1.429779e-06, 
    1.429775e-06, 1.429771e-06, 1.429767e-06, 1.429804e-06, 1.429806e-06, 
    1.429803e-06, 1.4298e-06, 1.429797e-06, 1.429793e-06, 1.429793e-06, 
    1.429792e-06, 1.42979e-06, 1.429788e-06, 1.429792e-06, 1.429788e-06, 
    1.429802e-06, 1.429795e-06, 1.429806e-06, 1.429803e-06, 1.4298e-06, 
    1.429801e-06, 1.429796e-06, 1.429795e-06, 1.429789e-06, 1.429792e-06, 
    1.429776e-06, 1.429783e-06, 1.429763e-06, 1.429769e-06, 1.429806e-06, 
    1.429804e-06, 1.429798e-06, 1.429801e-06, 1.429793e-06, 1.429791e-06, 
    1.429789e-06, 1.429787e-06, 1.429787e-06, 1.429785e-06, 1.429788e-06, 
    1.429786e-06, 1.429793e-06, 1.42979e-06, 1.429799e-06, 1.429797e-06, 
    1.429798e-06, 1.429799e-06, 1.429795e-06, 1.429792e-06, 1.429792e-06, 
    1.42979e-06, 1.429787e-06, 1.429793e-06, 1.429775e-06, 1.429786e-06, 
    1.429802e-06, 1.429799e-06, 1.429799e-06, 1.4298e-06, 1.429791e-06, 
    1.429794e-06, 1.429786e-06, 1.429788e-06, 1.429784e-06, 1.429786e-06, 
    1.429786e-06, 1.429789e-06, 1.42979e-06, 1.429794e-06, 1.429797e-06, 
    1.4298e-06, 1.429799e-06, 1.429796e-06, 1.429791e-06, 1.429787e-06, 
    1.429788e-06, 1.429784e-06, 1.429793e-06, 1.42979e-06, 1.429791e-06, 
    1.429787e-06, 1.429796e-06, 1.429789e-06, 1.429798e-06, 1.429797e-06, 
    1.429794e-06, 1.429789e-06, 1.429788e-06, 1.429787e-06, 1.429788e-06, 
    1.429791e-06, 1.429792e-06, 1.429794e-06, 1.429795e-06, 1.429797e-06, 
    1.429798e-06, 1.429797e-06, 1.429795e-06, 1.429791e-06, 1.429788e-06, 
    1.429783e-06, 1.429782e-06, 1.429778e-06, 1.429781e-06, 1.429775e-06, 
    1.42978e-06, 1.429771e-06, 1.429788e-06, 1.429781e-06, 1.429794e-06, 
    1.429793e-06, 1.42979e-06, 1.429784e-06, 1.429787e-06, 1.429783e-06, 
    1.429792e-06, 1.429796e-06, 1.429797e-06, 1.4298e-06, 1.429797e-06, 
    1.429798e-06, 1.429795e-06, 1.429796e-06, 1.429791e-06, 1.429794e-06, 
    1.429786e-06, 1.429784e-06, 1.429776e-06, 1.429771e-06, 1.429766e-06, 
    1.429764e-06, 1.429763e-06, 1.429763e-06 ;

 TOTLITN_1m =
  1.429816e-06, 1.429811e-06, 1.429812e-06, 1.429808e-06, 1.42981e-06, 
    1.429808e-06, 1.429815e-06, 1.429811e-06, 1.429813e-06, 1.429815e-06, 
    1.429802e-06, 1.429808e-06, 1.429795e-06, 1.429799e-06, 1.429788e-06, 
    1.429795e-06, 1.429787e-06, 1.429788e-06, 1.429783e-06, 1.429785e-06, 
    1.429778e-06, 1.429783e-06, 1.429775e-06, 1.429779e-06, 1.429779e-06, 
    1.429783e-06, 1.429807e-06, 1.429802e-06, 1.429807e-06, 1.429807e-06, 
    1.429807e-06, 1.42981e-06, 1.429812e-06, 1.429816e-06, 1.429815e-06, 
    1.429813e-06, 1.429806e-06, 1.429808e-06, 1.429803e-06, 1.429803e-06, 
    1.429797e-06, 1.4298e-06, 1.42979e-06, 1.429793e-06, 1.429785e-06, 
    1.429787e-06, 1.429785e-06, 1.429785e-06, 1.429785e-06, 1.429788e-06, 
    1.429786e-06, 1.429789e-06, 1.429799e-06, 1.429796e-06, 1.429805e-06, 
    1.429811e-06, 1.429815e-06, 1.429817e-06, 1.429817e-06, 1.429816e-06, 
    1.429813e-06, 1.429809e-06, 1.429807e-06, 1.429805e-06, 1.429803e-06, 
    1.429798e-06, 1.429795e-06, 1.429789e-06, 1.42979e-06, 1.429789e-06, 
    1.429787e-06, 1.429784e-06, 1.429784e-06, 1.429783e-06, 1.429789e-06, 
    1.429785e-06, 1.429791e-06, 1.429789e-06, 1.429803e-06, 1.429808e-06, 
    1.42981e-06, 1.429812e-06, 1.429817e-06, 1.429813e-06, 1.429815e-06, 
    1.429812e-06, 1.42981e-06, 1.429811e-06, 1.429805e-06, 1.429807e-06, 
    1.429795e-06, 1.4298e-06, 1.429787e-06, 1.42979e-06, 1.429786e-06, 
    1.429788e-06, 1.429785e-06, 1.429788e-06, 1.429783e-06, 1.429781e-06, 
    1.429782e-06, 1.429779e-06, 1.429788e-06, 1.429785e-06, 1.429811e-06, 
    1.42981e-06, 1.42981e-06, 1.429813e-06, 1.429813e-06, 1.429816e-06, 
    1.429813e-06, 1.429812e-06, 1.42981e-06, 1.429808e-06, 1.429806e-06, 
    1.429803e-06, 1.429799e-06, 1.429794e-06, 1.42979e-06, 1.429788e-06, 
    1.429789e-06, 1.429788e-06, 1.429789e-06, 1.42979e-06, 1.429782e-06, 
    1.429786e-06, 1.42978e-06, 1.42978e-06, 1.429783e-06, 1.42978e-06, 
    1.42981e-06, 1.429811e-06, 1.429814e-06, 1.429812e-06, 1.429816e-06, 
    1.429814e-06, 1.429812e-06, 1.429807e-06, 1.429806e-06, 1.429805e-06, 
    1.429803e-06, 1.4298e-06, 1.429795e-06, 1.429791e-06, 1.429787e-06, 
    1.429787e-06, 1.429787e-06, 1.429786e-06, 1.429788e-06, 1.429786e-06, 
    1.429785e-06, 1.429786e-06, 1.42978e-06, 1.429782e-06, 1.42978e-06, 
    1.429781e-06, 1.429811e-06, 1.429809e-06, 1.42981e-06, 1.429809e-06, 
    1.42981e-06, 1.429805e-06, 1.429804e-06, 1.429797e-06, 1.4298e-06, 
    1.429795e-06, 1.429799e-06, 1.429799e-06, 1.429795e-06, 1.429799e-06, 
    1.429791e-06, 1.429796e-06, 1.429786e-06, 1.429792e-06, 1.429786e-06, 
    1.429787e-06, 1.429785e-06, 1.429783e-06, 1.429781e-06, 1.429778e-06, 
    1.429779e-06, 1.429775e-06, 1.429807e-06, 1.429805e-06, 1.429805e-06, 
    1.429804e-06, 1.429802e-06, 1.429799e-06, 1.429794e-06, 1.429796e-06, 
    1.429792e-06, 1.429791e-06, 1.429797e-06, 1.429793e-06, 1.429804e-06, 
    1.429802e-06, 1.429803e-06, 1.429807e-06, 1.429795e-06, 1.429801e-06, 
    1.42979e-06, 1.429793e-06, 1.429784e-06, 1.429788e-06, 1.429779e-06, 
    1.429775e-06, 1.429771e-06, 1.429767e-06, 1.429804e-06, 1.429806e-06, 
    1.429803e-06, 1.4298e-06, 1.429797e-06, 1.429793e-06, 1.429793e-06, 
    1.429792e-06, 1.42979e-06, 1.429788e-06, 1.429792e-06, 1.429788e-06, 
    1.429802e-06, 1.429795e-06, 1.429806e-06, 1.429803e-06, 1.4298e-06, 
    1.429801e-06, 1.429796e-06, 1.429795e-06, 1.429789e-06, 1.429792e-06, 
    1.429776e-06, 1.429783e-06, 1.429763e-06, 1.429769e-06, 1.429806e-06, 
    1.429804e-06, 1.429798e-06, 1.429801e-06, 1.429793e-06, 1.429791e-06, 
    1.429789e-06, 1.429787e-06, 1.429787e-06, 1.429785e-06, 1.429788e-06, 
    1.429786e-06, 1.429793e-06, 1.42979e-06, 1.429799e-06, 1.429797e-06, 
    1.429798e-06, 1.429799e-06, 1.429795e-06, 1.429792e-06, 1.429792e-06, 
    1.42979e-06, 1.429787e-06, 1.429793e-06, 1.429775e-06, 1.429786e-06, 
    1.429802e-06, 1.429799e-06, 1.429799e-06, 1.4298e-06, 1.429791e-06, 
    1.429794e-06, 1.429786e-06, 1.429788e-06, 1.429784e-06, 1.429786e-06, 
    1.429786e-06, 1.429789e-06, 1.42979e-06, 1.429794e-06, 1.429797e-06, 
    1.4298e-06, 1.429799e-06, 1.429796e-06, 1.429791e-06, 1.429787e-06, 
    1.429788e-06, 1.429784e-06, 1.429793e-06, 1.42979e-06, 1.429791e-06, 
    1.429787e-06, 1.429796e-06, 1.429789e-06, 1.429798e-06, 1.429797e-06, 
    1.429794e-06, 1.429789e-06, 1.429788e-06, 1.429787e-06, 1.429788e-06, 
    1.429791e-06, 1.429792e-06, 1.429794e-06, 1.429795e-06, 1.429797e-06, 
    1.429798e-06, 1.429797e-06, 1.429795e-06, 1.429791e-06, 1.429788e-06, 
    1.429783e-06, 1.429782e-06, 1.429778e-06, 1.429781e-06, 1.429775e-06, 
    1.42978e-06, 1.429771e-06, 1.429788e-06, 1.429781e-06, 1.429794e-06, 
    1.429793e-06, 1.42979e-06, 1.429784e-06, 1.429787e-06, 1.429783e-06, 
    1.429792e-06, 1.429796e-06, 1.429797e-06, 1.4298e-06, 1.429797e-06, 
    1.429798e-06, 1.429795e-06, 1.429796e-06, 1.429791e-06, 1.429794e-06, 
    1.429786e-06, 1.429784e-06, 1.429776e-06, 1.429771e-06, 1.429766e-06, 
    1.429764e-06, 1.429763e-06, 1.429763e-06 ;

 TOTPFTC =
  0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174 ;

 TOTPFTN =
  0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.34459, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34452, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34455, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34452, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.3445, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.34449, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34456, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34455, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34455, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMC_1m =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.34459, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34452, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34455, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34452, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.3445, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.34449, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34456, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34455, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34455, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMN =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773748, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773758, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773745, 1.773744, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773754, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773736, 1.773739, 1.773755, 1.773754, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773752, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773751, 1.773751, 1.77375, 1.773748, 1.773747, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773751, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTSOMN_1m =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773748, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773758, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773745, 1.773744, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773754, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773736, 1.773739, 1.773755, 1.773754, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773752, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773751, 1.773751, 1.77375, 1.773748, 1.773747, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773751, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTVEGC =
  0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174 ;

 TOTVEGN =
  0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255 ;

 TREFMNAV =
  243.0873, 243.0906, 243.0899, 243.0925, 243.0911, 243.0928, 243.088, 
    243.0907, 243.089, 243.0876, 243.0974, 243.0926, 243.1026, 243.0995, 
    243.1073, 243.1021, 243.1083, 243.1072, 243.1107, 243.1097, 243.1142, 
    243.1112, 243.1166, 243.1135, 243.114, 243.1111, 243.0937, 243.0968, 
    243.0935, 243.0939, 243.0937, 243.0911, 243.0898, 243.0871, 243.0876, 
    243.0896, 243.0941, 243.0926, 243.0965, 243.0964, 243.1007, 243.0988, 
    243.1059, 243.1039, 243.1098, 243.1083, 243.1097, 243.1093, 243.1097, 
    243.1075, 243.1085, 243.1066, 243.0991, 243.1013, 243.0947, 243.0907, 
    243.0881, 243.0862, 243.0865, 243.087, 243.0896, 243.0921, 243.0939, 
    243.0952, 243.0964, 243.0999, 243.1019, 243.1063, 243.1056, 243.1069, 
    243.1082, 243.1103, 243.1099, 243.1108, 243.1069, 243.1095, 243.1051, 
    243.1063, 243.0965, 243.093, 243.0914, 243.0901, 243.0867, 243.089, 
    243.0881, 243.0903, 243.0917, 243.091, 243.0952, 243.0936, 243.1021, 
    243.0984, 243.108, 243.1057, 243.1086, 243.1071, 243.1096, 243.1074, 
    243.1112, 243.112, 243.1114, 243.1136, 243.1072, 243.1097, 243.091, 
    243.0911, 243.0916, 243.0893, 243.0892, 243.0871, 243.0889, 243.0897, 
    243.0918, 243.0929, 243.0941, 243.0965, 243.0993, 243.1031, 243.1059, 
    243.1077, 243.1066, 243.1076, 243.1065, 243.106, 243.1117, 243.1085, 
    243.1133, 243.1131, 243.1108, 243.1131, 243.0912, 243.0905, 243.0883, 
    243.09, 243.0869, 243.0886, 243.0896, 243.0936, 243.0945, 243.0952, 
    243.0968, 243.0988, 243.1024, 243.1054, 243.1082, 243.108, 243.1081, 
    243.1087, 243.1072, 243.109, 243.1092, 243.1085, 243.113, 243.1117, 
    243.1131, 243.1122, 243.0907, 243.0918, 243.0912, 243.0923, 243.0915, 
    243.0949, 243.0959, 243.1007, 243.0988, 243.1019, 243.0991, 243.0996, 
    243.1019, 243.0993, 243.1052, 243.1011, 243.1087, 243.1046, 243.109, 
    243.1082, 243.1095, 243.1106, 243.1121, 243.1147, 243.1141, 243.1163, 
    243.0934, 243.0948, 243.0947, 243.0961, 243.0972, 243.0995, 243.1032, 
    243.1019, 243.1044, 243.1049, 243.1011, 243.1034, 243.0957, 243.0969, 
    243.0962, 243.0935, 243.1021, 243.0977, 243.1059, 243.1035, 243.1105, 
    243.107, 243.1138, 243.1166, 243.1194, 243.1224, 243.0956, 243.0946, 
    243.0963, 243.0986, 243.1008, 243.1037, 243.104, 243.1045, 243.1059, 
    243.1071, 243.1046, 243.1074, 243.0971, 243.1025, 243.0943, 243.0967, 
    243.0985, 243.0977, 243.1017, 243.1026, 243.1064, 243.1045, 243.1159, 
    243.1108, 243.1248, 243.1209, 243.0943, 243.0956, 243.0999, 243.0979, 
    243.1039, 243.1053, 243.1065, 243.108, 243.1082, 243.1091, 243.1077, 
    243.1091, 243.1037, 243.1061, 243.0995, 243.1011, 243.1004, 243.0995, 
    243.1021, 243.1047, 243.1048, 243.1056, 243.1078, 243.1039, 243.1164, 
    243.1086, 243.097, 243.0993, 243.0997, 243.0988, 243.1052, 243.1029, 
    243.1091, 243.1074, 243.1102, 243.1088, 243.1086, 243.1068, 243.1057, 
    243.103, 243.1007, 243.099, 243.0994, 243.1013, 243.1048, 243.1082, 
    243.1075, 243.11, 243.1034, 243.1061, 243.1051, 243.1079, 243.1018, 
    243.1068, 243.1005, 243.1011, 243.1028, 243.1063, 243.1071, 243.1079, 
    243.1075, 243.1049, 243.1045, 243.1028, 243.1023, 243.101, 243.0998, 
    243.1009, 243.1019, 243.105, 243.1077, 243.1106, 243.1114, 243.1147, 
    243.1119, 243.1164, 243.1125, 243.1194, 243.1072, 243.1125, 243.1029, 
    243.104, 243.1058, 243.1101, 243.1078, 243.1105, 243.1045, 243.1013, 
    243.1006, 243.099, 243.1006, 243.1005, 243.102, 243.1015, 243.1051, 
    243.1031, 243.1086, 243.1105, 243.1161, 243.1194, 243.1229, 243.1244, 
    243.1249, 243.1251 ;

 TREFMNAV_R =
  243.0873, 243.0906, 243.0899, 243.0925, 243.0911, 243.0928, 243.088, 
    243.0907, 243.089, 243.0876, 243.0974, 243.0926, 243.1026, 243.0995, 
    243.1073, 243.1021, 243.1083, 243.1072, 243.1107, 243.1097, 243.1142, 
    243.1112, 243.1166, 243.1135, 243.114, 243.1111, 243.0937, 243.0968, 
    243.0935, 243.0939, 243.0937, 243.0911, 243.0898, 243.0871, 243.0876, 
    243.0896, 243.0941, 243.0926, 243.0965, 243.0964, 243.1007, 243.0988, 
    243.1059, 243.1039, 243.1098, 243.1083, 243.1097, 243.1093, 243.1097, 
    243.1075, 243.1085, 243.1066, 243.0991, 243.1013, 243.0947, 243.0907, 
    243.0881, 243.0862, 243.0865, 243.087, 243.0896, 243.0921, 243.0939, 
    243.0952, 243.0964, 243.0999, 243.1019, 243.1063, 243.1056, 243.1069, 
    243.1082, 243.1103, 243.1099, 243.1108, 243.1069, 243.1095, 243.1051, 
    243.1063, 243.0965, 243.093, 243.0914, 243.0901, 243.0867, 243.089, 
    243.0881, 243.0903, 243.0917, 243.091, 243.0952, 243.0936, 243.1021, 
    243.0984, 243.108, 243.1057, 243.1086, 243.1071, 243.1096, 243.1074, 
    243.1112, 243.112, 243.1114, 243.1136, 243.1072, 243.1097, 243.091, 
    243.0911, 243.0916, 243.0893, 243.0892, 243.0871, 243.0889, 243.0897, 
    243.0918, 243.0929, 243.0941, 243.0965, 243.0993, 243.1031, 243.1059, 
    243.1077, 243.1066, 243.1076, 243.1065, 243.106, 243.1117, 243.1085, 
    243.1133, 243.1131, 243.1108, 243.1131, 243.0912, 243.0905, 243.0883, 
    243.09, 243.0869, 243.0886, 243.0896, 243.0936, 243.0945, 243.0952, 
    243.0968, 243.0988, 243.1024, 243.1054, 243.1082, 243.108, 243.1081, 
    243.1087, 243.1072, 243.109, 243.1092, 243.1085, 243.113, 243.1117, 
    243.1131, 243.1122, 243.0907, 243.0918, 243.0912, 243.0923, 243.0915, 
    243.0949, 243.0959, 243.1007, 243.0988, 243.1019, 243.0991, 243.0996, 
    243.1019, 243.0993, 243.1052, 243.1011, 243.1087, 243.1046, 243.109, 
    243.1082, 243.1095, 243.1106, 243.1121, 243.1147, 243.1141, 243.1163, 
    243.0934, 243.0948, 243.0947, 243.0961, 243.0972, 243.0995, 243.1032, 
    243.1019, 243.1044, 243.1049, 243.1011, 243.1034, 243.0957, 243.0969, 
    243.0962, 243.0935, 243.1021, 243.0977, 243.1059, 243.1035, 243.1105, 
    243.107, 243.1138, 243.1166, 243.1194, 243.1224, 243.0956, 243.0946, 
    243.0963, 243.0986, 243.1008, 243.1037, 243.104, 243.1045, 243.1059, 
    243.1071, 243.1046, 243.1074, 243.0971, 243.1025, 243.0943, 243.0967, 
    243.0985, 243.0977, 243.1017, 243.1026, 243.1064, 243.1045, 243.1159, 
    243.1108, 243.1248, 243.1209, 243.0943, 243.0956, 243.0999, 243.0979, 
    243.1039, 243.1053, 243.1065, 243.108, 243.1082, 243.1091, 243.1077, 
    243.1091, 243.1037, 243.1061, 243.0995, 243.1011, 243.1004, 243.0995, 
    243.1021, 243.1047, 243.1048, 243.1056, 243.1078, 243.1039, 243.1164, 
    243.1086, 243.097, 243.0993, 243.0997, 243.0988, 243.1052, 243.1029, 
    243.1091, 243.1074, 243.1102, 243.1088, 243.1086, 243.1068, 243.1057, 
    243.103, 243.1007, 243.099, 243.0994, 243.1013, 243.1048, 243.1082, 
    243.1075, 243.11, 243.1034, 243.1061, 243.1051, 243.1079, 243.1018, 
    243.1068, 243.1005, 243.1011, 243.1028, 243.1063, 243.1071, 243.1079, 
    243.1075, 243.1049, 243.1045, 243.1028, 243.1023, 243.101, 243.0998, 
    243.1009, 243.1019, 243.105, 243.1077, 243.1106, 243.1114, 243.1147, 
    243.1119, 243.1164, 243.1125, 243.1194, 243.1072, 243.1125, 243.1029, 
    243.104, 243.1058, 243.1101, 243.1078, 243.1105, 243.1045, 243.1013, 
    243.1006, 243.099, 243.1006, 243.1005, 243.102, 243.1015, 243.1051, 
    243.1031, 243.1086, 243.1105, 243.1161, 243.1194, 243.1229, 243.1244, 
    243.1249, 243.1251 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  270.7703, 270.7681, 270.7685, 270.7668, 270.7678, 270.7667, 270.7698, 
    270.7681, 270.7692, 270.7701, 270.7636, 270.7668, 270.7602, 270.7622, 
    270.757, 270.7605, 270.7563, 270.7571, 270.7547, 270.7554, 270.7524, 
    270.7544, 270.7508, 270.7528, 270.7525, 270.7545, 270.7661, 270.764, 
    270.7662, 270.7659, 270.7661, 270.7678, 270.7686, 270.7704, 270.7701, 
    270.7688, 270.7658, 270.7668, 270.7642, 270.7643, 270.7614, 270.7627, 
    270.7579, 270.7593, 270.7553, 270.7563, 270.7554, 270.7557, 270.7554, 
    270.7569, 270.7562, 270.7575, 270.7625, 270.761, 270.7654, 270.7681, 
    270.7697, 270.771, 270.7708, 270.7705, 270.7688, 270.7671, 270.7659, 
    270.7651, 270.7643, 270.7619, 270.7606, 270.7577, 270.7582, 270.7573, 
    270.7564, 270.755, 270.7552, 270.7546, 270.7573, 270.7556, 270.7585, 
    270.7577, 270.7642, 270.7665, 270.7676, 270.7685, 270.7707, 270.7691, 
    270.7697, 270.7683, 270.7674, 270.7678, 270.7651, 270.7661, 270.7605, 
    270.7629, 270.7566, 270.7581, 270.7562, 270.7571, 270.7555, 270.757, 
    270.7544, 270.7539, 270.7542, 270.7527, 270.757, 270.7554, 270.7679, 
    270.7678, 270.7674, 270.769, 270.769, 270.7704, 270.7692, 270.7687, 
    270.7673, 270.7666, 270.7658, 270.7642, 270.7624, 270.7598, 270.758, 
    270.7567, 270.7575, 270.7568, 270.7576, 270.7579, 270.7541, 270.7562, 
    270.753, 270.7531, 270.7546, 270.7531, 270.7677, 270.7681, 270.7696, 
    270.7685, 270.7705, 270.7694, 270.7687, 270.7661, 270.7655, 270.765, 
    270.764, 270.7627, 270.7603, 270.7583, 270.7564, 270.7565, 270.7565, 
    270.7561, 270.7571, 270.7559, 270.7557, 270.7562, 270.7532, 270.754, 
    270.7531, 270.7537, 270.768, 270.7673, 270.7677, 270.767, 270.7675, 
    270.7653, 270.7646, 270.7614, 270.7627, 270.7606, 270.7625, 270.7621, 
    270.7606, 270.7624, 270.7584, 270.7611, 270.756, 270.7588, 270.7559, 
    270.7564, 270.7555, 270.7548, 270.7538, 270.752, 270.7524, 270.7509, 
    270.7662, 270.7654, 270.7654, 270.7644, 270.7637, 270.7622, 270.7597, 
    270.7607, 270.7589, 270.7586, 270.7612, 270.7596, 270.7647, 270.7639, 
    270.7644, 270.7662, 270.7605, 270.7634, 270.7579, 270.7596, 270.7549, 
    270.7572, 270.7527, 270.7508, 270.7489, 270.7468, 270.7648, 270.7654, 
    270.7643, 270.7628, 270.7614, 270.7595, 270.7592, 270.7589, 270.758, 
    270.7572, 270.7588, 270.757, 270.7638, 270.7602, 270.7657, 270.7641, 
    270.7629, 270.7634, 270.7607, 270.7601, 270.7576, 270.7589, 270.7513, 
    270.7546, 270.7451, 270.7478, 270.7657, 270.7648, 270.7619, 270.7633, 
    270.7593, 270.7583, 270.7575, 270.7565, 270.7564, 270.7558, 270.7568, 
    270.7558, 270.7594, 270.7578, 270.7622, 270.7612, 270.7617, 270.7622, 
    270.7605, 270.7588, 270.7587, 270.7581, 270.7567, 270.7593, 270.7509, 
    270.7562, 270.7639, 270.7623, 270.7621, 270.7627, 270.7584, 270.76, 
    270.7558, 270.7569, 270.7551, 270.756, 270.7562, 270.7573, 270.7581, 
    270.7599, 270.7614, 270.7626, 270.7623, 270.761, 270.7587, 270.7564, 
    270.7569, 270.7552, 270.7596, 270.7578, 270.7585, 270.7566, 270.7607, 
    270.7574, 270.7615, 270.7612, 270.76, 270.7577, 270.7571, 270.7566, 
    270.7569, 270.7586, 270.7589, 270.76, 270.7604, 270.7612, 270.762, 
    270.7613, 270.7606, 270.7586, 270.7568, 270.7548, 270.7543, 270.752, 
    270.7539, 270.7509, 270.7535, 270.7489, 270.7571, 270.7535, 270.7599, 
    270.7592, 270.758, 270.7551, 270.7567, 270.7549, 270.7589, 270.761, 
    270.7615, 270.7625, 270.7615, 270.7616, 270.7606, 270.7609, 270.7585, 
    270.7598, 270.7562, 270.7549, 270.7511, 270.7488, 270.7465, 270.7454, 
    270.7451, 270.745 ;

 TREFMXAV_R =
  270.7703, 270.7681, 270.7685, 270.7668, 270.7678, 270.7667, 270.7698, 
    270.7681, 270.7692, 270.7701, 270.7636, 270.7668, 270.7602, 270.7622, 
    270.757, 270.7605, 270.7563, 270.7571, 270.7547, 270.7554, 270.7524, 
    270.7544, 270.7508, 270.7528, 270.7525, 270.7545, 270.7661, 270.764, 
    270.7662, 270.7659, 270.7661, 270.7678, 270.7686, 270.7704, 270.7701, 
    270.7688, 270.7658, 270.7668, 270.7642, 270.7643, 270.7614, 270.7627, 
    270.7579, 270.7593, 270.7553, 270.7563, 270.7554, 270.7557, 270.7554, 
    270.7569, 270.7562, 270.7575, 270.7625, 270.761, 270.7654, 270.7681, 
    270.7697, 270.771, 270.7708, 270.7705, 270.7688, 270.7671, 270.7659, 
    270.7651, 270.7643, 270.7619, 270.7606, 270.7577, 270.7582, 270.7573, 
    270.7564, 270.755, 270.7552, 270.7546, 270.7573, 270.7556, 270.7585, 
    270.7577, 270.7642, 270.7665, 270.7676, 270.7685, 270.7707, 270.7691, 
    270.7697, 270.7683, 270.7674, 270.7678, 270.7651, 270.7661, 270.7605, 
    270.7629, 270.7566, 270.7581, 270.7562, 270.7571, 270.7555, 270.757, 
    270.7544, 270.7539, 270.7542, 270.7527, 270.757, 270.7554, 270.7679, 
    270.7678, 270.7674, 270.769, 270.769, 270.7704, 270.7692, 270.7687, 
    270.7673, 270.7666, 270.7658, 270.7642, 270.7624, 270.7598, 270.758, 
    270.7567, 270.7575, 270.7568, 270.7576, 270.7579, 270.7541, 270.7562, 
    270.753, 270.7531, 270.7546, 270.7531, 270.7677, 270.7681, 270.7696, 
    270.7685, 270.7705, 270.7694, 270.7687, 270.7661, 270.7655, 270.765, 
    270.764, 270.7627, 270.7603, 270.7583, 270.7564, 270.7565, 270.7565, 
    270.7561, 270.7571, 270.7559, 270.7557, 270.7562, 270.7532, 270.754, 
    270.7531, 270.7537, 270.768, 270.7673, 270.7677, 270.767, 270.7675, 
    270.7653, 270.7646, 270.7614, 270.7627, 270.7606, 270.7625, 270.7621, 
    270.7606, 270.7624, 270.7584, 270.7611, 270.756, 270.7588, 270.7559, 
    270.7564, 270.7555, 270.7548, 270.7538, 270.752, 270.7524, 270.7509, 
    270.7662, 270.7654, 270.7654, 270.7644, 270.7637, 270.7622, 270.7597, 
    270.7607, 270.7589, 270.7586, 270.7612, 270.7596, 270.7647, 270.7639, 
    270.7644, 270.7662, 270.7605, 270.7634, 270.7579, 270.7596, 270.7549, 
    270.7572, 270.7527, 270.7508, 270.7489, 270.7468, 270.7648, 270.7654, 
    270.7643, 270.7628, 270.7614, 270.7595, 270.7592, 270.7589, 270.758, 
    270.7572, 270.7588, 270.757, 270.7638, 270.7602, 270.7657, 270.7641, 
    270.7629, 270.7634, 270.7607, 270.7601, 270.7576, 270.7589, 270.7513, 
    270.7546, 270.7451, 270.7478, 270.7657, 270.7648, 270.7619, 270.7633, 
    270.7593, 270.7583, 270.7575, 270.7565, 270.7564, 270.7558, 270.7568, 
    270.7558, 270.7594, 270.7578, 270.7622, 270.7612, 270.7617, 270.7622, 
    270.7605, 270.7588, 270.7587, 270.7581, 270.7567, 270.7593, 270.7509, 
    270.7562, 270.7639, 270.7623, 270.7621, 270.7627, 270.7584, 270.76, 
    270.7558, 270.7569, 270.7551, 270.756, 270.7562, 270.7573, 270.7581, 
    270.7599, 270.7614, 270.7626, 270.7623, 270.761, 270.7587, 270.7564, 
    270.7569, 270.7552, 270.7596, 270.7578, 270.7585, 270.7566, 270.7607, 
    270.7574, 270.7615, 270.7612, 270.76, 270.7577, 270.7571, 270.7566, 
    270.7569, 270.7586, 270.7589, 270.76, 270.7604, 270.7612, 270.762, 
    270.7613, 270.7606, 270.7586, 270.7568, 270.7548, 270.7543, 270.752, 
    270.7539, 270.7509, 270.7535, 270.7489, 270.7571, 270.7535, 270.7599, 
    270.7592, 270.758, 270.7551, 270.7567, 270.7549, 270.7589, 270.761, 
    270.7615, 270.7625, 270.7615, 270.7616, 270.7606, 270.7609, 270.7585, 
    270.7598, 270.7562, 270.7549, 270.7511, 270.7488, 270.7465, 270.7454, 
    270.7451, 270.745 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  255.207, 255.2068, 255.2068, 255.2067, 255.2068, 255.2067, 255.2069, 
    255.2068, 255.2069, 255.2069, 255.2064, 255.2067, 255.2062, 255.2063, 
    255.2059, 255.2062, 255.2058, 255.2059, 255.2057, 255.2058, 255.2055, 
    255.2057, 255.2054, 255.2056, 255.2055, 255.2057, 255.2066, 255.2065, 
    255.2066, 255.2066, 255.2066, 255.2068, 255.2068, 255.207, 255.2069, 
    255.2068, 255.2066, 255.2067, 255.2065, 255.2065, 255.2063, 255.2064, 
    255.206, 255.2061, 255.2058, 255.2059, 255.2058, 255.2058, 255.2058, 
    255.2059, 255.2058, 255.2059, 255.2063, 255.2062, 255.2066, 255.2068, 
    255.2069, 255.207, 255.207, 255.207, 255.2068, 255.2067, 255.2066, 
    255.2065, 255.2065, 255.2063, 255.2062, 255.206, 255.206, 255.2059, 
    255.2059, 255.2057, 255.2058, 255.2057, 255.2059, 255.2058, 255.206, 
    255.206, 255.2065, 255.2067, 255.2067, 255.2068, 255.207, 255.2069, 
    255.2069, 255.2068, 255.2067, 255.2068, 255.2065, 255.2066, 255.2062, 
    255.2064, 255.2059, 255.206, 255.2058, 255.2059, 255.2058, 255.2059, 
    255.2057, 255.2056, 255.2057, 255.2056, 255.2059, 255.2058, 255.2068, 
    255.2068, 255.2067, 255.2068, 255.2069, 255.207, 255.2069, 255.2068, 
    255.2067, 255.2067, 255.2066, 255.2065, 255.2063, 255.2061, 255.206, 
    255.2059, 255.2059, 255.2059, 255.2059, 255.206, 255.2057, 255.2058, 
    255.2056, 255.2056, 255.2057, 255.2056, 255.2068, 255.2068, 255.2069, 
    255.2068, 255.207, 255.2069, 255.2068, 255.2066, 255.2066, 255.2065, 
    255.2065, 255.2064, 255.2062, 255.206, 255.2059, 255.2059, 255.2059, 
    255.2058, 255.2059, 255.2058, 255.2058, 255.2058, 255.2056, 255.2057, 
    255.2056, 255.2056, 255.2068, 255.2067, 255.2068, 255.2067, 255.2067, 
    255.2066, 255.2065, 255.2063, 255.2064, 255.2062, 255.2063, 255.2063, 
    255.2062, 255.2063, 255.206, 255.2062, 255.2058, 255.2061, 255.2058, 
    255.2059, 255.2058, 255.2057, 255.2056, 255.2055, 255.2055, 255.2054, 
    255.2066, 255.2066, 255.2066, 255.2065, 255.2065, 255.2063, 255.2061, 
    255.2062, 255.2061, 255.206, 255.2062, 255.2061, 255.2065, 255.2065, 
    255.2065, 255.2066, 255.2062, 255.2064, 255.206, 255.2061, 255.2057, 
    255.2059, 255.2056, 255.2054, 255.2052, 255.2051, 255.2065, 255.2066, 
    255.2065, 255.2064, 255.2063, 255.2061, 255.2061, 255.2061, 255.206, 
    255.2059, 255.2061, 255.2059, 255.2065, 255.2062, 255.2066, 255.2065, 
    255.2064, 255.2064, 255.2062, 255.2062, 255.2059, 255.2061, 255.2054, 
    255.2057, 255.2049, 255.2052, 255.2066, 255.2065, 255.2063, 255.2064, 
    255.2061, 255.206, 255.2059, 255.2059, 255.2059, 255.2058, 255.2059, 
    255.2058, 255.2061, 255.206, 255.2063, 255.2062, 255.2063, 255.2063, 
    255.2062, 255.206, 255.206, 255.206, 255.2059, 255.2061, 255.2054, 
    255.2058, 255.2065, 255.2063, 255.2063, 255.2064, 255.206, 255.2061, 
    255.2058, 255.2059, 255.2057, 255.2058, 255.2058, 255.2059, 255.206, 
    255.2061, 255.2063, 255.2063, 255.2063, 255.2062, 255.206, 255.2059, 
    255.2059, 255.2058, 255.2061, 255.206, 255.206, 255.2059, 255.2062, 
    255.2059, 255.2063, 255.2062, 255.2061, 255.206, 255.2059, 255.2059, 
    255.2059, 255.206, 255.2061, 255.2061, 255.2062, 255.2062, 255.2063, 
    255.2063, 255.2062, 255.206, 255.2059, 255.2057, 255.2057, 255.2055, 
    255.2057, 255.2054, 255.2056, 255.2052, 255.2059, 255.2056, 255.2061, 
    255.2061, 255.206, 255.2057, 255.2059, 255.2057, 255.2061, 255.2062, 
    255.2063, 255.2063, 255.2063, 255.2063, 255.2062, 255.2062, 255.206, 
    255.2061, 255.2058, 255.2057, 255.2054, 255.2052, 255.205, 255.205, 
    255.2049, 255.2049 ;

 TSAI =
  0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173 ;

 TSA_R =
  255.207, 255.2068, 255.2068, 255.2067, 255.2068, 255.2067, 255.2069, 
    255.2068, 255.2069, 255.2069, 255.2064, 255.2067, 255.2062, 255.2063, 
    255.2059, 255.2062, 255.2058, 255.2059, 255.2057, 255.2058, 255.2055, 
    255.2057, 255.2054, 255.2056, 255.2055, 255.2057, 255.2066, 255.2065, 
    255.2066, 255.2066, 255.2066, 255.2068, 255.2068, 255.207, 255.2069, 
    255.2068, 255.2066, 255.2067, 255.2065, 255.2065, 255.2063, 255.2064, 
    255.206, 255.2061, 255.2058, 255.2059, 255.2058, 255.2058, 255.2058, 
    255.2059, 255.2058, 255.2059, 255.2063, 255.2062, 255.2066, 255.2068, 
    255.2069, 255.207, 255.207, 255.207, 255.2068, 255.2067, 255.2066, 
    255.2065, 255.2065, 255.2063, 255.2062, 255.206, 255.206, 255.2059, 
    255.2059, 255.2057, 255.2058, 255.2057, 255.2059, 255.2058, 255.206, 
    255.206, 255.2065, 255.2067, 255.2067, 255.2068, 255.207, 255.2069, 
    255.2069, 255.2068, 255.2067, 255.2068, 255.2065, 255.2066, 255.2062, 
    255.2064, 255.2059, 255.206, 255.2058, 255.2059, 255.2058, 255.2059, 
    255.2057, 255.2056, 255.2057, 255.2056, 255.2059, 255.2058, 255.2068, 
    255.2068, 255.2067, 255.2068, 255.2069, 255.207, 255.2069, 255.2068, 
    255.2067, 255.2067, 255.2066, 255.2065, 255.2063, 255.2061, 255.206, 
    255.2059, 255.2059, 255.2059, 255.2059, 255.206, 255.2057, 255.2058, 
    255.2056, 255.2056, 255.2057, 255.2056, 255.2068, 255.2068, 255.2069, 
    255.2068, 255.207, 255.2069, 255.2068, 255.2066, 255.2066, 255.2065, 
    255.2065, 255.2064, 255.2062, 255.206, 255.2059, 255.2059, 255.2059, 
    255.2058, 255.2059, 255.2058, 255.2058, 255.2058, 255.2056, 255.2057, 
    255.2056, 255.2056, 255.2068, 255.2067, 255.2068, 255.2067, 255.2067, 
    255.2066, 255.2065, 255.2063, 255.2064, 255.2062, 255.2063, 255.2063, 
    255.2062, 255.2063, 255.206, 255.2062, 255.2058, 255.2061, 255.2058, 
    255.2059, 255.2058, 255.2057, 255.2056, 255.2055, 255.2055, 255.2054, 
    255.2066, 255.2066, 255.2066, 255.2065, 255.2065, 255.2063, 255.2061, 
    255.2062, 255.2061, 255.206, 255.2062, 255.2061, 255.2065, 255.2065, 
    255.2065, 255.2066, 255.2062, 255.2064, 255.206, 255.2061, 255.2057, 
    255.2059, 255.2056, 255.2054, 255.2052, 255.2051, 255.2065, 255.2066, 
    255.2065, 255.2064, 255.2063, 255.2061, 255.2061, 255.2061, 255.206, 
    255.2059, 255.2061, 255.2059, 255.2065, 255.2062, 255.2066, 255.2065, 
    255.2064, 255.2064, 255.2062, 255.2062, 255.2059, 255.2061, 255.2054, 
    255.2057, 255.2049, 255.2052, 255.2066, 255.2065, 255.2063, 255.2064, 
    255.2061, 255.206, 255.2059, 255.2059, 255.2059, 255.2058, 255.2059, 
    255.2058, 255.2061, 255.206, 255.2063, 255.2062, 255.2063, 255.2063, 
    255.2062, 255.206, 255.206, 255.206, 255.2059, 255.2061, 255.2054, 
    255.2058, 255.2065, 255.2063, 255.2063, 255.2064, 255.206, 255.2061, 
    255.2058, 255.2059, 255.2057, 255.2058, 255.2058, 255.2059, 255.206, 
    255.2061, 255.2063, 255.2063, 255.2063, 255.2062, 255.206, 255.2059, 
    255.2059, 255.2058, 255.2061, 255.206, 255.206, 255.2059, 255.2062, 
    255.2059, 255.2063, 255.2062, 255.2061, 255.206, 255.2059, 255.2059, 
    255.2059, 255.206, 255.2061, 255.2061, 255.2062, 255.2062, 255.2063, 
    255.2063, 255.2062, 255.206, 255.2059, 255.2057, 255.2057, 255.2055, 
    255.2057, 255.2054, 255.2056, 255.2052, 255.2059, 255.2056, 255.2061, 
    255.2061, 255.206, 255.2057, 255.2059, 255.2057, 255.2061, 255.2062, 
    255.2063, 255.2063, 255.2063, 255.2063, 255.2062, 255.2062, 255.206, 
    255.2061, 255.2058, 255.2057, 255.2054, 255.2052, 255.205, 255.205, 
    255.2049, 255.2049 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  253.6972, 253.699, 253.6987, 253.7002, 253.6994, 253.7003, 253.6976, 
    253.6991, 253.6981, 253.6973, 253.703, 253.7003, 253.7061, 253.7043, 
    253.7088, 253.7058, 253.7095, 253.7088, 253.7109, 253.7103, 253.713, 
    253.7112, 253.7144, 253.7126, 253.7128, 253.7111, 253.7009, 253.7027, 
    253.7007, 253.701, 253.7009, 253.6994, 253.6986, 253.697, 253.6973, 
    253.6985, 253.7011, 253.7002, 253.7025, 253.7025, 253.705, 253.7038, 
    253.7081, 253.7069, 253.7103, 253.7095, 253.7103, 253.7101, 253.7103, 
    253.709, 253.7096, 253.7084, 253.704, 253.7053, 253.7015, 253.6991, 
    253.6976, 253.6965, 253.6967, 253.697, 253.6985, 253.6999, 253.701, 
    253.7017, 253.7025, 253.7045, 253.7057, 253.7083, 253.7078, 253.7086, 
    253.7094, 253.7106, 253.7104, 253.711, 253.7086, 253.7102, 253.7076, 
    253.7083, 253.7025, 253.7005, 253.6995, 253.6987, 253.6968, 253.6981, 
    253.6976, 253.6989, 253.6997, 253.6993, 253.7018, 253.7008, 253.7058, 
    253.7036, 253.7093, 253.7079, 253.7096, 253.7088, 253.7102, 253.7089, 
    253.7112, 253.7117, 253.7113, 253.7126, 253.7088, 253.7103, 253.6993, 
    253.6993, 253.6997, 253.6983, 253.6982, 253.697, 253.6981, 253.6985, 
    253.6998, 253.7004, 253.7011, 253.7025, 253.7041, 253.7064, 253.708, 
    253.7091, 253.7085, 253.709, 253.7084, 253.7081, 253.7115, 253.7095, 
    253.7125, 253.7123, 253.711, 253.7123, 253.6994, 253.699, 253.6977, 
    253.6987, 253.6969, 253.6979, 253.6985, 253.7008, 253.7013, 253.7018, 
    253.7027, 253.7039, 253.7059, 253.7077, 253.7094, 253.7093, 253.7094, 
    253.7097, 253.7088, 253.7099, 253.71, 253.7096, 253.7123, 253.7115, 
    253.7123, 253.7118, 253.6991, 253.6998, 253.6994, 253.7001, 253.6996, 
    253.7016, 253.7022, 253.705, 253.7039, 253.7057, 253.7041, 253.7043, 
    253.7057, 253.7041, 253.7076, 253.7052, 253.7097, 253.7073, 253.7099, 
    253.7094, 253.7102, 253.7109, 253.7117, 253.7133, 253.7129, 253.7143, 
    253.7007, 253.7015, 253.7015, 253.7023, 253.7029, 253.7043, 253.7065, 
    253.7057, 253.7072, 253.7075, 253.7052, 253.7066, 253.7021, 253.7028, 
    253.7024, 253.7008, 253.7058, 253.7032, 253.708, 253.7066, 253.7108, 
    253.7087, 253.7127, 253.7144, 253.7161, 253.7179, 253.702, 253.7014, 
    253.7024, 253.7037, 253.705, 253.7067, 253.7069, 253.7072, 253.708, 
    253.7087, 253.7073, 253.7089, 253.7029, 253.7061, 253.7012, 253.7026, 
    253.7037, 253.7032, 253.7056, 253.7061, 253.7083, 253.7072, 253.714, 
    253.711, 253.7194, 253.717, 253.7012, 253.702, 253.7045, 253.7033, 
    253.7068, 253.7077, 253.7084, 253.7093, 253.7094, 253.7099, 253.7091, 
    253.7099, 253.7067, 253.7081, 253.7043, 253.7052, 253.7048, 253.7043, 
    253.7058, 253.7073, 253.7074, 253.7079, 253.7092, 253.7069, 253.7143, 
    253.7096, 253.7028, 253.7042, 253.7044, 253.7039, 253.7076, 253.7063, 
    253.7099, 253.7089, 253.7106, 253.7098, 253.7096, 253.7086, 253.7079, 
    253.7063, 253.705, 253.7039, 253.7042, 253.7053, 253.7074, 253.7094, 
    253.709, 253.7104, 253.7066, 253.7082, 253.7076, 253.7092, 253.7056, 
    253.7086, 253.7049, 253.7052, 253.7062, 253.7083, 253.7088, 253.7093, 
    253.709, 253.7075, 253.7072, 253.7062, 253.7059, 253.7051, 253.7045, 
    253.7051, 253.7057, 253.7075, 253.7091, 253.7109, 253.7113, 253.7133, 
    253.7116, 253.7143, 253.7119, 253.7161, 253.7088, 253.712, 253.7063, 
    253.7069, 253.708, 253.7105, 253.7092, 253.7108, 253.7072, 253.7054, 
    253.7049, 253.704, 253.7049, 253.7048, 253.7057, 253.7055, 253.7075, 
    253.7064, 253.7096, 253.7108, 253.7141, 253.7161, 253.7183, 253.7192, 
    253.7195, 253.7196,
  255.2279, 255.2296, 255.2293, 255.2307, 255.2299, 255.2308, 255.2282, 
    255.2297, 255.2288, 255.228, 255.2333, 255.2307, 255.2362, 255.2345, 
    255.2387, 255.2359, 255.2393, 255.2387, 255.2407, 255.2401, 255.2426, 
    255.241, 255.244, 255.2422, 255.2425, 255.2409, 255.2313, 255.233, 
    255.2312, 255.2314, 255.2313, 255.2299, 255.2292, 255.2278, 255.228, 
    255.2291, 255.2315, 255.2307, 255.2328, 255.2328, 255.2351, 255.2341, 
    255.238, 255.2369, 255.2401, 255.2393, 255.2401, 255.2399, 255.2401, 
    255.2389, 255.2394, 255.2384, 255.2343, 255.2354, 255.2319, 255.2297, 
    255.2283, 255.2273, 255.2274, 255.2277, 255.2291, 255.2304, 255.2314, 
    255.2321, 255.2328, 255.2347, 255.2358, 255.2382, 255.2378, 255.2385, 
    255.2392, 255.2404, 255.2402, 255.2407, 255.2385, 255.24, 255.2376, 
    255.2382, 255.2328, 255.2309, 255.23, 255.2293, 255.2275, 255.2288, 
    255.2283, 255.2295, 255.2302, 255.2298, 255.2321, 255.2312, 255.2359, 
    255.2339, 255.2392, 255.2379, 255.2395, 255.2387, 255.24, 255.2388, 
    255.2409, 255.2414, 255.2411, 255.2423, 255.2387, 255.2401, 255.2298, 
    255.2299, 255.2302, 255.2289, 255.2289, 255.2277, 255.2287, 255.2292, 
    255.2303, 255.2309, 255.2315, 255.2328, 255.2343, 255.2364, 255.238, 
    255.239, 255.2384, 255.2389, 255.2383, 255.238, 255.2412, 255.2394, 
    255.2421, 255.242, 255.2407, 255.242, 255.2299, 255.2296, 255.2284, 
    255.2293, 255.2276, 255.2286, 255.2291, 255.2312, 255.2317, 255.2321, 
    255.233, 255.2341, 255.236, 255.2377, 255.2393, 255.2392, 255.2392, 
    255.2395, 255.2387, 255.2397, 255.2399, 255.2394, 255.242, 255.2412, 
    255.242, 255.2415, 255.2297, 255.2303, 255.23, 255.2306, 255.2301, 
    255.232, 255.2325, 255.2351, 255.2341, 255.2358, 255.2343, 255.2345, 
    255.2358, 255.2344, 255.2376, 255.2354, 255.2396, 255.2373, 255.2397, 
    255.2393, 255.24, 255.2406, 255.2414, 255.2429, 255.2426, 255.2438, 
    255.2312, 255.2319, 255.2318, 255.2326, 255.2332, 255.2345, 255.2365, 
    255.2358, 255.2372, 255.2375, 255.2353, 255.2366, 255.2324, 255.2331, 
    255.2327, 255.2312, 255.2359, 255.2335, 255.238, 255.2367, 255.2405, 
    255.2386, 255.2424, 255.244, 255.2455, 255.2473, 255.2323, 255.2318, 
    255.2327, 255.234, 255.2352, 255.2368, 255.2369, 255.2372, 255.238, 
    255.2386, 255.2373, 255.2388, 255.2332, 255.2361, 255.2316, 255.2329, 
    255.2339, 255.2335, 255.2357, 255.2362, 255.2383, 255.2372, 255.2436, 
    255.2407, 255.2487, 255.2464, 255.2316, 255.2323, 255.2347, 255.2336, 
    255.2369, 255.2377, 255.2383, 255.2392, 255.2393, 255.2398, 255.239, 
    255.2397, 255.2368, 255.2381, 255.2345, 255.2353, 255.2349, 255.2345, 
    255.2359, 255.2373, 255.2374, 255.2378, 255.239, 255.2369, 255.2439, 
    255.2395, 255.2331, 255.2344, 255.2346, 255.2341, 255.2376, 255.2363, 
    255.2398, 255.2388, 255.2404, 255.2396, 255.2395, 255.2385, 255.2379, 
    255.2364, 255.2351, 255.2342, 255.2344, 255.2355, 255.2374, 255.2393, 
    255.2389, 255.2402, 255.2366, 255.2381, 255.2375, 255.2391, 255.2357, 
    255.2385, 255.235, 255.2353, 255.2363, 255.2382, 255.2387, 255.2391, 
    255.2389, 255.2375, 255.2372, 255.2363, 255.236, 255.2353, 255.2346, 
    255.2352, 255.2358, 255.2375, 255.239, 255.2406, 255.241, 255.2429, 
    255.2413, 255.2439, 255.2417, 255.2455, 255.2387, 255.2417, 255.2363, 
    255.2369, 255.2379, 255.2403, 255.2391, 255.2406, 255.2372, 255.2355, 
    255.2351, 255.2342, 255.2351, 255.235, 255.2358, 255.2356, 255.2375, 
    255.2365, 255.2395, 255.2406, 255.2437, 255.2456, 255.2476, 255.2485, 
    255.2487, 255.2488,
  257.2929, 257.2943, 257.2941, 257.2952, 257.2946, 257.2953, 257.2932, 
    257.2944, 257.2936, 257.2931, 257.2973, 257.2952, 257.2996, 257.2982, 
    257.3017, 257.2994, 257.3022, 257.3017, 257.3033, 257.3028, 257.3049, 
    257.3035, 257.306, 257.3046, 257.3048, 257.3035, 257.2957, 257.2971, 
    257.2956, 257.2958, 257.2957, 257.2946, 257.294, 257.2928, 257.293, 
    257.2939, 257.2959, 257.2952, 257.2969, 257.2969, 257.2988, 257.2979, 
    257.3011, 257.3002, 257.3029, 257.3022, 257.3028, 257.3026, 257.3028, 
    257.3018, 257.3022, 257.3014, 257.2981, 257.299, 257.2961, 257.2944, 
    257.2933, 257.2924, 257.2926, 257.2928, 257.2939, 257.295, 257.2958, 
    257.2963, 257.2969, 257.2984, 257.2993, 257.3013, 257.3009, 257.3015, 
    257.3021, 257.3031, 257.3029, 257.3033, 257.3015, 257.3027, 257.3008, 
    257.3013, 257.2969, 257.2954, 257.2947, 257.2941, 257.2927, 257.2936, 
    257.2932, 257.2942, 257.2948, 257.2945, 257.2964, 257.2956, 257.2994, 
    257.2978, 257.302, 257.301, 257.3023, 257.3016, 257.3028, 257.3018, 
    257.3035, 257.3039, 257.3036, 257.3046, 257.3017, 257.3028, 257.2945, 
    257.2946, 257.2948, 257.2938, 257.2937, 257.2928, 257.2936, 257.2939, 
    257.2949, 257.2953, 257.2958, 257.2969, 257.2981, 257.2998, 257.3011, 
    257.3019, 257.3014, 257.3018, 257.3014, 257.3011, 257.3037, 257.3022, 
    257.3045, 257.3044, 257.3033, 257.3044, 257.2946, 257.2943, 257.2933, 
    257.2941, 257.2927, 257.2935, 257.2939, 257.2956, 257.296, 257.2964, 
    257.2971, 257.2979, 257.2995, 257.3009, 257.3022, 257.3021, 257.3021, 
    257.3024, 257.3017, 257.3025, 257.3026, 257.3023, 257.3044, 257.3037, 
    257.3044, 257.304, 257.2944, 257.2949, 257.2946, 257.2951, 257.2947, 
    257.2962, 257.2967, 257.2988, 257.2979, 257.2993, 257.2981, 257.2983, 
    257.2993, 257.2982, 257.3008, 257.299, 257.3024, 257.3005, 257.3025, 
    257.3022, 257.3027, 257.3033, 257.3039, 257.3051, 257.3048, 257.3059, 
    257.2956, 257.2962, 257.2961, 257.2968, 257.2972, 257.2982, 257.2999, 
    257.2993, 257.3004, 257.3007, 257.2989, 257.3, 257.2966, 257.2971, 
    257.2968, 257.2956, 257.2994, 257.2975, 257.3011, 257.3, 257.3032, 
    257.3016, 257.3047, 257.306, 257.3073, 257.3087, 257.2965, 257.2961, 
    257.2968, 257.2979, 257.2988, 257.3001, 257.3002, 257.3005, 257.3011, 
    257.3016, 257.3005, 257.3018, 257.2972, 257.2996, 257.2959, 257.297, 
    257.2978, 257.2975, 257.2992, 257.2996, 257.3013, 257.3004, 257.3057, 
    257.3033, 257.3099, 257.308, 257.296, 257.2965, 257.2984, 257.2975, 
    257.3002, 257.3008, 257.3014, 257.3021, 257.3022, 257.3026, 257.3019, 
    257.3025, 257.3001, 257.3012, 257.2982, 257.299, 257.2986, 257.2982, 
    257.2994, 257.3005, 257.3006, 257.301, 257.302, 257.3002, 257.3059, 
    257.3023, 257.2971, 257.2982, 257.2983, 257.2979, 257.3008, 257.2997, 
    257.3026, 257.3018, 257.303, 257.3024, 257.3023, 257.3015, 257.301, 
    257.2998, 257.2988, 257.298, 257.2982, 257.299, 257.3006, 257.3021, 
    257.3018, 257.3029, 257.3, 257.3012, 257.3007, 257.302, 257.2993, 
    257.3015, 257.2987, 257.299, 257.2997, 257.3013, 257.3017, 257.302, 
    257.3018, 257.3007, 257.3005, 257.2997, 257.2995, 257.2989, 257.2984, 
    257.2988, 257.2993, 257.3007, 257.3019, 257.3033, 257.3036, 257.3051, 
    257.3038, 257.3059, 257.3041, 257.3073, 257.3017, 257.3041, 257.2998, 
    257.3002, 257.3011, 257.303, 257.302, 257.3032, 257.3005, 257.299, 
    257.2987, 257.298, 257.2987, 257.2987, 257.2993, 257.2991, 257.3007, 
    257.2999, 257.3023, 257.3032, 257.3058, 257.3073, 257.309, 257.3097, 
    257.3099, 257.31,
  259.7985, 259.7993, 259.7992, 259.7998, 259.7995, 259.7999, 259.7987, 
    259.7993, 259.7989, 259.7986, 259.8011, 259.7999, 259.8024, 259.8016, 
    259.8037, 259.8023, 259.804, 259.8037, 259.8047, 259.8044, 259.8056, 
    259.8048, 259.8063, 259.8054, 259.8055, 259.8047, 259.8001, 259.8009, 
    259.8001, 259.8002, 259.8001, 259.7995, 259.7991, 259.7985, 259.7986, 
    259.7991, 259.8002, 259.7998, 259.8008, 259.8008, 259.8019, 259.8014, 
    259.8033, 259.8028, 259.8044, 259.804, 259.8044, 259.8042, 259.8044, 
    259.8038, 259.804, 259.8035, 259.8015, 259.8021, 259.8004, 259.7993, 
    259.7987, 259.7982, 259.7983, 259.7984, 259.7991, 259.7997, 259.8002, 
    259.8005, 259.8008, 259.8018, 259.8023, 259.8034, 259.8032, 259.8036, 
    259.8039, 259.8045, 259.8044, 259.8047, 259.8036, 259.8043, 259.8031, 
    259.8034, 259.8009, 259.8, 259.7995, 259.7992, 259.7984, 259.799, 
    259.7987, 259.7993, 259.7996, 259.7994, 259.8005, 259.8001, 259.8023, 
    259.8013, 259.8039, 259.8033, 259.804, 259.8036, 259.8043, 259.8037, 
    259.8047, 259.805, 259.8048, 259.8055, 259.8037, 259.8044, 259.7994, 
    259.7995, 259.7996, 259.799, 259.799, 259.7985, 259.7989, 259.7991, 
    259.7996, 259.7999, 259.8002, 259.8008, 259.8016, 259.8026, 259.8033, 
    259.8038, 259.8035, 259.8038, 259.8035, 259.8033, 259.8049, 259.804, 
    259.8054, 259.8053, 259.8047, 259.8053, 259.7995, 259.7993, 259.7988, 
    259.7992, 259.7984, 259.7989, 259.7991, 259.8001, 259.8003, 259.8005, 
    259.8009, 259.8015, 259.8024, 259.8032, 259.804, 259.8039, 259.8039, 
    259.8041, 259.8037, 259.8041, 259.8042, 259.804, 259.8053, 259.8049, 
    259.8053, 259.8051, 259.7994, 259.7997, 259.7995, 259.7998, 259.7996, 
    259.8004, 259.8007, 259.8019, 259.8015, 259.8022, 259.8015, 259.8017, 
    259.8022, 259.8016, 259.8031, 259.8021, 259.8041, 259.803, 259.8042, 
    259.804, 259.8043, 259.8046, 259.805, 259.8058, 259.8056, 259.8062, 
    259.8, 259.8004, 259.8004, 259.8008, 259.801, 259.8016, 259.8026, 
    259.8022, 259.8029, 259.8031, 259.802, 259.8026, 259.8007, 259.801, 
    259.8008, 259.8001, 259.8023, 259.8011, 259.8033, 259.8027, 259.8046, 
    259.8036, 259.8055, 259.8063, 259.8071, 259.808, 259.8006, 259.8004, 
    259.8008, 259.8014, 259.802, 259.8027, 259.8028, 259.8029, 259.8033, 
    259.8036, 259.803, 259.8037, 259.801, 259.8024, 259.8003, 259.8009, 
    259.8014, 259.8012, 259.8022, 259.8025, 259.8034, 259.8029, 259.8061, 
    259.8047, 259.8087, 259.8075, 259.8003, 259.8006, 259.8017, 259.8012, 
    259.8028, 259.8032, 259.8035, 259.8039, 259.804, 259.8042, 259.8038, 
    259.8042, 259.8027, 259.8034, 259.8016, 259.802, 259.8018, 259.8016, 
    259.8023, 259.803, 259.803, 259.8033, 259.8038, 259.8028, 259.8062, 
    259.804, 259.801, 259.8016, 259.8017, 259.8015, 259.8031, 259.8025, 
    259.8042, 259.8037, 259.8045, 259.8041, 259.804, 259.8036, 259.8033, 
    259.8026, 259.8019, 259.8015, 259.8016, 259.8021, 259.803, 259.804, 
    259.8037, 259.8044, 259.8027, 259.8034, 259.8031, 259.8039, 259.8022, 
    259.8036, 259.8019, 259.802, 259.8025, 259.8034, 259.8036, 259.8039, 
    259.8037, 259.8031, 259.8029, 259.8025, 259.8024, 259.802, 259.8017, 
    259.802, 259.8022, 259.8031, 259.8038, 259.8046, 259.8048, 259.8058, 
    259.805, 259.8062, 259.8051, 259.8071, 259.8037, 259.8051, 259.8025, 
    259.8028, 259.8033, 259.8045, 259.8039, 259.8046, 259.8029, 259.8021, 
    259.8019, 259.8015, 259.8019, 259.8019, 259.8023, 259.8022, 259.8031, 
    259.8026, 259.804, 259.8046, 259.8061, 259.8071, 259.8081, 259.8085, 
    259.8087, 259.8087,
  262.0123, 262.0125, 262.0125, 262.0127, 262.0126, 262.0127, 262.0124, 
    262.0125, 262.0124, 262.0124, 262.013, 262.0127, 262.0133, 262.0131, 
    262.0137, 262.0133, 262.0138, 262.0137, 262.0139, 262.0139, 262.0142, 
    262.014, 262.0144, 262.0142, 262.0142, 262.014, 262.0127, 262.0129, 
    262.0127, 262.0128, 262.0127, 262.0126, 262.0125, 262.0123, 262.0124, 
    262.0125, 262.0128, 262.0127, 262.0129, 262.0129, 262.0132, 262.0131, 
    262.0136, 262.0134, 262.0139, 262.0138, 262.0139, 262.0138, 262.0139, 
    262.0137, 262.0138, 262.0136, 262.0131, 262.0132, 262.0128, 262.0125, 
    262.0124, 262.0123, 262.0123, 262.0123, 262.0125, 262.0126, 262.0128, 
    262.0128, 262.0129, 262.0132, 262.0133, 262.0136, 262.0135, 262.0136, 
    262.0138, 262.0139, 262.0139, 262.0139, 262.0136, 262.0139, 262.0135, 
    262.0136, 262.0129, 262.0127, 262.0126, 262.0125, 262.0123, 262.0124, 
    262.0124, 262.0125, 262.0126, 262.0125, 262.0128, 262.0127, 262.0133, 
    262.0131, 262.0137, 262.0136, 262.0138, 262.0137, 262.0139, 262.0137, 
    262.014, 262.014, 262.014, 262.0142, 262.0137, 262.0139, 262.0125, 
    262.0126, 262.0126, 262.0125, 262.0125, 262.0123, 262.0124, 262.0125, 
    262.0126, 262.0127, 262.0128, 262.0129, 262.0131, 262.0134, 262.0136, 
    262.0137, 262.0136, 262.0137, 262.0136, 262.0136, 262.014, 262.0138, 
    262.0142, 262.0141, 262.0139, 262.0141, 262.0126, 262.0125, 262.0124, 
    262.0125, 262.0123, 262.0124, 262.0125, 262.0127, 262.0128, 262.0128, 
    262.0129, 262.0131, 262.0133, 262.0135, 262.0138, 262.0137, 262.0137, 
    262.0138, 262.0137, 262.0138, 262.0138, 262.0138, 262.0141, 262.014, 
    262.0141, 262.0141, 262.0125, 262.0126, 262.0126, 262.0126, 262.0126, 
    262.0128, 262.0129, 262.0132, 262.0131, 262.0133, 262.0131, 262.0131, 
    262.0133, 262.0131, 262.0135, 262.0132, 262.0138, 262.0135, 262.0138, 
    262.0138, 262.0139, 262.0139, 262.0141, 262.0143, 262.0142, 262.0144, 
    262.0127, 262.0128, 262.0128, 262.0129, 262.013, 262.0131, 262.0134, 
    262.0133, 262.0135, 262.0135, 262.0132, 262.0134, 262.0129, 262.0129, 
    262.0129, 262.0127, 262.0133, 262.013, 262.0136, 262.0134, 262.0139, 
    262.0137, 262.0142, 262.0144, 262.0146, 262.0149, 262.0128, 262.0128, 
    262.0129, 262.0131, 262.0132, 262.0134, 262.0134, 262.0135, 262.0136, 
    262.0137, 262.0135, 262.0137, 262.013, 262.0133, 262.0128, 262.0129, 
    262.0131, 262.013, 262.0133, 262.0133, 262.0136, 262.0135, 262.0143, 
    262.0139, 262.0151, 262.0148, 262.0128, 262.0128, 262.0132, 262.013, 
    262.0134, 262.0135, 262.0136, 262.0137, 262.0138, 262.0138, 262.0137, 
    262.0138, 262.0134, 262.0136, 262.0131, 262.0132, 262.0132, 262.0131, 
    262.0133, 262.0135, 262.0135, 262.0135, 262.0137, 262.0134, 262.0144, 
    262.0138, 262.0129, 262.0131, 262.0132, 262.0131, 262.0135, 262.0134, 
    262.0138, 262.0137, 262.0139, 262.0138, 262.0138, 262.0136, 262.0136, 
    262.0134, 262.0132, 262.0131, 262.0131, 262.0132, 262.0135, 262.0138, 
    262.0137, 262.0139, 262.0134, 262.0136, 262.0135, 262.0137, 262.0133, 
    262.0136, 262.0132, 262.0132, 262.0134, 262.0136, 262.0137, 262.0137, 
    262.0137, 262.0135, 262.0135, 262.0134, 262.0133, 262.0132, 262.0132, 
    262.0132, 262.0133, 262.0135, 262.0137, 262.0139, 262.014, 262.0143, 
    262.014, 262.0144, 262.0141, 262.0146, 262.0137, 262.0141, 262.0134, 
    262.0134, 262.0136, 262.0139, 262.0137, 262.0139, 262.0135, 262.0132, 
    262.0132, 262.0131, 262.0132, 262.0132, 262.0133, 262.0133, 262.0135, 
    262.0134, 262.0138, 262.0139, 262.0144, 262.0146, 262.015, 262.0151, 
    262.0151, 262.0151,
  262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993,
  263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.1108, 263.1231, 263.1208, 263.1306, 263.1252, 263.1316, 263.1133, 
    263.1236, 263.1171, 263.112, 263.1497, 263.1311, 263.1691, 263.1572, 
    263.187, 263.1672, 263.1909, 263.1864, 263.1999, 263.196, 263.2133, 
    263.2017, 263.2222, 263.2105, 263.2123, 263.2013, 263.1349, 263.1474, 
    263.1341, 263.1359, 263.1351, 263.1253, 263.1203, 263.1099, 263.1118, 
    263.1194, 263.1367, 263.1309, 263.1456, 263.1453, 263.1616, 263.1542, 
    263.1817, 263.1739, 263.1962, 263.1906, 263.196, 263.1943, 263.196, 
    263.1878, 263.1913, 263.1841, 263.1556, 263.164, 263.139, 263.1238, 
    263.1138, 263.1066, 263.1076, 263.1096, 263.1195, 263.1288, 263.1359, 
    263.1406, 263.1452, 263.1592, 263.1667, 263.1832, 263.1803, 263.1853, 
    263.1901, 263.1981, 263.1968, 263.2003, 263.1852, 263.1952, 263.1786, 
    263.1832, 263.1464, 263.1324, 263.1264, 263.1212, 263.1084, 263.1172, 
    263.1138, 263.1221, 263.1273, 263.1247, 263.1407, 263.1345, 263.1671, 
    263.1531, 263.1895, 263.1809, 263.1916, 263.1862, 263.1955, 263.1871, 
    263.2016, 263.2047, 263.2026, 263.2109, 263.1866, 263.196, 263.1247, 
    263.1251, 263.127, 263.1183, 263.1178, 263.1099, 263.1169, 263.12, 
    263.1276, 263.1321, 263.1364, 263.1458, 263.1563, 263.1709, 263.1814, 
    263.1884, 263.1842, 263.1879, 263.1837, 263.1817, 263.2036, 263.1913, 
    263.2097, 263.2087, 263.2004, 263.2088, 263.1254, 263.1229, 263.1144, 
    263.1211, 263.109, 263.1158, 263.1196, 263.1346, 263.1379, 263.1409, 
    263.1469, 263.1546, 263.1681, 263.1798, 263.1904, 263.1896, 263.1899, 
    263.1922, 263.1864, 263.1932, 263.1943, 263.1913, 263.2086, 263.2036, 
    263.2087, 263.2055, 263.1237, 263.1278, 263.1256, 263.1298, 263.1268, 
    263.1398, 263.1437, 263.1619, 263.1545, 263.1663, 263.1557, 263.1576, 
    263.1667, 263.1562, 263.1791, 263.1636, 263.1923, 263.1769, 263.1933, 
    263.1903, 263.1952, 263.1996, 263.205, 263.2151, 263.2128, 263.2212, 
    263.1339, 263.1392, 263.1388, 263.1443, 263.1484, 263.1573, 263.1714, 
    263.1661, 263.1759, 263.1779, 263.163, 263.1721, 263.1428, 263.1475, 
    263.1447, 263.1343, 263.1673, 263.1504, 263.1816, 263.1725, 263.1989, 
    263.1858, 263.2115, 263.2224, 263.2327, 263.2447, 263.1421, 263.1385, 
    263.145, 263.1538, 263.1621, 263.173, 263.1742, 263.1762, 263.1815, 
    263.1859, 263.1768, 263.187, 263.1485, 263.1688, 263.1371, 263.1467, 
    263.1533, 263.1504, 263.1655, 263.1691, 263.1834, 263.176, 263.2197, 
    263.2004, 263.2538, 263.2389, 263.1373, 263.1421, 263.1589, 263.1509, 
    263.1738, 263.1794, 263.1839, 263.1897, 263.1903, 263.1937, 263.1881, 
    263.1935, 263.1731, 263.1823, 263.157, 263.1631, 263.1603, 263.1572, 
    263.1668, 263.177, 263.1772, 263.1805, 263.1895, 263.1739, 263.2221, 
    263.1924, 263.1474, 263.1566, 263.158, 263.1544, 263.1788, 263.17, 
    263.1936, 263.1873, 263.1977, 263.1925, 263.1918, 263.1851, 263.181, 
    263.1704, 263.1618, 263.1549, 263.1565, 263.164, 263.1776, 263.1904, 
    263.1876, 263.1969, 263.1721, 263.1826, 263.1785, 263.189, 263.166, 
    263.1855, 263.1609, 263.1631, 263.1698, 263.1833, 263.1862, 263.1894, 
    263.1874, 263.1779, 263.1764, 263.1696, 263.1678, 263.1626, 263.1584, 
    263.1623, 263.1664, 263.1779, 263.1884, 263.1996, 263.2024, 263.2154, 
    263.2047, 263.2223, 263.2073, 263.2332, 263.1867, 263.2069, 263.1701, 
    263.1741, 263.1813, 263.1978, 263.189, 263.1993, 263.1764, 263.1643, 
    263.1612, 263.1553, 263.1613, 263.1608, 263.1665, 263.1647, 263.1783, 
    263.171, 263.1917, 263.1992, 263.2203, 263.2332, 263.2464, 263.2522, 
    263.2539, 263.2547 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.5952, 253.596, 253.5959, 253.5965, 253.5961, 253.5966, 253.5954, 
    253.596, 253.5956, 253.5953, 253.5977, 253.5965, 253.599, 253.5983, 
    253.6002, 253.5989, 253.6004, 253.6002, 253.6011, 253.6008, 253.6019, 
    253.6012, 253.6025, 253.6017, 253.6019, 253.6012, 253.5968, 253.5976, 
    253.5967, 253.5968, 253.5968, 253.5961, 253.5958, 253.5952, 253.5953, 
    253.5958, 253.5969, 253.5965, 253.5975, 253.5975, 253.5985, 253.5981, 
    253.5998, 253.5993, 253.6008, 253.6004, 253.6008, 253.6007, 253.6008, 
    253.6003, 253.6005, 253.6, 253.5981, 253.5987, 253.597, 253.596, 
    253.5954, 253.5949, 253.595, 253.5951, 253.5958, 253.5964, 253.5968, 
    253.5972, 253.5975, 253.5983, 253.5988, 253.5999, 253.5997, 253.6001, 
    253.6004, 253.6009, 253.6008, 253.6011, 253.6001, 253.6007, 253.5996, 
    253.5999, 253.5975, 253.5966, 253.5962, 253.5959, 253.595, 253.5956, 
    253.5954, 253.5959, 253.5963, 253.5961, 253.5972, 253.5968, 253.5989, 
    253.598, 253.6004, 253.5998, 253.6005, 253.6001, 253.6008, 253.6002, 
    253.6012, 253.6014, 253.6012, 253.6018, 253.6002, 253.6008, 253.5961, 
    253.5961, 253.5963, 253.5957, 253.5957, 253.5951, 253.5956, 253.5958, 
    253.5963, 253.5966, 253.5969, 253.5975, 253.5982, 253.5991, 253.5998, 
    253.6003, 253.6, 253.6003, 253.6, 253.5999, 253.6013, 253.6005, 253.6017, 
    253.6016, 253.6011, 253.6016, 253.5962, 253.596, 253.5954, 253.5959, 
    253.5951, 253.5955, 253.5958, 253.5968, 253.597, 253.5972, 253.5976, 
    253.5981, 253.599, 253.5997, 253.6004, 253.6004, 253.6004, 253.6005, 
    253.6002, 253.6006, 253.6007, 253.6005, 253.6016, 253.6013, 253.6016, 
    253.6014, 253.5961, 253.5963, 253.5962, 253.5965, 253.5963, 253.5971, 
    253.5974, 253.5985, 253.5981, 253.5988, 253.5981, 253.5983, 253.5988, 
    253.5982, 253.5997, 253.5986, 253.6005, 253.5995, 253.6006, 253.6004, 
    253.6007, 253.601, 253.6014, 253.6021, 253.6019, 253.6025, 253.5967, 
    253.5971, 253.597, 253.5974, 253.5977, 253.5983, 253.5992, 253.5988, 
    253.5995, 253.5996, 253.5986, 253.5992, 253.5973, 253.5976, 253.5974, 
    253.5967, 253.5989, 253.5978, 253.5998, 253.5992, 253.601, 253.6001, 
    253.6018, 253.6025, 253.6032, 253.604, 253.5973, 253.597, 253.5974, 
    253.598, 253.5986, 253.5993, 253.5993, 253.5995, 253.5998, 253.6001, 
    253.5995, 253.6002, 253.5977, 253.599, 253.5969, 253.5975, 253.598, 
    253.5978, 253.5988, 253.599, 253.5999, 253.5995, 253.6023, 253.6011, 
    253.6046, 253.6036, 253.5969, 253.5973, 253.5984, 253.5978, 253.5993, 
    253.5997, 253.6, 253.6004, 253.6004, 253.6006, 253.6003, 253.6006, 
    253.5993, 253.5999, 253.5982, 253.5986, 253.5984, 253.5983, 253.5989, 
    253.5995, 253.5995, 253.5998, 253.6003, 253.5993, 253.6025, 253.6005, 
    253.5976, 253.5982, 253.5983, 253.5981, 253.5997, 253.5991, 253.6006, 
    253.6002, 253.6009, 253.6006, 253.6005, 253.6001, 253.5998, 253.5991, 
    253.5985, 253.5981, 253.5982, 253.5987, 253.5996, 253.6004, 253.6002, 
    253.6008, 253.5992, 253.5999, 253.5996, 253.6003, 253.5988, 253.6001, 
    253.5985, 253.5986, 253.5991, 253.5999, 253.6001, 253.6003, 253.6002, 
    253.5996, 253.5995, 253.5991, 253.5989, 253.5986, 253.5983, 253.5986, 
    253.5988, 253.5996, 253.6003, 253.601, 253.6012, 253.6021, 253.6013, 
    253.6025, 253.6015, 253.6032, 253.6001, 253.6015, 253.5991, 253.5993, 
    253.5998, 253.6009, 253.6003, 253.601, 253.5995, 253.5987, 253.5985, 
    253.5981, 253.5985, 253.5985, 253.5989, 253.5987, 253.5996, 253.5992, 
    253.6005, 253.601, 253.6024, 253.6033, 253.6041, 253.6045, 253.6046, 
    253.6047 ;

 TWS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 T_SCALAR =
  0.145703, 0.145702, 0.1457022, 0.1457013, 0.1457018, 0.1457012, 0.1457028, 
    0.1457019, 0.1457025, 0.1457029, 0.1456998, 0.1457013, 0.1456983, 
    0.1456992, 0.145697, 0.1456984, 0.1456967, 0.145697, 0.1456961, 
    0.1456963, 0.1456952, 0.145696, 0.1456947, 0.1456954, 0.1456953, 
    0.145696, 0.145701, 0.1457, 0.145701, 0.1457009, 0.145701, 0.1457018, 
    0.1457022, 0.1457031, 0.1457029, 0.1457023, 0.1457008, 0.1457013, 
    0.1457001, 0.1457001, 0.1456989, 0.1456994, 0.1456973, 0.1456979, 
    0.1456963, 0.1456967, 0.1456964, 0.1456965, 0.1456964, 0.1456969, 
    0.1456967, 0.1456972, 0.1456993, 0.1456987, 0.1457006, 0.1457019, 
    0.1457027, 0.1457034, 0.1457033, 0.1457031, 0.1457023, 0.1457015, 
    0.1457009, 0.1457005, 0.1457001, 0.1456991, 0.1456985, 0.1456972, 
    0.1456974, 0.1456971, 0.1456968, 0.1456962, 0.1456963, 0.1456961, 
    0.1456971, 0.1456964, 0.1456976, 0.1456972, 0.1457001, 0.1457012, 
    0.1457017, 0.1457021, 0.1457032, 0.1457025, 0.1457027, 0.145702, 
    0.1457016, 0.1457018, 0.1457005, 0.145701, 0.1456985, 0.1456995, 
    0.1456968, 0.1456974, 0.1456967, 0.145697, 0.1456964, 0.145697, 0.145696, 
    0.1456958, 0.1456959, 0.1456954, 0.145697, 0.1456964, 0.1457018, 
    0.1457018, 0.1457016, 0.1457024, 0.1457024, 0.1457031, 0.1457025, 
    0.1457022, 0.1457016, 0.1457012, 0.1457009, 0.1457001, 0.1456993, 
    0.1456982, 0.1456974, 0.1456969, 0.1456972, 0.1456969, 0.1456972, 
    0.1456973, 0.1456959, 0.1456967, 0.1456954, 0.1456955, 0.1456961, 
    0.1456955, 0.1457018, 0.145702, 0.1457027, 0.1457021, 0.1457032, 
    0.1457026, 0.1457023, 0.145701, 0.1457007, 0.1457005, 0.1457, 0.1456994, 
    0.1456984, 0.1456975, 0.1456967, 0.1456968, 0.1456968, 0.1456966, 
    0.145697, 0.1456966, 0.1456965, 0.1456967, 0.1456955, 0.1456958, 
    0.1456955, 0.1456957, 0.1457019, 0.1457016, 0.1457018, 0.1457014, 
    0.1457016, 0.1457006, 0.1457003, 0.1456988, 0.1456994, 0.1456985, 
    0.1456993, 0.1456992, 0.1456985, 0.1456993, 0.1456975, 0.1456987, 
    0.1456966, 0.1456977, 0.1456965, 0.1456967, 0.1456964, 0.1456961, 
    0.1456957, 0.1456951, 0.1456953, 0.1456947, 0.1457011, 0.1457006, 
    0.1457007, 0.1457002, 0.1456999, 0.1456992, 0.1456981, 0.1456985, 
    0.1456978, 0.1456976, 0.1456988, 0.1456981, 0.1457003, 0.1457, 0.1457002, 
    0.145701, 0.1456984, 0.1456997, 0.1456974, 0.145698, 0.1456961, 
    0.1456971, 0.1456953, 0.1456947, 0.1456941, 0.1456934, 0.1457004, 
    0.1457007, 0.1457002, 0.1456995, 0.1456988, 0.145698, 0.1456979, 
    0.1456978, 0.1456974, 0.145697, 0.1456977, 0.145697, 0.1456999, 
    0.1456983, 0.1457008, 0.1457, 0.1456995, 0.1456997, 0.1456986, 0.1456983, 
    0.1456972, 0.1456978, 0.1456948, 0.1456961, 0.145693, 0.1456937, 
    0.1457008, 0.1457004, 0.1456991, 0.1456997, 0.145698, 0.1456975, 
    0.1456972, 0.1456968, 0.1456967, 0.1456965, 0.1456969, 0.1456965, 
    0.145698, 0.1456973, 0.1456992, 0.1456987, 0.145699, 0.1456992, 
    0.1456985, 0.1456977, 0.1456977, 0.1456974, 0.1456968, 0.1456979, 
    0.1456947, 0.1456966, 0.1457, 0.1456992, 0.1456991, 0.1456994, 0.1456975, 
    0.1456982, 0.1456965, 0.145697, 0.1456962, 0.1456966, 0.1456966, 
    0.1456971, 0.1456974, 0.1456982, 0.1456988, 0.1456994, 0.1456992, 
    0.1456987, 0.1456976, 0.1456967, 0.1456969, 0.1456963, 0.1456981, 
    0.1456973, 0.1456976, 0.1456968, 0.1456985, 0.1456971, 0.1456989, 
    0.1456987, 0.1456982, 0.1456972, 0.145697, 0.1456968, 0.1456969, 
    0.1456976, 0.1456978, 0.1456982, 0.1456984, 0.1456988, 0.1456991, 
    0.1456988, 0.1456985, 0.1456976, 0.1456969, 0.1456961, 0.1456959, 
    0.1456951, 0.1456958, 0.1456947, 0.1456956, 0.145694, 0.145697, 
    0.1456956, 0.1456982, 0.1456979, 0.1456974, 0.1456962, 0.1456968, 
    0.1456961, 0.1456978, 0.1456987, 0.1456989, 0.1456993, 0.1456989, 
    0.1456989, 0.1456985, 0.1456986, 0.1456976, 0.1456981, 0.1456966, 
    0.1456961, 0.1456948, 0.145694, 0.1456933, 0.145693, 0.145693, 0.1456929,
  0.1513271, 0.1513317, 0.1513308, 0.1513345, 0.1513325, 0.1513349, 
    0.1513281, 0.1513319, 0.1513295, 0.1513276, 0.1513415, 0.1513347, 
    0.151349, 0.1513445, 0.1513558, 0.1513482, 0.1513574, 0.1513557, 
    0.151361, 0.1513595, 0.1513661, 0.1513617, 0.1513697, 0.1513651, 
    0.1513658, 0.1513615, 0.1513361, 0.1513406, 0.1513358, 0.1513365, 
    0.1513362, 0.1513325, 0.1513306, 0.1513269, 0.1513276, 0.1513303, 
    0.1513368, 0.1513346, 0.1513402, 0.1513401, 0.1513462, 0.1513434, 
    0.1513538, 0.1513509, 0.1513595, 0.1513573, 0.1513594, 0.1513588, 
    0.1513594, 0.1513562, 0.1513576, 0.1513548, 0.1513439, 0.1513471, 
    0.1513376, 0.1513319, 0.1513283, 0.1513256, 0.151326, 0.1513267, 
    0.1513304, 0.1513339, 0.1513365, 0.1513383, 0.15134, 0.1513451, 0.151348, 
    0.1513544, 0.1513533, 0.1513552, 0.1513571, 0.1513602, 0.1513597, 
    0.1513611, 0.1513552, 0.1513591, 0.1513527, 0.1513544, 0.1513402, 
    0.1513352, 0.1513329, 0.151331, 0.1513263, 0.1513295, 0.1513283, 
    0.1513314, 0.1513333, 0.1513323, 0.1513383, 0.151336, 0.1513482, 
    0.1513429, 0.1513569, 0.1513535, 0.1513577, 0.1513556, 0.1513592, 
    0.1513559, 0.1513616, 0.1513628, 0.151362, 0.1513653, 0.1513558, 
    0.1513594, 0.1513323, 0.1513325, 0.1513332, 0.1513299, 0.1513297, 
    0.1513268, 0.1513294, 0.1513305, 0.1513334, 0.1513351, 0.1513367, 
    0.1513402, 0.1513441, 0.1513497, 0.1513537, 0.1513565, 0.1513548, 
    0.1513563, 0.1513546, 0.1513539, 0.1513624, 0.1513576, 0.1513648, 
    0.1513644, 0.1513611, 0.1513645, 0.1513326, 0.1513317, 0.1513285, 
    0.151331, 0.1513265, 0.151329, 0.1513304, 0.151336, 0.1513373, 0.1513384, 
    0.1513407, 0.1513436, 0.1513486, 0.1513531, 0.1513572, 0.1513569, 
    0.151357, 0.1513579, 0.1513557, 0.1513583, 0.1513587, 0.1513576, 
    0.1513644, 0.1513624, 0.1513644, 0.1513632, 0.151332, 0.1513335, 
    0.1513327, 0.1513342, 0.1513331, 0.1513379, 0.1513394, 0.1513462, 
    0.1513435, 0.151348, 0.151344, 0.1513446, 0.151348, 0.1513442, 0.1513528, 
    0.1513468, 0.151358, 0.1513519, 0.1513584, 0.1513572, 0.1513591, 
    0.1513608, 0.151363, 0.1513669, 0.151366, 0.1513694, 0.1513358, 
    0.1513377, 0.1513376, 0.1513397, 0.1513412, 0.1513446, 0.1513499, 
    0.1513479, 0.1513517, 0.1513524, 0.1513467, 0.1513502, 0.1513391, 
    0.1513408, 0.1513398, 0.1513359, 0.1513483, 0.1513419, 0.1513538, 
    0.1513503, 0.1513606, 0.1513554, 0.1513655, 0.1513698, 0.151374, 
    0.1513787, 0.1513388, 0.1513375, 0.1513399, 0.1513432, 0.1513464, 
    0.1513505, 0.151351, 0.1513518, 0.1513538, 0.1513555, 0.151352, 
    0.1513559, 0.1513411, 0.1513489, 0.151337, 0.1513405, 0.151343, 0.151342, 
    0.1513477, 0.151349, 0.1513545, 0.1513517, 0.1513686, 0.1513611, 
    0.1513825, 0.1513764, 0.151337, 0.1513389, 0.1513451, 0.1513422, 
    0.1513508, 0.1513529, 0.1513547, 0.1513569, 0.1513572, 0.1513585, 
    0.1513564, 0.1513584, 0.1513505, 0.1513541, 0.1513445, 0.1513468, 
    0.1513457, 0.1513446, 0.1513482, 0.151352, 0.1513521, 0.1513533, 
    0.1513566, 0.1513509, 0.1513695, 0.1513578, 0.1513408, 0.1513443, 
    0.1513448, 0.1513435, 0.1513527, 0.1513494, 0.1513585, 0.151356, 
    0.1513601, 0.1513581, 0.1513578, 0.1513552, 0.1513536, 0.1513495, 
    0.1513463, 0.1513437, 0.1513443, 0.1513471, 0.1513522, 0.1513572, 
    0.1513561, 0.1513598, 0.1513502, 0.1513541, 0.1513526, 0.1513567, 
    0.1513478, 0.1513551, 0.151346, 0.1513468, 0.1513493, 0.1513544, 
    0.1513556, 0.1513568, 0.1513561, 0.1513524, 0.1513518, 0.1513493, 
    0.1513485, 0.1513466, 0.151345, 0.1513464, 0.151348, 0.1513524, 
    0.1513564, 0.1513608, 0.1513619, 0.1513669, 0.1513627, 0.1513695, 
    0.1513636, 0.151374, 0.1513557, 0.1513636, 0.1513495, 0.151351, 
    0.1513536, 0.15136, 0.1513567, 0.1513606, 0.1513518, 0.1513471, 
    0.1513461, 0.1513438, 0.1513461, 0.1513459, 0.1513481, 0.1513474, 
    0.1513526, 0.1513498, 0.1513577, 0.1513606, 0.151369, 0.1513741, 
    0.1513795, 0.1513818, 0.1513826, 0.1513829,
  0.1611689, 0.1611748, 0.1611737, 0.1611784, 0.1611758, 0.1611789, 
    0.1611702, 0.161175, 0.161172, 0.1611695, 0.1611875, 0.1611786, 
    0.1611972, 0.1611914, 0.1612061, 0.1611962, 0.1612081, 0.1612059, 
    0.1612128, 0.1612108, 0.1612195, 0.1612137, 0.1612242, 0.1612181, 
    0.161219, 0.1612135, 0.1611805, 0.1611864, 0.1611801, 0.161181, 
    0.1611806, 0.1611759, 0.1611734, 0.1611686, 0.1611695, 0.161173, 
    0.1611814, 0.1611786, 0.1611858, 0.1611856, 0.1611935, 0.16119, 
    0.1612035, 0.1611996, 0.1612109, 0.161208, 0.1612107, 0.1612099, 
    0.1612107, 0.1612066, 0.1612083, 0.1612047, 0.1611906, 0.1611947, 
    0.1611825, 0.161175, 0.1611704, 0.161167, 0.1611675, 0.1611684, 
    0.1611731, 0.1611776, 0.161181, 0.1611833, 0.1611856, 0.1611922, 
    0.1611959, 0.1612042, 0.1612028, 0.1612053, 0.1612077, 0.1612118, 
    0.1612111, 0.1612129, 0.1612053, 0.1612103, 0.161202, 0.1612042, 
    0.1611859, 0.1611793, 0.1611763, 0.1611739, 0.1611678, 0.161172, 
    0.1611704, 0.1611744, 0.1611769, 0.1611757, 0.1611834, 0.1611803, 
    0.1611962, 0.1611893, 0.1612075, 0.1612031, 0.1612085, 0.1612058, 
    0.1612104, 0.1612062, 0.1612136, 0.1612152, 0.1612141, 0.1612184, 
    0.161206, 0.1612107, 0.1611756, 0.1611758, 0.1611768, 0.1611725, 
    0.1611723, 0.1611685, 0.1611719, 0.1611733, 0.161177, 0.1611792, 
    0.1611813, 0.1611858, 0.1611909, 0.1611981, 0.1612034, 0.1612069, 
    0.1612048, 0.1612066, 0.1612045, 0.1612035, 0.1612146, 0.1612083, 
    0.1612178, 0.1612173, 0.161213, 0.1612173, 0.1611759, 0.1611748, 
    0.1611707, 0.1611739, 0.1611681, 0.1611713, 0.1611731, 0.1611803, 
    0.161182, 0.1611834, 0.1611864, 0.1611901, 0.1611967, 0.1612025, 
    0.1612079, 0.1612075, 0.1612076, 0.1612088, 0.1612059, 0.1612093, 
    0.1612099, 0.1612084, 0.1612172, 0.1612147, 0.1612173, 0.1612156, 
    0.1611752, 0.1611771, 0.1611761, 0.161178, 0.1611766, 0.1611829, 
    0.1611847, 0.1611936, 0.16119, 0.1611958, 0.1611907, 0.1611916, 
    0.1611959, 0.161191, 0.1612021, 0.1611944, 0.1612089, 0.161201, 
    0.1612093, 0.1612079, 0.1612104, 0.1612125, 0.1612154, 0.1612205, 
    0.1612193, 0.1612237, 0.1611801, 0.1611826, 0.1611824, 0.1611851, 
    0.1611871, 0.1611914, 0.1611984, 0.1611958, 0.1612006, 0.1612016, 
    0.1611943, 0.1611987, 0.1611843, 0.1611866, 0.1611853, 0.1611802, 
    0.1611963, 0.161188, 0.1612034, 0.1611989, 0.1612122, 0.1612055, 
    0.1612187, 0.1612242, 0.1612297, 0.1612359, 0.161184, 0.1611823, 
    0.1611854, 0.1611897, 0.1611938, 0.1611992, 0.1611998, 0.1612008, 
    0.1612034, 0.1612056, 0.161201, 0.1612062, 0.161187, 0.1611971, 
    0.1611816, 0.1611862, 0.1611895, 0.1611881, 0.1611955, 0.1611972, 
    0.1612043, 0.1612007, 0.1612228, 0.1612129, 0.1612408, 0.1612329, 
    0.1611817, 0.161184, 0.1611922, 0.1611883, 0.1611996, 0.1612023, 
    0.1612047, 0.1612075, 0.1612079, 0.1612096, 0.1612068, 0.1612095, 
    0.1611992, 0.1612038, 0.1611913, 0.1611943, 0.161193, 0.1611914, 
    0.1611961, 0.1612011, 0.1612013, 0.1612029, 0.1612071, 0.1611996, 
    0.1612239, 0.1612086, 0.1611866, 0.161191, 0.1611918, 0.16119, 0.1612021, 
    0.1611977, 0.1612095, 0.1612063, 0.1612116, 0.161209, 0.1612086, 
    0.1612052, 0.1612031, 0.1611979, 0.1611936, 0.1611903, 0.1611911, 
    0.1611947, 0.1612014, 0.1612079, 0.1612064, 0.1612112, 0.1611988, 
    0.1612039, 0.1612019, 0.1612072, 0.1611957, 0.1612052, 0.1611933, 
    0.1611943, 0.1611976, 0.1612042, 0.1612058, 0.1612073, 0.1612064, 
    0.1612016, 0.1612009, 0.1611975, 0.1611966, 0.1611941, 0.161192, 
    0.1611939, 0.1611959, 0.1612016, 0.1612068, 0.1612126, 0.161214, 
    0.1612205, 0.1612151, 0.1612239, 0.1612162, 0.1612297, 0.1612059, 
    0.1612162, 0.1611978, 0.1611998, 0.1612033, 0.1612116, 0.1612072, 
    0.1612123, 0.1612008, 0.1611948, 0.1611934, 0.1611905, 0.1611934, 
    0.1611932, 0.161196, 0.1611951, 0.1612018, 0.1611982, 0.1612086, 
    0.1612123, 0.1612232, 0.1612299, 0.1612369, 0.16124, 0.1612409, 0.1612413,
  0.1753678, 0.1753722, 0.1753714, 0.1753749, 0.175373, 0.1753753, 0.1753688, 
    0.1753724, 0.1753701, 0.1753683, 0.1753818, 0.1753751, 0.1753892, 
    0.1753848, 0.175396, 0.1753885, 0.1753976, 0.1753959, 0.1754012, 
    0.1753997, 0.1754065, 0.175402, 0.1754102, 0.1754054, 0.1754061, 
    0.1754018, 0.1753765, 0.1753809, 0.1753762, 0.1753769, 0.1753766, 
    0.175373, 0.1753712, 0.1753676, 0.1753682, 0.1753709, 0.1753772, 
    0.1753751, 0.1753805, 0.1753804, 0.1753864, 0.1753837, 0.1753941, 
    0.1753911, 0.1753998, 0.1753976, 0.1753997, 0.175399, 0.1753997, 
    0.1753964, 0.1753978, 0.175395, 0.1753842, 0.1753873, 0.175378, 
    0.1753724, 0.1753689, 0.1753664, 0.1753667, 0.1753674, 0.1753709, 
    0.1753743, 0.1753769, 0.1753786, 0.1753803, 0.1753854, 0.1753883, 
    0.1753946, 0.1753935, 0.1753954, 0.1753974, 0.1754005, 0.1754, 0.1754014, 
    0.1753954, 0.1753993, 0.1753929, 0.1753946, 0.1753806, 0.1753756, 
    0.1753734, 0.1753716, 0.175367, 0.1753701, 0.1753689, 0.1753719, 
    0.1753738, 0.1753729, 0.1753787, 0.1753764, 0.1753884, 0.1753832, 
    0.1753971, 0.1753938, 0.1753979, 0.1753958, 0.1753995, 0.1753962, 
    0.1754019, 0.1754031, 0.1754023, 0.1754056, 0.175396, 0.1753996, 
    0.1753728, 0.175373, 0.1753737, 0.1753705, 0.1753703, 0.1753675, 
    0.1753701, 0.1753711, 0.1753739, 0.1753755, 0.1753771, 0.1753805, 
    0.1753844, 0.1753899, 0.175394, 0.1753967, 0.175395, 0.1753965, 
    0.1753949, 0.1753941, 0.1754027, 0.1753978, 0.1754051, 0.1754047, 
    0.1754014, 0.1754048, 0.1753731, 0.1753722, 0.1753691, 0.1753715, 
    0.1753672, 0.1753696, 0.175371, 0.1753764, 0.1753777, 0.1753787, 
    0.175381, 0.1753838, 0.1753888, 0.1753933, 0.1753975, 0.1753972, 
    0.1753973, 0.1753982, 0.1753959, 0.1753986, 0.175399, 0.1753978, 
    0.1754047, 0.1754027, 0.1754047, 0.1754035, 0.1753725, 0.175374, 
    0.1753732, 0.1753747, 0.1753736, 0.1753783, 0.1753797, 0.1753865, 
    0.1753837, 0.1753882, 0.1753842, 0.1753849, 0.1753882, 0.1753844, 
    0.175393, 0.1753871, 0.1753982, 0.1753921, 0.1753986, 0.1753975, 
    0.1753994, 0.1754011, 0.1754033, 0.1754073, 0.1754064, 0.1754098, 
    0.1753762, 0.1753781, 0.175378, 0.17538, 0.1753815, 0.1753848, 0.1753901, 
    0.1753881, 0.1753919, 0.1753926, 0.175387, 0.1753904, 0.1753794, 
    0.1753811, 0.1753801, 0.1753763, 0.1753885, 0.1753822, 0.175394, 
    0.1753905, 0.1754008, 0.1753956, 0.1754058, 0.1754102, 0.1754145, 
    0.1754194, 0.1753792, 0.1753779, 0.1753803, 0.1753835, 0.1753866, 
    0.1753908, 0.1753912, 0.175392, 0.175394, 0.1753957, 0.1753922, 
    0.1753962, 0.1753814, 0.1753891, 0.1753773, 0.1753808, 0.1753833, 
    0.1753822, 0.1753879, 0.1753893, 0.1753947, 0.1753919, 0.1754091, 
    0.1754014, 0.1754233, 0.175417, 0.1753774, 0.1753792, 0.1753854, 
    0.1753824, 0.175391, 0.1753932, 0.175395, 0.1753972, 0.1753974, 
    0.1753988, 0.1753966, 0.1753987, 0.1753908, 0.1753943, 0.1753847, 
    0.175387, 0.175386, 0.1753848, 0.1753884, 0.1753922, 0.1753924, 
    0.1753936, 0.1753969, 0.1753911, 0.1754099, 0.1753981, 0.1753812, 
    0.1753845, 0.1753851, 0.1753838, 0.175393, 0.1753896, 0.1753987, 
    0.1753963, 0.1754003, 0.1753983, 0.175398, 0.1753954, 0.1753938, 
    0.1753897, 0.1753865, 0.175384, 0.1753846, 0.1753873, 0.1753924, 
    0.1753974, 0.1753963, 0.1754, 0.1753904, 0.1753944, 0.1753928, 0.1753969, 
    0.1753881, 0.1753954, 0.1753862, 0.175387, 0.1753895, 0.1753946, 
    0.1753958, 0.175397, 0.1753963, 0.1753926, 0.175392, 0.1753895, 
    0.1753887, 0.1753868, 0.1753852, 0.1753867, 0.1753882, 0.1753926, 
    0.1753966, 0.1754011, 0.1754022, 0.1754073, 0.175403, 0.17541, 0.1754039, 
    0.1754145, 0.1753959, 0.1754039, 0.1753897, 0.1753912, 0.1753939, 
    0.1754003, 0.1753969, 0.1754009, 0.175392, 0.1753874, 0.1753863, 
    0.1753841, 0.1753863, 0.1753862, 0.1753883, 0.1753876, 0.1753928, 
    0.17539, 0.175398, 0.1754009, 0.1754094, 0.1754147, 0.1754202, 0.1754226, 
    0.1754234, 0.1754237,
  0.1899663, 0.1899676, 0.1899674, 0.1899685, 0.1899679, 0.1899686, 
    0.1899666, 0.1899677, 0.189967, 0.1899665, 0.1899706, 0.1899685, 
    0.189973, 0.1899715, 0.1899752, 0.1899727, 0.1899758, 0.1899752, 
    0.189977, 0.1899765, 0.1899788, 0.1899772, 0.1899801, 0.1899784, 
    0.1899787, 0.1899772, 0.1899689, 0.1899703, 0.1899689, 0.189969, 
    0.189969, 0.1899679, 0.1899673, 0.1899662, 0.1899664, 0.1899672, 
    0.1899691, 0.1899685, 0.1899702, 0.1899701, 0.1899721, 0.1899712, 
    0.1899746, 0.1899736, 0.1899765, 0.1899757, 0.1899765, 0.1899762, 
    0.1899765, 0.1899754, 0.1899758, 0.1899749, 0.1899713, 0.1899724, 
    0.1899694, 0.1899677, 0.1899666, 0.1899659, 0.189966, 0.1899662, 
    0.1899672, 0.1899683, 0.1899691, 0.1899696, 0.1899701, 0.1899717, 
    0.1899727, 0.1899748, 0.1899744, 0.189975, 0.1899757, 0.1899767, 
    0.1899766, 0.189977, 0.189975, 0.1899763, 0.1899742, 0.1899748, 
    0.1899702, 0.1899687, 0.189968, 0.1899674, 0.1899661, 0.189967, 
    0.1899666, 0.1899675, 0.1899681, 0.1899678, 0.1899696, 0.1899689, 
    0.1899727, 0.189971, 0.1899756, 0.1899745, 0.1899759, 0.1899752, 
    0.1899764, 0.1899753, 0.1899772, 0.1899776, 0.1899773, 0.1899785, 
    0.1899752, 0.1899764, 0.1899678, 0.1899679, 0.1899681, 0.1899671, 
    0.1899671, 0.1899662, 0.189967, 0.1899673, 0.1899681, 0.1899686, 
    0.1899691, 0.1899702, 0.1899714, 0.1899732, 0.1899745, 0.1899755, 
    0.1899749, 0.1899754, 0.1899748, 0.1899746, 0.1899775, 0.1899758, 
    0.1899783, 0.1899782, 0.189977, 0.1899782, 0.1899679, 0.1899676, 
    0.1899667, 0.1899674, 0.1899661, 0.1899668, 0.1899672, 0.1899689, 
    0.1899693, 0.1899696, 0.1899703, 0.1899712, 0.1899728, 0.1899743, 
    0.1899757, 0.1899756, 0.1899756, 0.1899759, 0.1899752, 0.1899761, 
    0.1899762, 0.1899758, 0.1899782, 0.1899775, 0.1899782, 0.1899778, 
    0.1899677, 0.1899682, 0.1899679, 0.1899684, 0.189968, 0.1899695, 
    0.1899699, 0.1899721, 0.1899712, 0.1899726, 0.1899714, 0.1899716, 
    0.1899726, 0.1899714, 0.1899742, 0.1899723, 0.189976, 0.1899739, 
    0.1899761, 0.1899757, 0.1899763, 0.1899769, 0.1899777, 0.1899791, 
    0.1899788, 0.18998, 0.1899688, 0.1899694, 0.1899694, 0.18997, 0.1899705, 
    0.1899716, 0.1899733, 0.1899726, 0.1899738, 0.1899741, 0.1899722, 
    0.1899734, 0.1899698, 0.1899704, 0.1899701, 0.1899689, 0.1899727, 
    0.1899707, 0.1899746, 0.1899734, 0.1899769, 0.1899751, 0.1899786, 
    0.1899801, 0.1899817, 0.1899834, 0.1899698, 0.1899694, 0.1899701, 
    0.1899711, 0.1899721, 0.1899735, 0.1899736, 0.1899739, 0.1899746, 
    0.1899751, 0.1899739, 0.1899753, 0.1899705, 0.1899729, 0.1899692, 
    0.1899703, 0.1899711, 0.1899707, 0.1899725, 0.189973, 0.1899748, 
    0.1899739, 0.1899797, 0.189977, 0.1899849, 0.1899826, 0.1899692, 
    0.1899698, 0.1899717, 0.1899708, 0.1899736, 0.1899743, 0.1899749, 
    0.1899756, 0.1899757, 0.1899762, 0.1899754, 0.1899761, 0.1899735, 
    0.1899747, 0.1899715, 0.1899723, 0.1899719, 0.1899716, 0.1899727, 
    0.189974, 0.189974, 0.1899744, 0.1899755, 0.1899736, 0.18998, 0.1899759, 
    0.1899704, 0.1899714, 0.1899716, 0.1899712, 0.1899742, 0.1899731, 
    0.1899761, 0.1899753, 0.1899767, 0.189976, 0.1899759, 0.189975, 
    0.1899745, 0.1899731, 0.1899721, 0.1899713, 0.1899715, 0.1899724, 
    0.189974, 0.1899757, 0.1899753, 0.1899766, 0.1899734, 0.1899747, 
    0.1899742, 0.1899755, 0.1899726, 0.189975, 0.189972, 0.1899723, 
    0.1899731, 0.1899747, 0.1899752, 0.1899756, 0.1899753, 0.1899741, 
    0.1899739, 0.1899731, 0.1899728, 0.1899722, 0.1899717, 0.1899721, 
    0.1899726, 0.1899741, 0.1899754, 0.1899769, 0.1899773, 0.1899791, 
    0.1899776, 0.18998, 0.1899779, 0.1899817, 0.1899752, 0.1899779, 
    0.1899731, 0.1899736, 0.1899745, 0.1899767, 0.1899755, 0.1899769, 
    0.1899739, 0.1899724, 0.189972, 0.1899713, 0.189972, 0.189972, 0.1899727, 
    0.1899725, 0.1899741, 0.1899732, 0.1899759, 0.1899769, 0.1899798, 
    0.1899817, 0.1899837, 0.1899846, 0.1899849, 0.189985,
  0.1973253, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 
    0.1973252, 0.1973252, 0.1973252, 0.1973253, 0.1973251, 0.1973252, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 0.1973251, 
    0.1973251, 0.1973252, 0.1973252, 0.1973253, 0.1973253, 0.1973252, 
    0.1973251, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973252, 0.1973252, 0.1973253, 0.1973253, 0.1973253, 
    0.1973252, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973252, 0.1973252, 0.1973252, 0.1973253, 0.1973252, 
    0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 
    0.1973252, 0.1973253, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 0.1973252, 
    0.1973252, 0.1973252, 0.1973253, 0.1973252, 0.1973252, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973252, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973252, 0.1973252, 0.1973253, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973254, 0.1973252, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973252, 0.1973251, 0.1973252, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973252, 0.1973252, 0.1973253, 0.1973253, 
    0.1973254, 0.1973254,
  0.1984806, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984806, 0.1984805, 0.1984805, 0.1984806, 0.1984805, 0.1984805, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984803, 0.1984804, 0.1984803, 0.1984803, 
    0.1984803, 0.1984804, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984805, 0.1984806, 0.1984806, 0.1984805, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984804, 0.1984805, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984805, 0.1984804, 
    0.1984805, 0.1984805, 0.1984806, 0.1984806, 0.1984806, 0.1984806, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984806, 0.1984805, 
    0.1984806, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984804, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984803, 
    0.1984804, 0.1984804, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984806, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984803, 0.1984803, 0.1984804, 0.1984803, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984806, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984803, 0.1984804, 0.1984803, 0.1984804, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984804, 0.1984805, 0.1984804, 0.1984805, 0.1984804, 
    0.1984804, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984803, 
    0.1984803, 0.1984803, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984804, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984803, 0.1984803, 0.1984803, 0.1984803, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984805, 0.1984804, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984803, 0.1984804, 0.1984803, 0.1984803, 
    0.1984805, 0.1984805, 0.1984804, 0.1984805, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984803, 0.1984804, 0.1984805, 0.1984805, 0.1984804, 0.1984805, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984805, 
    0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984803, 0.1984804, 0.1984803, 0.1984803, 0.1984803, 
    0.1984804, 0.1984803, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984805, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984803, 0.1984803, 0.1984803, 0.1984803, 
    0.1984803, 0.1984803,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  5.611732, 5.611785, 5.611775, 5.611816, 5.611794, 5.611821, 5.611743, 
    5.611786, 5.611759, 5.611738, 5.611895, 5.611818, 5.611979, 5.61193, 
    5.612058, 5.611971, 5.612076, 5.612057, 5.612118, 5.612101, 5.612175, 
    5.612126, 5.612216, 5.612164, 5.612172, 5.612124, 5.611835, 5.611886, 
    5.611832, 5.611839, 5.611836, 5.611794, 5.611772, 5.611729, 5.611737, 
    5.611769, 5.611843, 5.611818, 5.611881, 5.61188, 5.611948, 5.611917, 
    5.612036, 5.612001, 5.612102, 5.612076, 5.6121, 5.612093, 5.6121, 
    5.612063, 5.612079, 5.612047, 5.611923, 5.611959, 5.611853, 5.611786, 
    5.611745, 5.611715, 5.611719, 5.611727, 5.611769, 5.611809, 5.61184, 
    5.61186, 5.61188, 5.611937, 5.611969, 5.612042, 5.61203, 5.612051, 
    5.612074, 5.61211, 5.612104, 5.612119, 5.612051, 5.612096, 5.612022, 
    5.612042, 5.611881, 5.611825, 5.611798, 5.611777, 5.611722, 5.61176, 
    5.611745, 5.611781, 5.611803, 5.611792, 5.61186, 5.611834, 5.611971, 
    5.611912, 5.612071, 5.612032, 5.612081, 5.612056, 5.612098, 5.612061, 
    5.612125, 5.612139, 5.612129, 5.612167, 5.612058, 5.6121, 5.611792, 
    5.611794, 5.611802, 5.611764, 5.611762, 5.611729, 5.611759, 5.611772, 
    5.611804, 5.611824, 5.611842, 5.611882, 5.611926, 5.611988, 5.612035, 
    5.612066, 5.612047, 5.612064, 5.612045, 5.612036, 5.612134, 5.612079, 
    5.612161, 5.612157, 5.612119, 5.612157, 5.611795, 5.611784, 5.611748, 
    5.611777, 5.611725, 5.611753, 5.61177, 5.611834, 5.611848, 5.611861, 
    5.611887, 5.611919, 5.611976, 5.612027, 5.612075, 5.612072, 5.612073, 
    5.612083, 5.612057, 5.612088, 5.612092, 5.612079, 5.612156, 5.612134, 
    5.612157, 5.612143, 5.611788, 5.611805, 5.611796, 5.611814, 5.611801, 
    5.611856, 5.611872, 5.611949, 5.611918, 5.611968, 5.611924, 5.611931, 
    5.611968, 5.611927, 5.612023, 5.611956, 5.612083, 5.612012, 5.612088, 
    5.612075, 5.612097, 5.612116, 5.612141, 5.612185, 5.612175, 5.612212, 
    5.611831, 5.611853, 5.611852, 5.611876, 5.611893, 5.61193, 5.61199, 
    5.611968, 5.61201, 5.612018, 5.611955, 5.611993, 5.611868, 5.611888, 
    5.611877, 5.611833, 5.611972, 5.6119, 5.612035, 5.611995, 5.612113, 
    5.612054, 5.612169, 5.612216, 5.612263, 5.612314, 5.611866, 5.611851, 
    5.611878, 5.611915, 5.611951, 5.611997, 5.612002, 5.61201, 5.612035, 
    5.612055, 5.612013, 5.61206, 5.611891, 5.611979, 5.611845, 5.611884, 
    5.611913, 5.611901, 5.611966, 5.61198, 5.612043, 5.61201, 5.612204, 
    5.612119, 5.612356, 5.612289, 5.611845, 5.611866, 5.611937, 5.611903, 
    5.612, 5.612025, 5.612046, 5.612072, 5.612075, 5.61209, 5.612065, 
    5.612089, 5.611997, 5.612039, 5.611929, 5.611955, 5.611944, 5.61193, 
    5.611971, 5.612013, 5.612015, 5.61203, 5.612067, 5.612001, 5.612212, 
    5.612081, 5.611889, 5.611927, 5.611934, 5.611918, 5.612023, 5.611984, 
    5.61209, 5.612062, 5.612108, 5.612085, 5.612081, 5.612051, 5.612032, 
    5.611986, 5.611949, 5.611921, 5.611928, 5.611959, 5.612016, 5.612075, 
    5.612062, 5.612104, 5.611993, 5.61204, 5.612021, 5.612069, 5.611967, 
    5.61205, 5.611946, 5.611955, 5.611983, 5.612041, 5.612057, 5.61207, 
    5.612062, 5.612018, 5.612011, 5.611983, 5.611975, 5.611954, 5.611935, 
    5.611952, 5.611969, 5.612019, 5.612066, 5.612116, 5.612129, 5.612184, 
    5.612137, 5.612213, 5.612146, 5.612262, 5.612057, 5.612147, 5.611985, 
    5.612002, 5.612033, 5.612107, 5.612069, 5.612114, 5.612011, 5.611959, 
    5.611947, 5.611922, 5.611948, 5.611946, 5.61197, 5.611962, 5.61202, 
    5.611989, 5.612081, 5.612114, 5.612208, 5.612264, 5.612323, 5.612349, 
    5.612357, 5.61236 ;

 URBAN_AC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 URBAN_HEAT =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 VOCFLXT =
  6.476429e-15, 6.475229e-15, 6.475457e-15, 6.474503e-15, 6.475024e-15, 
    6.474405e-15, 6.476176e-15, 6.475191e-15, 6.475813e-15, 6.476308e-15, 
    6.472684e-15, 6.474457e-15, 6.470752e-15, 6.471895e-15, 6.468998e-15, 
    6.470942e-15, 6.468602e-15, 6.469031e-15, 6.467687e-15, 6.46807e-15, 
    6.466401e-15, 6.46751e-15, 6.465502e-15, 6.466654e-15, 6.466482e-15, 
    6.46755e-15, 6.474079e-15, 6.472911e-15, 6.474153e-15, 6.473985e-15, 
    6.474056e-15, 6.475021e-15, 6.475522e-15, 6.476506e-15, 6.476323e-15, 
    6.475592e-15, 6.473909e-15, 6.474465e-15, 6.473022e-15, 6.473053e-15, 
    6.471464e-15, 6.472181e-15, 6.469498e-15, 6.470255e-15, 6.468054e-15, 
    6.46861e-15, 6.468084e-15, 6.46824e-15, 6.468082e-15, 6.468896e-15, 
    6.468548e-15, 6.469258e-15, 6.472051e-15, 6.471236e-15, 6.473681e-15, 
    6.475188e-15, 6.476137e-15, 6.476827e-15, 6.47673e-15, 6.476548e-15, 
    6.475588e-15, 6.474668e-15, 6.473974e-15, 6.473515e-15, 6.473058e-15, 
    6.471737e-15, 6.47099e-15, 6.469356e-15, 6.469632e-15, 6.469151e-15, 
    6.468664e-15, 6.467874e-15, 6.468001e-15, 6.467658e-15, 6.469149e-15, 
    6.468165e-15, 6.469793e-15, 6.46935e-15, 6.473011e-15, 6.474312e-15, 
    6.474931e-15, 6.475416e-15, 6.476656e-15, 6.475804e-15, 6.476141e-15, 
    6.475323e-15, 6.474813e-15, 6.475062e-15, 6.473502e-15, 6.47411e-15, 
    6.470946e-15, 6.472307e-15, 6.468721e-15, 6.469574e-15, 6.468514e-15, 
    6.469051e-15, 6.468137e-15, 6.468959e-15, 6.467524e-15, 6.467221e-15, 
    6.46743e-15, 6.466603e-15, 6.469007e-15, 6.468091e-15, 6.475072e-15, 
    6.475032e-15, 6.474837e-15, 6.475698e-15, 6.475747e-15, 6.476514e-15, 
    6.475824e-15, 6.475537e-15, 6.474778e-15, 6.474343e-15, 6.473925e-15, 
    6.473007e-15, 6.471995e-15, 6.47056e-15, 6.469519e-15, 6.468826e-15, 
    6.469246e-15, 6.468876e-15, 6.469292e-15, 6.469484e-15, 6.46734e-15, 
    6.468549e-15, 6.466721e-15, 6.46682e-15, 6.467653e-15, 6.466809e-15, 
    6.475003e-15, 6.475236e-15, 6.47607e-15, 6.475417e-15, 6.476597e-15, 
    6.475946e-15, 6.475577e-15, 6.474115e-15, 6.473775e-15, 6.473485e-15, 
    6.472894e-15, 6.472145e-15, 6.470837e-15, 6.469689e-15, 6.468633e-15, 
    6.468709e-15, 6.468683e-15, 6.468455e-15, 6.469029e-15, 6.468359e-15, 
    6.468254e-15, 6.468541e-15, 6.466834e-15, 6.46732e-15, 6.466822e-15, 
    6.467136e-15, 6.475158e-15, 6.474763e-15, 6.474977e-15, 6.474578e-15, 
    6.474865e-15, 6.473609e-15, 6.473232e-15, 6.471453e-15, 6.472164e-15, 
    6.471012e-15, 6.472041e-15, 6.471862e-15, 6.471006e-15, 6.47198e-15, 
    6.469767e-15, 6.471295e-15, 6.468446e-15, 6.469998e-15, 6.46835e-15, 
    6.468637e-15, 6.468154e-15, 6.467731e-15, 6.467184e-15, 6.466199e-15, 
    6.466424e-15, 6.465588e-15, 6.474166e-15, 6.473661e-15, 6.473691e-15, 
    6.473153e-15, 6.472758e-15, 6.471885e-15, 6.470504e-15, 6.471018e-15, 
    6.470058e-15, 6.46987e-15, 6.471321e-15, 6.470444e-15, 6.473312e-15, 
    6.472863e-15, 6.47312e-15, 6.474135e-15, 6.470919e-15, 6.472576e-15, 
    6.469505e-15, 6.470398e-15, 6.467793e-15, 6.469101e-15, 6.466551e-15, 
    6.4655e-15, 6.464448e-15, 6.463297e-15, 6.47337e-15, 6.473714e-15, 
    6.473084e-15, 6.47224e-15, 6.471416e-15, 6.470346e-15, 6.470229e-15, 
    6.470033e-15, 6.469506e-15, 6.469072e-15, 6.469985e-15, 6.468962e-15, 
    6.472787e-15, 6.470769e-15, 6.473858e-15, 6.472946e-15, 6.472283e-15, 
    6.47256e-15, 6.471073e-15, 6.470729e-15, 6.469334e-15, 6.470046e-15, 
    6.465772e-15, 6.467661e-15, 6.462376e-15, 6.463857e-15, 6.473839e-15, 
    6.473364e-15, 6.471737e-15, 6.472508e-15, 6.470267e-15, 6.469722e-15, 
    6.469268e-15, 6.468711e-15, 6.46864e-15, 6.468309e-15, 6.468854e-15, 
    6.468325e-15, 6.470344e-15, 6.469438e-15, 6.471905e-15, 6.471313e-15, 
    6.47158e-15, 6.471885e-15, 6.470947e-15, 6.469973e-15, 6.469929e-15, 
    6.469621e-15, 6.468795e-15, 6.470257e-15, 6.46557e-15, 6.468499e-15, 
    6.472849e-15, 6.471968e-15, 6.471815e-15, 6.472161e-15, 6.469777e-15, 
    6.470644e-15, 6.468314e-15, 6.468937e-15, 6.46791e-15, 6.468422e-15, 
    6.468498e-15, 6.469152e-15, 6.469566e-15, 6.470608e-15, 6.47145e-15, 
    6.472107e-15, 6.471953e-15, 6.47123e-15, 6.469908e-15, 6.468644e-15, 
    6.468924e-15, 6.467988e-15, 6.47043e-15, 6.469416e-15, 6.469815e-15, 
    6.468771e-15, 6.471037e-15, 6.469176e-15, 6.471521e-15, 6.471311e-15, 
    6.47066e-15, 6.469363e-15, 6.469042e-15, 6.468741e-15, 6.468922e-15, 
    6.46987e-15, 6.470016e-15, 6.470671e-15, 6.470863e-15, 6.471355e-15, 
    6.471773e-15, 6.471397e-15, 6.471006e-15, 6.46986e-15, 6.468843e-15, 
    6.467728e-15, 6.467447e-15, 6.466204e-15, 6.467246e-15, 6.465558e-15, 
    6.46704e-15, 6.464454e-15, 6.469034e-15, 6.467039e-15, 6.470623e-15, 
    6.470231e-15, 6.469544e-15, 6.467927e-15, 6.468776e-15, 6.467772e-15, 
    6.470021e-15, 6.471217e-15, 6.471499e-15, 6.472072e-15, 6.471486e-15, 
    6.471532e-15, 6.470974e-15, 6.471152e-15, 6.469822e-15, 6.470536e-15, 
    6.468506e-15, 6.467775e-15, 6.465684e-15, 6.46442e-15, 6.4631e-15, 
    6.462531e-15, 6.462355e-15, 6.462283e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 WF =
  7.122544, 7.149283, 7.144082, 7.16561, 7.153701, 7.167743, 7.127964, 
    7.150341, 7.136054, 7.124956, 7.207006, 7.166563, 7.249272, 7.223327, 
    7.288661, 7.245221, 7.297448, 7.28742, 7.31767, 7.308995, 7.34776, 
    7.321677, 7.367941, 7.341532, 7.345653, 7.320815, 7.174701, 7.201955, 
    7.173086, 7.176967, 7.175229, 7.153944, 7.143112, 7.120512, 7.124614, 
    7.14122, 7.178713, 7.166083, 7.197978, 7.197258, 7.232886, 7.216805, 
    7.276908, 7.259789, 7.309357, 7.296864, 7.308767, 7.305158, 7.308814, 
    7.2905, 7.298341, 7.282247, 7.219811, 7.238111, 7.183631, 7.150853, 
    7.128942, 7.113416, 7.115609, 7.119789, 7.141317, 7.161605, 7.176858, 
    7.187074, 7.197154, 7.227691, 7.243929, 7.280366, 7.273793, 7.284941, 
    7.295623, 7.313566, 7.310613, 7.318523, 7.284657, 7.307146, 7.270048, 
    7.280178, 7.199844, 7.169491, 7.15651, 7.14508, 7.117295, 7.136471, 
    7.128906, 7.146924, 7.158385, 7.152717, 7.187354, 7.17392, 7.244892, 
    7.214255, 7.294376, 7.275143, 7.298994, 7.286819, 7.307687, 7.288904, 
    7.321473, 7.328574, 7.32372, 7.342398, 7.287862, 7.308762, 7.152556, 
    7.15348, 7.157791, 7.138855, 7.1377, 7.120398, 7.135796, 7.142357, 
    7.159054, 7.168809, 7.178069, 7.198462, 7.221282, 7.253304, 7.276388, 
    7.29189, 7.282385, 7.290776, 7.281394, 7.277002, 7.325909, 7.298412, 
    7.339709, 7.337421, 7.318709, 7.337679, 7.15413, 7.148812, 7.130359, 
    7.144797, 7.118516, 7.133212, 7.141669, 7.174189, 7.181296, 7.187876, 
    7.200896, 7.217627, 7.247047, 7.272731, 7.296247, 7.294523, 7.295129, 
    7.300385, 7.287365, 7.302524, 7.305066, 7.298414, 7.337114, 7.326043, 
    7.337372, 7.330163, 7.150541, 7.159494, 7.154655, 7.16371, 7.157339, 
    7.185496, 7.193939, 7.233564, 7.217294, 7.243216, 7.219928, 7.224047, 
    7.244041, 7.221189, 7.271303, 7.237278, 7.300589, 7.266483, 7.302729, 
    7.296145, 7.307054, 7.31683, 7.329152, 7.351915, 7.346642, 7.365717, 
    7.172675, 7.18413, 7.183131, 7.19514, 7.20403, 7.22334, 7.254385, 
    7.242702, 7.264173, 7.268486, 7.235877, 7.255875, 7.191813, 7.202122, 
    7.19599, 7.173573, 7.245379, 7.208451, 7.276768, 7.256678, 7.315434, 
    7.286158, 7.343737, 7.368434, 7.39178, 7.419083, 7.190399, 7.182607, 
    7.196572, 7.215911, 7.23392, 7.2579, 7.260363, 7.26486, 7.276533, 
    7.286354, 7.266273, 7.288818, 7.204496, 7.248596, 7.179654, 7.200346, 
    7.214775, 7.208452, 7.24137, 7.249142, 7.280789, 7.264421, 7.362324, 
    7.318882, 7.439955, 7.405961, 7.179884, 7.190377, 7.226976, 7.209546, 
    7.259508, 7.271844, 7.281893, 7.294738, 7.296133, 7.303754, 7.291267, 
    7.303264, 7.257951, 7.278175, 7.222797, 7.236239, 7.230056, 7.223272, 
    7.244226, 7.266587, 7.267081, 7.27426, 7.294493, 7.259712, 7.367917, 
    7.300918, 7.201832, 7.222081, 7.224996, 7.217141, 7.270606, 7.251196, 
    7.30357, 7.28939, 7.31264, 7.301078, 7.299377, 7.284554, 7.275334, 
    7.252082, 7.233211, 7.218282, 7.221752, 7.238159, 7.26796, 7.296252, 
    7.290045, 7.310871, 7.255876, 7.278889, 7.269983, 7.293226, 7.242388, 
    7.285615, 7.231366, 7.236113, 7.250811, 7.280441, 7.287033, 7.294047, 
    7.289721, 7.268721, 7.265292, 7.250457, 7.246358, 7.23508, 7.225747, 
    7.23427, 7.243227, 7.268736, 7.291776, 7.316967, 7.323148, 7.352646, 
    7.328605, 7.368288, 7.334507, 7.393075, 7.288149, 7.333547, 7.251486, 
    7.260295, 7.276235, 7.312928, 7.293117, 7.316298, 7.265159, 7.238718, 
    7.231908, 7.219186, 7.2322, 7.231141, 7.243609, 7.239602, 7.269585, 
    7.253468, 7.29933, 7.316119, 7.363711, 7.392994, 7.422918, 7.43615, 
    7.440183, 7.441868 ;

 WIND =
  5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932 ;

 WOODC =
  0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  0.0002000768, 0.0002000343, 0.0002000423, 0.0002000088, 0.0002000271, 
    0.0002000054, 0.0002000678, 0.0002000329, 0.0002000549, 0.0002000725, 
    0.0001999457, 0.0002000073, 0.0001998799, 0.0001999189, 0.0001998204, 
    0.0001998863, 0.000199807, 0.0001998216, 0.0001997761, 0.0001997891, 
    0.0001997326, 0.0001997701, 0.0001997023, 0.0001997412, 0.0001997353, 
    0.0001997715, 0.0001999941, 0.0001999536, 0.0001999967, 0.0001999909, 
    0.0001999933, 0.0002000269, 0.0002000445, 0.0002000796, 0.000200073, 
    0.000200047, 0.0001999882, 0.0002000076, 0.0001999576, 0.0001999587, 
    0.0001999042, 0.0001999287, 0.0001998374, 0.0001998631, 0.0001997885, 
    0.0001998073, 0.0001997895, 0.0001997948, 0.0001997894, 0.000199817, 
    0.0001998052, 0.0001998293, 0.0001999243, 0.0001998964, 0.0001999803, 
    0.0002000327, 0.0002000663, 0.0002000911, 0.0002000876, 0.000200081, 
    0.0002000469, 0.0002000146, 0.0001999906, 0.0001999746, 0.0001999589, 
    0.0001999134, 0.000199888, 0.0001998325, 0.0001998419, 0.0001998256, 
    0.0001998091, 0.0001997824, 0.0001997867, 0.0001997751, 0.0001998256, 
    0.0001997922, 0.0001998474, 0.0001998324, 0.000199957, 0.0002000022, 
    0.0002000237, 0.0002000408, 0.0002000849, 0.0002000545, 0.0002000665, 
    0.0002000376, 0.0002000197, 0.0002000284, 0.0001999742, 0.0001999953, 
    0.0001998865, 0.000199933, 0.0001998111, 0.00019984, 0.0001998041, 
    0.0001998223, 0.0001997913, 0.0001998191, 0.0001997706, 0.0001997603, 
    0.0001997674, 0.0001997395, 0.0001998208, 0.0001997897, 0.0002000288, 
    0.0002000274, 0.0002000205, 0.0002000508, 0.0002000525, 0.0002000799, 
    0.0002000553, 0.0002000451, 0.0002000185, 0.0002000033, 0.0001999888, 
    0.0001999571, 0.0001999223, 0.0001998734, 0.0001998381, 0.0001998146, 
    0.0001998289, 0.0001998163, 0.0001998305, 0.000199837, 0.0001997643, 
    0.0001998052, 0.0001997435, 0.0001997468, 0.0001997749, 0.0001997464, 
    0.0002000263, 0.0002000345, 0.000200064, 0.0002000409, 0.0002000829, 
    0.0002000596, 0.0002000465, 0.0001999953, 0.0001999836, 0.0001999736, 
    0.0001999532, 0.0001999275, 0.0001998828, 0.0001998439, 0.0001998081, 
    0.0001998107, 0.0001998098, 0.0001998021, 0.0001998215, 0.0001997988, 
    0.0001997953, 0.000199805, 0.0001997473, 0.0001997637, 0.0001997469, 
    0.0001997575, 0.0002000318, 0.000200018, 0.0002000255, 0.0002000115, 
    0.0002000215, 0.0001999778, 0.0001999648, 0.0001999038, 0.0001999281, 
    0.0001998888, 0.0001999239, 0.0001999178, 0.0001998885, 0.0001999219, 
    0.0001998464, 0.0001998984, 0.0001998018, 0.0001998542, 0.0001997985, 
    0.0001998083, 0.0001997919, 0.0001997776, 0.0001997591, 0.0001997258, 
    0.0001997334, 0.0001997052, 0.0001999972, 0.0001999796, 0.0001999807, 
    0.0001999621, 0.0001999485, 0.0001999186, 0.0001998715, 0.000199889, 
    0.0001998564, 0.00019985, 0.0001998994, 0.0001998694, 0.0001999676, 
    0.0001999521, 0.000199961, 0.0001999961, 0.0001998856, 0.0001999422, 
    0.0001998376, 0.0001998679, 0.0001997797, 0.0001998239, 0.0001997377, 
    0.0001997022, 0.0001996668, 0.0001996279, 0.0001999696, 0.0001999815, 
    0.0001999598, 0.0001999307, 0.0001999026, 0.0001998661, 0.0001998622, 
    0.0001998555, 0.0001998377, 0.000199823, 0.0001998538, 0.0001998192, 
    0.0001999494, 0.0001998805, 0.0001999865, 0.0001999549, 0.0001999322, 
    0.0001999417, 0.0001998909, 0.0001998792, 0.0001998318, 0.000199856, 
    0.0001997113, 0.0001997752, 0.0001995969, 0.0001996468, 0.0001999858, 
    0.0001999694, 0.0001999135, 0.00019994, 0.0001998635, 0.000199845, 
    0.0001998296, 0.0001998107, 0.0001998083, 0.0001997971, 0.0001998156, 
    0.0001997977, 0.0001998661, 0.0001998354, 0.0001999193, 0.0001998991, 
    0.0001999082, 0.0001999186, 0.0001998867, 0.0001998535, 0.000199852, 
    0.0001998416, 0.0001998133, 0.0001998632, 0.0001997044, 0.0001998034, 
    0.0001999517, 0.0001999214, 0.0001999162, 0.0001999281, 0.0001998469, 
    0.0001998763, 0.0001997973, 0.0001998184, 0.0001997836, 0.000199801, 
    0.0001998035, 0.0001998257, 0.0001998397, 0.0001998751, 0.0001999037, 
    0.0001999262, 0.0001999209, 0.0001998963, 0.0001998513, 0.0001998084, 
    0.0001998179, 0.0001997863, 0.000199869, 0.0001998346, 0.0001998481, 
    0.0001998128, 0.0001998897, 0.0001998263, 0.0001999062, 0.000199899, 
    0.0001998768, 0.0001998327, 0.000199822, 0.0001998117, 0.0001998179, 
    0.00019985, 0.000199855, 0.0001998772, 0.0001998837, 0.0001999005, 
    0.0001999148, 0.0001999019, 0.0001998886, 0.0001998497, 0.0001998152, 
    0.0001997775, 0.000199768, 0.0001997259, 0.0001997611, 0.000199704, 
    0.000199754, 0.0001996668, 0.0001998216, 0.000199754, 0.0001998756, 
    0.0001998622, 0.0001998389, 0.0001997841, 0.0001998129, 0.0001997789, 
    0.0001998551, 0.0001998958, 0.0001999054, 0.000199925, 0.000199905, 
    0.0001999066, 0.0001998875, 0.0001998936, 0.0001998484, 0.0001998726, 
    0.0001998038, 0.000199779, 0.0001997084, 0.0001996658, 0.0001996214, 
    0.0001996022, 0.0001995963, 0.0001995939 ;

 W_SCALAR =
  0.626114, 0.6277712, 0.6274492, 0.6287847, 0.6280439, 0.6289183, 0.62645, 
    0.627837, 0.6269517, 0.6262631, 0.631373, 0.6288443, 0.6339937, 0.632385, 
    0.6364222, 0.6337437, 0.6369616, 0.6363448, 0.6381996, 0.6376686, 
    0.6400383, 0.6384447, 0.6412646, 0.6396578, 0.6399094, 0.6383921, 
    0.6293533, 0.6310586, 0.6292523, 0.6294956, 0.6293864, 0.6280593, 
    0.6273901, 0.6259871, 0.6262419, 0.6272722, 0.629605, 0.6288134, 
    0.630807, 0.630762, 0.632978, 0.6319793, 0.6356981, 0.6346422, 0.6376907, 
    0.6369248, 0.6376548, 0.6374335, 0.6376576, 0.6365342, 0.6370156, 
    0.6360265, 0.6321665, 0.6333022, 0.6299121, 0.6278697, 0.6265109, 
    0.625546, 0.6256825, 0.6259426, 0.6272783, 0.6285328, 0.629488, 
    0.6301267, 0.6307555, 0.6326579, 0.6336632, 0.6359116, 0.6355059, 
    0.6361929, 0.6368486, 0.6379488, 0.6377677, 0.6382523, 0.6361746, 
    0.6375559, 0.6352749, 0.6358992, 0.6309272, 0.629027, 0.6282191, 
    0.6275111, 0.6257874, 0.626978, 0.6265088, 0.6276246, 0.6283333, 
    0.6279829, 0.6301441, 0.6293043, 0.6337228, 0.6318215, 0.6367721, 
    0.6355892, 0.6370555, 0.6363074, 0.6375889, 0.6364356, 0.6384325, 
    0.638867, 0.6385701, 0.6397099, 0.6363717, 0.6376548, 0.627973, 
    0.6280302, 0.6282964, 0.6271258, 0.6270541, 0.6259801, 0.6269357, 
    0.6273425, 0.6283743, 0.6289844, 0.629564, 0.6308375, 0.6322584, 
    0.6342425, 0.6356659, 0.6366192, 0.6360347, 0.6365507, 0.6359739, 
    0.6357034, 0.6387042, 0.6370202, 0.639546, 0.6394063, 0.6382638, 
    0.6394221, 0.6280704, 0.6277413, 0.6265987, 0.627493, 0.6258631, 
    0.6267758, 0.6273003, 0.629322, 0.6297656, 0.630177, 0.630989, 0.6320305, 
    0.6338555, 0.6354411, 0.6368867, 0.6367808, 0.6368181, 0.6371409, 
    0.6363412, 0.6372721, 0.6374283, 0.6370199, 0.6393877, 0.6387116, 
    0.6394034, 0.6389633, 0.6278483, 0.6284018, 0.6281027, 0.628665, 
    0.628269, 0.6300293, 0.6305566, 0.6330211, 0.63201, 0.6336185, 0.6321735, 
    0.6324297, 0.6336712, 0.6322516, 0.6353538, 0.6332517, 0.6371534, 
    0.6350575, 0.6372846, 0.6368804, 0.6375495, 0.6381486, 0.6389017, 
    0.6402902, 0.6399688, 0.641129, 0.6292263, 0.6299434, 0.6298802, 
    0.6306302, 0.6311846, 0.6323853, 0.6343088, 0.6335858, 0.6349127, 
    0.635179, 0.6331629, 0.6344012, 0.6304231, 0.6310667, 0.6306834, 
    0.629283, 0.6337526, 0.6314608, 0.6356894, 0.6344503, 0.6380632, 
    0.6362679, 0.6397918, 0.6412956, 0.6427084, 0.644358, 0.6303345, 
    0.6298475, 0.6307193, 0.6319249, 0.633042, 0.6345259, 0.6346776, 
    0.6349554, 0.6356745, 0.6362789, 0.6350433, 0.6364304, 0.6312163, 
    0.6339513, 0.6296633, 0.6309562, 0.6318538, 0.63146, 0.6335031, 
    0.6339842, 0.6359374, 0.634928, 0.6409247, 0.6382753, 0.645612, 
    0.6435664, 0.6296772, 0.6303328, 0.6326118, 0.6315279, 0.6346248, 
    0.635386, 0.6360044, 0.6367946, 0.6368797, 0.6373476, 0.6365809, 
    0.6373174, 0.6345291, 0.6357759, 0.6323513, 0.6331858, 0.6328019, 
    0.6323808, 0.63368, 0.6350628, 0.6350921, 0.6355352, 0.6367835, 
    0.6346374, 0.6412666, 0.6371772, 0.6310472, 0.6323085, 0.6324883, 0.632, 
    0.6353098, 0.6341115, 0.6373363, 0.6364655, 0.6378918, 0.6371832, 
    0.637079, 0.6361682, 0.635601, 0.6341665, 0.6329982, 0.6320708, 
    0.6322864, 0.633305, 0.6351473, 0.6368876, 0.6365066, 0.6377835, 
    0.6344005, 0.6358203, 0.6352718, 0.6367014, 0.6335666, 0.6362373, 
    0.6328831, 0.6331775, 0.6340877, 0.6359167, 0.6363207, 0.6367522, 
    0.6364859, 0.635194, 0.6349822, 0.6340656, 0.6338125, 0.6331134, 
    0.6325345, 0.6330635, 0.6336189, 0.6351945, 0.6366128, 0.6381571, 
    0.6385347, 0.6403366, 0.6388703, 0.6412894, 0.6392335, 0.64279, 
    0.6363915, 0.6391725, 0.634129, 0.6346734, 0.6356574, 0.6379111, 
    0.6366947, 0.638117, 0.6349738, 0.6333402, 0.6329169, 0.6321272, 
    0.6329349, 0.6328692, 0.6336417, 0.6333935, 0.6352468, 0.6342516, 
    0.6370764, 0.6381058, 0.6410075, 0.642783, 0.6445873, 0.6453831, 
    0.6456251, 0.6457263,
  0.5467896, 0.5488337, 0.5484365, 0.5500841, 0.5491702, 0.5502488, 
    0.5472041, 0.5489149, 0.5478229, 0.5469736, 0.5532776, 0.5501575, 
    0.5565122, 0.5545264, 0.5595103, 0.5562034, 0.5601763, 0.5594147, 
    0.5617052, 0.5610493, 0.5639763, 0.5620078, 0.5654912, 0.5635062, 
    0.563817, 0.5619429, 0.5507856, 0.5528895, 0.5506609, 0.5509611, 
    0.5508264, 0.5491892, 0.5483637, 0.5466332, 0.5469474, 0.5482183, 
    0.551096, 0.5501195, 0.5525792, 0.5525237, 0.5552585, 0.5540259, 
    0.5586162, 0.5573127, 0.5610767, 0.5601309, 0.5610324, 0.560759, 
    0.5610359, 0.5596485, 0.5602431, 0.5590217, 0.5542569, 0.5556586, 
    0.5514749, 0.5489553, 0.5472792, 0.5460892, 0.5462575, 0.5465783, 
    0.5482258, 0.5497732, 0.5509517, 0.5517396, 0.5525157, 0.5548633, 
    0.5561041, 0.5588798, 0.558379, 0.5592272, 0.5600367, 0.5613955, 
    0.5611718, 0.5617703, 0.5592046, 0.5609102, 0.5580937, 0.5588645, 
    0.5527274, 0.550383, 0.5493863, 0.5485129, 0.5463869, 0.5478554, 
    0.5472766, 0.548653, 0.5495272, 0.5490948, 0.5517612, 0.550725, 
    0.5561776, 0.553831, 0.5599423, 0.5584818, 0.5602922, 0.5593686, 
    0.5609509, 0.5595269, 0.5619928, 0.5625294, 0.5621628, 0.5635706, 
    0.5594479, 0.5610324, 0.5490828, 0.5491533, 0.5494817, 0.5480376, 
    0.5479492, 0.5466246, 0.5478032, 0.548305, 0.5495778, 0.5503303, 
    0.5510455, 0.5526168, 0.5543703, 0.5568193, 0.5585765, 0.5597535, 
    0.5590318, 0.559669, 0.5589567, 0.5586227, 0.5623285, 0.5602487, 
    0.5633681, 0.5631956, 0.5617845, 0.5632151, 0.5492028, 0.548797, 
    0.5473875, 0.5484906, 0.5464803, 0.5476059, 0.5482529, 0.5507469, 
    0.5512942, 0.5518018, 0.5528038, 0.554089, 0.5563414, 0.5582989, 
    0.5600838, 0.5599531, 0.5599991, 0.5603977, 0.5594103, 0.5605597, 
    0.5607526, 0.5602483, 0.5631725, 0.5623376, 0.563192, 0.5626484, 
    0.5489289, 0.5496116, 0.5492427, 0.5499364, 0.5494478, 0.5516195, 
    0.5522702, 0.5553115, 0.5540637, 0.556049, 0.5542654, 0.5545816, 
    0.556114, 0.5543618, 0.5581912, 0.5555962, 0.5604132, 0.5578253, 
    0.5605752, 0.5600761, 0.5609024, 0.5616422, 0.5625723, 0.5642874, 
    0.5638904, 0.5653237, 0.5506288, 0.5515136, 0.5514356, 0.552361, 
    0.5530451, 0.5545269, 0.5569011, 0.5560086, 0.5576466, 0.5579753, 
    0.5554866, 0.5570152, 0.5521054, 0.5528997, 0.5524267, 0.5506988, 
    0.5562145, 0.5533859, 0.5586056, 0.5570757, 0.5615367, 0.5593197, 
    0.5636718, 0.5655294, 0.567275, 0.5693137, 0.5519961, 0.5513952, 
    0.5524709, 0.5539586, 0.5553374, 0.5571691, 0.5573564, 0.5576993, 
    0.5585871, 0.5593334, 0.5578079, 0.5595204, 0.5530841, 0.5564598, 
    0.5511681, 0.5527633, 0.5538709, 0.553385, 0.5559065, 0.5565004, 
    0.5589117, 0.5576655, 0.5650712, 0.5617986, 0.5708637, 0.5683354, 
    0.5511852, 0.551994, 0.5548064, 0.5534688, 0.5572913, 0.558231, 
    0.5589944, 0.5599701, 0.5600753, 0.5606531, 0.5597062, 0.5606156, 
    0.557173, 0.5587122, 0.554485, 0.5555149, 0.5550411, 0.5545214, 
    0.5561249, 0.5578319, 0.5578681, 0.5584152, 0.5599563, 0.5573067, 
    0.5654936, 0.5604425, 0.5528756, 0.5544321, 0.554654, 0.5540513, 
    0.5581368, 0.5566576, 0.560639, 0.5595638, 0.5613251, 0.5604501, 
    0.5603213, 0.5591968, 0.5584964, 0.5567254, 0.5552832, 0.5541387, 
    0.5544049, 0.5556619, 0.5579363, 0.5600849, 0.5596145, 0.5611913, 
    0.5570143, 0.5587671, 0.55809, 0.559855, 0.5559849, 0.5592818, 0.5551413, 
    0.5555047, 0.5566282, 0.5588861, 0.5593849, 0.5599178, 0.559589, 
    0.5579939, 0.5577323, 0.5566008, 0.5562884, 0.5554256, 0.554711, 
    0.555364, 0.5560495, 0.5579945, 0.5597456, 0.5616527, 0.5621191, 
    0.5643448, 0.5625335, 0.5655218, 0.562982, 0.5673758, 0.5594723, 
    0.5629068, 0.5566792, 0.5573511, 0.558566, 0.5613488, 0.5598468, 
    0.5616032, 0.557722, 0.5557054, 0.555183, 0.5542084, 0.5552053, 
    0.5551242, 0.5560777, 0.5557713, 0.558059, 0.5568305, 0.5603182, 
    0.5615892, 0.5651736, 0.5673673, 0.5695971, 0.5705807, 0.57088, 0.571005,
  0.514181, 0.516431, 0.5159937, 0.5178076, 0.5168014, 0.517989, 0.5146372, 
    0.5165204, 0.5153183, 0.5143835, 0.5213248, 0.5178885, 0.5248888, 
    0.5227006, 0.5281937, 0.5245485, 0.528928, 0.5280883, 0.5306142, 
    0.5298908, 0.5331194, 0.530948, 0.5347911, 0.5326009, 0.5329437, 
    0.5308763, 0.5185801, 0.5208973, 0.5184428, 0.5187734, 0.518625, 
    0.5168223, 0.5159136, 0.5140088, 0.5143547, 0.5157536, 0.518922, 
    0.5178466, 0.5205554, 0.5204943, 0.5235071, 0.5221491, 0.527208, 
    0.525771, 0.529921, 0.528878, 0.5298721, 0.5295706, 0.529876, 0.5283461, 
    0.5290017, 0.527655, 0.5224035, 0.523948, 0.5193393, 0.5165648, 
    0.5147199, 0.5134102, 0.5135954, 0.5139484, 0.5157617, 0.5174654, 
    0.5187631, 0.5196308, 0.5204855, 0.5230717, 0.524439, 0.5274985, 
    0.5269464, 0.5278815, 0.5287742, 0.5302725, 0.530026, 0.5306859, 
    0.5278566, 0.5297374, 0.526632, 0.5274817, 0.5207186, 0.5181367, 
    0.5170394, 0.5160778, 0.5137378, 0.515354, 0.514717, 0.5162321, 
    0.5171944, 0.5167184, 0.5196545, 0.5185134, 0.52452, 0.5219344, 
    0.5286701, 0.5270597, 0.5290559, 0.5280374, 0.5297823, 0.528212, 
    0.5309314, 0.5315233, 0.5311189, 0.5326718, 0.5281249, 0.5298721, 
    0.5167052, 0.5167828, 0.5171444, 0.5155546, 0.5154573, 0.5139994, 
    0.5152966, 0.5158489, 0.5172502, 0.5180788, 0.5188663, 0.5205969, 
    0.5225285, 0.5252272, 0.5271642, 0.5284618, 0.5276662, 0.5283687, 
    0.5275834, 0.5272152, 0.5313016, 0.5290079, 0.5324485, 0.5322582, 
    0.5307016, 0.5322797, 0.5168373, 0.5163905, 0.5148391, 0.5160533, 
    0.5138406, 0.5150794, 0.5157917, 0.5185375, 0.5191402, 0.5196993, 
    0.5208029, 0.5222186, 0.5247006, 0.5268581, 0.5288261, 0.5286819, 
    0.5287327, 0.5291722, 0.5280834, 0.5293509, 0.5295636, 0.5290075, 
    0.5322328, 0.5313117, 0.5322542, 0.5316545, 0.5165358, 0.5172874, 
    0.5168813, 0.5176449, 0.517107, 0.5194985, 0.5202151, 0.5235656, 
    0.5221908, 0.5243783, 0.522413, 0.5227614, 0.5244499, 0.5225192, 
    0.5267394, 0.5238793, 0.5291893, 0.5263361, 0.529368, 0.5288175, 
    0.5297288, 0.5305446, 0.5315706, 0.5334628, 0.5330247, 0.5346062, 
    0.5184075, 0.5193818, 0.5192959, 0.5203151, 0.5210686, 0.5227011, 
    0.5253174, 0.5243338, 0.5261391, 0.5265014, 0.5237585, 0.5254431, 
    0.5200336, 0.5209085, 0.5203875, 0.5184845, 0.5245607, 0.5214441, 
    0.5271962, 0.5255099, 0.5304283, 0.5279836, 0.5327836, 0.5348333, 
    0.53676, 0.5390108, 0.5199133, 0.5192514, 0.5204362, 0.522075, 0.5235941, 
    0.5256128, 0.5258191, 0.5261972, 0.5271759, 0.5279986, 0.5263168, 
    0.5282048, 0.5211116, 0.524831, 0.5190013, 0.5207582, 0.5219783, 
    0.521443, 0.5242213, 0.5248758, 0.5275337, 0.5261599, 0.5343276, 
    0.5307172, 0.5407226, 0.5379306, 0.5190201, 0.5199109, 0.5230091, 
    0.5215353, 0.5257474, 0.5267833, 0.5276249, 0.5287007, 0.5288167, 
    0.5294538, 0.5284097, 0.5294125, 0.5256171, 0.5273138, 0.522655, 
    0.5237897, 0.5232677, 0.5226951, 0.5244619, 0.5263433, 0.5263833, 
    0.5269864, 0.5286854, 0.5257645, 0.5347937, 0.5292216, 0.5208819, 
    0.5225966, 0.5228412, 0.5221772, 0.5266795, 0.525049, 0.5294383, 
    0.5282527, 0.5301949, 0.5292299, 0.529088, 0.527848, 0.5270758, 
    0.5251238, 0.5235345, 0.5222734, 0.5225667, 0.5239518, 0.5264584, 
    0.5288273, 0.5283086, 0.5300474, 0.5254422, 0.5273743, 0.5266278, 
    0.5285739, 0.5243077, 0.5279418, 0.5233781, 0.5237785, 0.5250166, 
    0.5275055, 0.5280554, 0.528643, 0.5282804, 0.5265219, 0.5262336, 
    0.5249864, 0.5246422, 0.5236913, 0.522904, 0.5236234, 0.5243788, 
    0.5265225, 0.5284531, 0.5305563, 0.5310706, 0.533526, 0.5315278, 
    0.5348248, 0.5320225, 0.5368713, 0.5281518, 0.5319395, 0.5250729, 
    0.5258134, 0.5271526, 0.5302211, 0.5285647, 0.5305016, 0.5262223, 
    0.5239997, 0.523424, 0.5223501, 0.5234485, 0.5233592, 0.5244099, 
    0.5240723, 0.5265937, 0.5252396, 0.5290845, 0.5304863, 0.5344406, 
    0.5368619, 0.5393238, 0.54041, 0.5407405, 0.5408787,
  0.507081, 0.5094717, 0.5090069, 0.5109348, 0.5098653, 0.5111277, 0.5075657, 
    0.5095666, 0.5082893, 0.5072961, 0.5146752, 0.5110208, 0.5184684, 
    0.5161392, 0.5219887, 0.5181062, 0.5227712, 0.5218765, 0.5245687, 
    0.5237975, 0.5272405, 0.5249246, 0.5290242, 0.5266873, 0.5270531, 
    0.5248482, 0.5117561, 0.5142204, 0.5116101, 0.5119616, 0.5118038, 
    0.5098875, 0.5089218, 0.5068982, 0.5072655, 0.5087517, 0.5121196, 
    0.5109763, 0.5138568, 0.5137918, 0.5169976, 0.5155523, 0.5209385, 
    0.5194079, 0.5238296, 0.522718, 0.5237775, 0.5234562, 0.5237817, 
    0.5221511, 0.5228498, 0.5214148, 0.5158231, 0.5174669, 0.5125633, 
    0.5096138, 0.5076535, 0.5062624, 0.5064591, 0.506834, 0.5087604, 
    0.510571, 0.5119506, 0.5128734, 0.5137824, 0.5165341, 0.5179896, 
    0.521248, 0.5206599, 0.5216561, 0.5226073, 0.5242044, 0.5239415, 
    0.5246451, 0.5216296, 0.523634, 0.5203249, 0.5212302, 0.5140304, 
    0.5112847, 0.5101182, 0.5090963, 0.5066103, 0.5083272, 0.5076504, 
    0.5092602, 0.5102831, 0.5097771, 0.5128986, 0.5116852, 0.5180759, 
    0.5153238, 0.5224963, 0.5207806, 0.5229076, 0.5218222, 0.5236818, 
    0.5220082, 0.5249069, 0.525538, 0.5251068, 0.526763, 0.5219154, 
    0.5237775, 0.509763, 0.5098455, 0.5102298, 0.5085403, 0.5084369, 
    0.5068881, 0.5082662, 0.508853, 0.5103422, 0.5112231, 0.5120604, 
    0.5139009, 0.5159561, 0.5188288, 0.5208918, 0.5222744, 0.5214266, 
    0.5221751, 0.5213384, 0.5209461, 0.5253016, 0.5228564, 0.5265248, 
    0.5263218, 0.5246619, 0.5263447, 0.5099034, 0.5094286, 0.5077801, 
    0.5090702, 0.5067194, 0.5080355, 0.5087922, 0.5117108, 0.5123517, 
    0.5129462, 0.51412, 0.5156263, 0.5182681, 0.5205658, 0.5226626, 0.522509, 
    0.5225631, 0.5230315, 0.5218713, 0.523222, 0.5234487, 0.5228559, 
    0.5262946, 0.5253124, 0.5263175, 0.525678, 0.5095829, 0.5103818, 
    0.5099502, 0.5107619, 0.5101901, 0.5127326, 0.5134948, 0.5170599, 
    0.5155967, 0.517925, 0.5158332, 0.5162039, 0.5180013, 0.5159461, 
    0.5204393, 0.5173937, 0.5230497, 0.5200098, 0.5232402, 0.5226535, 
    0.5236247, 0.5244945, 0.5255885, 0.5276068, 0.5271394, 0.5288268, 
    0.5115726, 0.5126086, 0.5125172, 0.5136012, 0.5144027, 0.5161397, 
    0.5189249, 0.5178776, 0.5197999, 0.5201859, 0.5172652, 0.5190588, 
    0.5133017, 0.5142323, 0.5136781, 0.5116544, 0.5181192, 0.5148022, 
    0.5209259, 0.5191298, 0.5243706, 0.5217649, 0.5268822, 0.5290691, 
    0.531126, 0.5335299, 0.5131738, 0.5124699, 0.51373, 0.5154734, 0.5170902, 
    0.5192394, 0.5194592, 0.5198618, 0.5209044, 0.5217809, 0.5199893, 
    0.5220006, 0.5144485, 0.5184069, 0.5122039, 0.5140725, 0.5153706, 
    0.514801, 0.5177578, 0.5184546, 0.5212855, 0.5198221, 0.5285296, 
    0.5246785, 0.5353591, 0.5323761, 0.512224, 0.5131713, 0.5164675, 
    0.5148993, 0.5193828, 0.5204861, 0.5213827, 0.522529, 0.5226526, 
    0.5233316, 0.5222189, 0.5232877, 0.519244, 0.5210513, 0.5160906, 
    0.5172983, 0.5167427, 0.5161333, 0.518014, 0.5200175, 0.5200601, 
    0.5207024, 0.5225127, 0.519401, 0.529027, 0.5230841, 0.5142041, 
    0.5160285, 0.5162888, 0.5155821, 0.5203755, 0.5186391, 0.5233151, 
    0.5220516, 0.5241216, 0.523093, 0.5229418, 0.5216204, 0.5207977, 
    0.5187187, 0.5170267, 0.5156846, 0.5159967, 0.5174709, 0.52014, 0.522664, 
    0.5221112, 0.5239643, 0.5190578, 0.5211157, 0.5203205, 0.5223938, 
    0.5178498, 0.5217203, 0.5168603, 0.5172865, 0.5186046, 0.5212555, 
    0.5218414, 0.5224675, 0.5220811, 0.5202077, 0.5199006, 0.5185725, 
    0.5182059, 0.5171937, 0.5163556, 0.5171214, 0.5179255, 0.5202084, 
    0.5222652, 0.5245069, 0.5250553, 0.5276743, 0.5255428, 0.5290601, 
    0.5260704, 0.5312447, 0.5219441, 0.5259819, 0.5186645, 0.519453, 
    0.5208795, 0.5241495, 0.522384, 0.5244486, 0.5198885, 0.5175219, 
    0.5169091, 0.5157663, 0.5169352, 0.5168402, 0.5179586, 0.5175992, 
    0.5202841, 0.518842, 0.522938, 0.5244322, 0.5286501, 0.5312347, 
    0.5338643, 0.5350251, 0.5353783, 0.535526,
  0.5310283, 0.5334976, 0.5330174, 0.5350101, 0.5339045, 0.5352095, 
    0.5315287, 0.5335958, 0.532276, 0.5312504, 0.5388804, 0.535099, 0.542811, 
    0.5403967, 0.5464641, 0.5424354, 0.5472769, 0.5463476, 0.5491447, 
    0.5483431, 0.5519236, 0.5495147, 0.5537806, 0.551348, 0.5517285, 
    0.5494353, 0.5358595, 0.5384095, 0.5357085, 0.536072, 0.5359088, 
    0.5339274, 0.5329295, 0.5308394, 0.5312188, 0.5327538, 0.5362355, 
    0.5350531, 0.5380331, 0.5379658, 0.5412862, 0.5397888, 0.5453737, 
    0.5437855, 0.5483766, 0.5472215, 0.5483223, 0.5479885, 0.5483267, 
    0.5466328, 0.5473585, 0.5458682, 0.5400692, 0.5417727, 0.5366945, 
    0.5336446, 0.5316194, 0.5301831, 0.5303861, 0.5307732, 0.5327628, 
    0.534634, 0.5360606, 0.5370153, 0.5379561, 0.5408059, 0.5423146, 
    0.5456951, 0.5450845, 0.5461187, 0.5471066, 0.548766, 0.5484928, 
    0.5492241, 0.5460913, 0.5481732, 0.5447369, 0.5456765, 0.5382128, 
    0.535372, 0.5341659, 0.5331097, 0.5305423, 0.5323152, 0.5316162, 
    0.5332791, 0.5343363, 0.5338134, 0.5370414, 0.5357862, 0.542404, 
    0.5395521, 0.5469913, 0.5452098, 0.5474184, 0.5462912, 0.5482229, 
    0.5464844, 0.5494963, 0.5501525, 0.5497041, 0.5514268, 0.546388, 
    0.5483224, 0.5337988, 0.533884, 0.5342813, 0.5325354, 0.5324286, 
    0.5308291, 0.5322522, 0.5328584, 0.5343975, 0.5353082, 0.5361742, 
    0.5380787, 0.540207, 0.5431848, 0.5453253, 0.5467609, 0.5458805, 
    0.5466577, 0.5457889, 0.5453817, 0.5499067, 0.5473652, 0.5511789, 
    0.5509678, 0.5492416, 0.5509916, 0.5339439, 0.5334532, 0.5317501, 
    0.5330828, 0.5306549, 0.5320139, 0.5327955, 0.5358126, 0.5364755, 
    0.5370907, 0.5383056, 0.5398654, 0.5426033, 0.5449869, 0.547164, 
    0.5470045, 0.5470606, 0.5475472, 0.5463421, 0.5477451, 0.5479807, 
    0.5473649, 0.5509395, 0.5499179, 0.5509633, 0.5502981, 0.5336127, 
    0.5344384, 0.5339922, 0.5348313, 0.5342402, 0.5368697, 0.5376584, 
    0.5413507, 0.5398347, 0.5422475, 0.5400797, 0.5404638, 0.5423266, 
    0.5401968, 0.5448556, 0.5416968, 0.5475662, 0.5444099, 0.5477641, 
    0.5471546, 0.5481636, 0.5490676, 0.550205, 0.5523049, 0.5518185, 
    0.5535751, 0.5356696, 0.5367413, 0.5366468, 0.5377685, 0.5385983, 
    0.5403972, 0.5432844, 0.5421984, 0.5441922, 0.5445926, 0.5415636, 
    0.5434232, 0.5374586, 0.5384219, 0.5378482, 0.5357543, 0.5424489, 
    0.5390118, 0.5453607, 0.543497, 0.5489387, 0.5462317, 0.5515508, 
    0.5538274, 0.5559705, 0.5584776, 0.5373262, 0.5365978, 0.5379019, 
    0.5397071, 0.5413823, 0.5436107, 0.5438387, 0.5442564, 0.5453383, 
    0.5462483, 0.5443886, 0.5464764, 0.5386456, 0.5427473, 0.5363227, 
    0.5382564, 0.5396006, 0.5390107, 0.5420743, 0.5427967, 0.545734, 
    0.5442152, 0.5532655, 0.5492588, 0.560387, 0.5572739, 0.5363435, 
    0.5373236, 0.5407369, 0.5391124, 0.5437594, 0.5449042, 0.5458349, 
    0.5470252, 0.5471537, 0.5478591, 0.5467032, 0.5478134, 0.5436154, 
    0.5454908, 0.5403464, 0.541598, 0.5410221, 0.5403906, 0.5423399, 
    0.5444179, 0.5444621, 0.5451287, 0.5470083, 0.5437782, 0.5537835, 
    0.5476019, 0.5383927, 0.5402821, 0.5405517, 0.5398197, 0.5447894, 
    0.542988, 0.5478418, 0.5465294, 0.54868, 0.5476112, 0.547454, 0.5460817, 
    0.5452276, 0.5430706, 0.5413164, 0.5399258, 0.5402491, 0.5417768, 
    0.544545, 0.5471654, 0.5465913, 0.5485165, 0.5434223, 0.5455577, 
    0.5447323, 0.5468848, 0.5421696, 0.5461854, 0.5411439, 0.5415856, 
    0.5429522, 0.5457028, 0.5463112, 0.5469614, 0.5465601, 0.5446153, 
    0.5442966, 0.542919, 0.5425388, 0.5414894, 0.540621, 0.5414145, 
    0.5422481, 0.544616, 0.5467513, 0.5490805, 0.5496506, 0.5523751, 
    0.5501575, 0.553818, 0.5507063, 0.5560942, 0.5464178, 0.5506142, 
    0.5430143, 0.5438323, 0.5453125, 0.548709, 0.5468747, 0.5490199, 
    0.5442841, 0.5418296, 0.5411946, 0.5400104, 0.5412216, 0.5411231, 
    0.5422824, 0.5419098, 0.5446946, 0.5431985, 0.5474501, 0.5490029, 
    0.553391, 0.5560839, 0.5588266, 0.5600382, 0.560407, 0.5605612,
  0.5352148, 0.5380582, 0.5375048, 0.5398021, 0.5385271, 0.5400322, 
    0.5357906, 0.5381713, 0.5366509, 0.5354704, 0.5442732, 0.5399046, 
    0.5488271, 0.5460284, 0.5530713, 0.5483913, 0.5540172, 0.5529357, 
    0.5561931, 0.5552589, 0.5594364, 0.5566245, 0.5616076, 0.5587641, 
    0.5592086, 0.556532, 0.5407822, 0.5437285, 0.5406079, 0.5410275, 
    0.5408392, 0.5385535, 0.5374035, 0.5349976, 0.535434, 0.5372011, 
    0.5412163, 0.5398516, 0.5432934, 0.5432155, 0.5470589, 0.5453244, 
    0.5518032, 0.5499581, 0.5552979, 0.5539527, 0.5552347, 0.5548458, 
    0.5552398, 0.5532675, 0.5541121, 0.5523781, 0.5456492, 0.5476228, 
    0.5417464, 0.5382274, 0.535895, 0.5342428, 0.5344762, 0.5349215, 
    0.5372114, 0.5393682, 0.5410145, 0.542117, 0.5432043, 0.5465024, 
    0.5482512, 0.5521768, 0.5514671, 0.5526695, 0.5538189, 0.5557517, 
    0.5554333, 0.5562858, 0.5526375, 0.5550609, 0.5510631, 0.5521552, 
    0.5435011, 0.5402196, 0.5388284, 0.5376112, 0.5346558, 0.536696, 
    0.5358914, 0.5378063, 0.5390249, 0.538422, 0.5421472, 0.5406976, 
    0.5483549, 0.5450505, 0.5536848, 0.5516127, 0.554182, 0.5528702, 
    0.5551189, 0.5530949, 0.5566031, 0.5573686, 0.5568455, 0.558856, 
    0.5529828, 0.5552348, 0.5384052, 0.5385035, 0.5389615, 0.5369496, 
    0.5368266, 0.5349857, 0.5366235, 0.5373217, 0.5390955, 0.5401461, 
    0.5411456, 0.5433461, 0.5458087, 0.5492607, 0.551747, 0.5534166, 
    0.5523924, 0.5532966, 0.5522859, 0.5518125, 0.5570818, 0.5541201, 
    0.5585666, 0.5583201, 0.5563061, 0.5583479, 0.5385725, 0.5380069, 
    0.5360455, 0.5375802, 0.5347854, 0.5363491, 0.5372493, 0.5407281, 
    0.5414935, 0.5422041, 0.5436084, 0.5454132, 0.5485861, 0.5513536, 
    0.5538858, 0.5537, 0.5537654, 0.554332, 0.5529294, 0.5545623, 0.5548368, 
    0.5541196, 0.5582871, 0.5570949, 0.5583149, 0.5575384, 0.5381907, 
    0.5391427, 0.5386282, 0.5395958, 0.5389141, 0.5419488, 0.5428602, 
    0.5471337, 0.5453777, 0.5481734, 0.5456613, 0.5461061, 0.5482651, 
    0.5457968, 0.551201, 0.5475348, 0.554354, 0.5506832, 0.5545844, 
    0.5538749, 0.5550498, 0.5561033, 0.5574298, 0.5598819, 0.5593136, 
    0.5613672, 0.5405631, 0.5418006, 0.5416914, 0.5429875, 0.5439469, 
    0.546029, 0.5493764, 0.5481164, 0.5504304, 0.5508955, 0.5473804, 
    0.5495375, 0.5426292, 0.5437428, 0.5430796, 0.5406608, 0.5484069, 
    0.5444253, 0.5517881, 0.5496231, 0.555953, 0.5528008, 0.5590008, 
    0.5616624, 0.5641723, 0.5671139, 0.5424762, 0.5416348, 0.5431416, 
    0.5452299, 0.5471702, 0.5497551, 0.5500198, 0.5505049, 0.551762, 
    0.5528202, 0.5506585, 0.5530856, 0.5440016, 0.5487531, 0.541317, 
    0.5435515, 0.5451066, 0.544424, 0.5479724, 0.5488104, 0.5522221, 
    0.5504571, 0.5610051, 0.5563262, 0.5693584, 0.5657008, 0.541341, 
    0.5424732, 0.5464224, 0.5445417, 0.5499278, 0.5512575, 0.5523394, 
    0.5537242, 0.5538737, 0.5546951, 0.5533494, 0.5546418, 0.5497606, 
    0.5519393, 0.5459701, 0.5474203, 0.5467528, 0.5460213, 0.5482805, 
    0.5506925, 0.5507438, 0.5515184, 0.5537045, 0.5499496, 0.5616111, 
    0.5543956, 0.543709, 0.5458956, 0.5462079, 0.5453603, 0.5511241, 
    0.5490324, 0.554675, 0.5531472, 0.5556515, 0.5544064, 0.5542234, 
    0.5526264, 0.5516334, 0.5491282, 0.5470939, 0.5454831, 0.5458574, 
    0.5476276, 0.5508401, 0.5538874, 0.5532192, 0.555461, 0.5495364, 
    0.5520171, 0.5510578, 0.5535609, 0.5480831, 0.552747, 0.546894, 0.547406, 
    0.5489909, 0.5521858, 0.5528933, 0.5536499, 0.553183, 0.5509218, 
    0.5505516, 0.5489523, 0.5485112, 0.5472944, 0.5462882, 0.5472076, 
    0.548174, 0.5509226, 0.5534053, 0.5561183, 0.5567831, 0.5599639, 
    0.5573744, 0.5616514, 0.5580148, 0.5643173, 0.5530174, 0.5579073, 
    0.549063, 0.5500124, 0.5517321, 0.5556853, 0.5535491, 0.5560476, 
    0.550537, 0.5476888, 0.5469527, 0.545581, 0.546984, 0.5468699, 0.5482138, 
    0.5477818, 0.5510139, 0.5492766, 0.5542188, 0.5560278, 0.5611519, 
    0.5643051, 0.5675238, 0.5689481, 0.569382, 0.5695634,
  0.5840928, 0.5875039, 0.586839, 0.5896025, 0.5880677, 0.5898799, 0.5847825, 
    0.5876398, 0.585814, 0.5843988, 0.5950066, 0.5897262, 0.6005461, 
    0.5971375, 0.6057423, 0.6000144, 0.606905, 0.6055759, 0.6095858, 
    0.6084337, 0.6135982, 0.6101183, 0.6162958, 0.6127648, 0.6133156, 
    0.610004, 0.5907843, 0.5943465, 0.5905741, 0.5910804, 0.5908531, 
    0.5880995, 0.5867173, 0.5838327, 0.5843552, 0.5864743, 0.5913082, 
    0.5896623, 0.5938194, 0.5937251, 0.598391, 0.5962822, 0.6041864, 
    0.6019276, 0.6084818, 0.6068256, 0.6084039, 0.6079248, 0.6084102, 
    0.6059834, 0.6070218, 0.6048914, 0.5966766, 0.5990776, 0.5919484, 
    0.5877073, 0.5849076, 0.5829297, 0.5832089, 0.5837415, 0.5864867, 
    0.5890799, 0.5910646, 0.5923963, 0.5937116, 0.5977138, 0.5998436, 
    0.6046445, 0.6037745, 0.605249, 0.6066612, 0.6090413, 0.6086487, 
    0.6097001, 0.6052098, 0.6081898, 0.6032797, 0.6046181, 0.594071, 
    0.5901058, 0.5884302, 0.5869668, 0.5834236, 0.5858681, 0.5849032, 
    0.5872012, 0.5886666, 0.5879413, 0.5924327, 0.5906823, 0.59997, 
    0.5959496, 0.6064963, 0.6039529, 0.6071077, 0.6054955, 0.6082612, 
    0.6057714, 0.6100919, 0.6110377, 0.6103912, 0.6128787, 0.6056337, 
    0.608404, 0.5879211, 0.5880393, 0.5885903, 0.5861724, 0.5860248, 
    0.5838185, 0.5857811, 0.5866191, 0.5887516, 0.5900171, 0.5912228, 
    0.5938833, 0.5968704, 0.6010756, 0.6041175, 0.6061666, 0.6049091, 
    0.6060191, 0.6047784, 0.6041978, 0.6106831, 0.6070315, 0.6125202, 
    0.6122149, 0.6097252, 0.6122493, 0.5881223, 0.5874423, 0.585088, 
    0.5869296, 0.5835787, 0.585452, 0.5865321, 0.590719, 0.591643, 0.5925015, 
    0.5942009, 0.5963899, 0.600252, 0.6036355, 0.6067434, 0.606515, 
    0.6065954, 0.6072922, 0.6055681, 0.6075758, 0.6079137, 0.607031, 
    0.612174, 0.6106993, 0.6122084, 0.6112476, 0.5876632, 0.5888084, 
    0.5881893, 0.5893542, 0.5885333, 0.5921929, 0.593295, 0.598482, 
    0.5963468, 0.5997487, 0.5966913, 0.5972318, 0.5998605, 0.596856, 
    0.6034486, 0.5989705, 0.6073193, 0.6028146, 0.607603, 0.6067299, 
    0.6081761, 0.6094749, 0.6111133, 0.614151, 0.6134459, 0.6159966, 0.59052, 
    0.5920138, 0.5918819, 0.5934491, 0.5946111, 0.5971382, 0.6012169, 
    0.5996793, 0.6025052, 0.6030744, 0.5987824, 0.6014137, 0.5930157, 
    0.5943638, 0.5935606, 0.5906379, 0.6000335, 0.5951911, 0.6041679, 
    0.6015183, 0.6092895, 0.6054103, 0.6130582, 0.616364, 0.6194943, 
    0.6231793, 0.5928306, 0.5918136, 0.5936357, 0.5961673, 0.5985264, 
    0.6016796, 0.6020031, 0.6025964, 0.604136, 0.6054341, 0.6027843, 0.60576, 
    0.5946774, 0.6004558, 0.5914298, 0.5941321, 0.5960177, 0.5951895, 
    0.5995038, 0.6005259, 0.6047, 0.6025379, 0.6155463, 0.60975, 0.626003, 
    0.6214069, 0.5914588, 0.592827, 0.5976164, 0.5953322, 0.6018906, 
    0.6035177, 0.604844, 0.6065447, 0.6067286, 0.6077392, 0.6060841, 
    0.6076736, 0.6016863, 0.6043533, 0.5970665, 0.5988309, 0.5980184, 
    0.5971288, 0.5998793, 0.602826, 0.6028888, 0.6038374, 0.6065205, 
    0.6019173, 0.6163, 0.6073705, 0.5943229, 0.596976, 0.5973556, 0.5963256, 
    0.6033544, 0.6007968, 0.6077145, 0.6058357, 0.6089177, 0.6073838, 
    0.6071586, 0.6051962, 0.6039782, 0.6009138, 0.5984336, 0.5964748, 
    0.5969296, 0.5990835, 0.6030067, 0.6067454, 0.6059241, 0.6086828, 
    0.6014123, 0.6044487, 0.6032732, 0.6063439, 0.5996386, 0.6053442, 
    0.5981902, 0.5988135, 0.6007461, 0.6046556, 0.6055239, 0.6064534, 
    0.6058795, 0.6031066, 0.6026536, 0.6006989, 0.6001608, 0.5986777, 
    0.5974532, 0.598572, 0.5997495, 0.6031076, 0.6061528, 0.6094934, 
    0.6103141, 0.6142528, 0.6110448, 0.6163503, 0.6118369, 0.6196755, 
    0.6056762, 0.611704, 0.6008341, 0.6019941, 0.6040992, 0.6089593, 
    0.6063294, 0.6094062, 0.6026358, 0.5991581, 0.5982616, 0.5965938, 
    0.5982998, 0.5981608, 0.5997981, 0.5992714, 0.6032195, 0.601095, 
    0.6071531, 0.6093818, 0.6157289, 0.6196603, 0.6236942, 0.6254861, 
    0.6260327, 0.6262615,
  0.662225, 0.6677868, 0.6666974, 0.6712427, 0.6687127, 0.6717014, 0.6633441, 
    0.6680099, 0.665023, 0.6627212, 0.680266, 0.671447, 0.6897113, 0.683875, 
    0.6987641, 0.6887957, 0.7008164, 0.698471, 0.7055875, 0.7035305, 
    0.7128335, 0.706542, 0.7177785, 0.7113178, 0.712319, 0.7063369, 
    0.6732004, 0.6791539, 0.6728516, 0.6736922, 0.6733146, 0.6687649, 
    0.6664983, 0.6618037, 0.6626505, 0.6661009, 0.674071, 0.6713414, 
    0.6782679, 0.6781096, 0.6860121, 0.6824228, 0.6960331, 0.6920994, 
    0.703616, 0.700676, 0.7034774, 0.7026249, 0.7034885, 0.6991888, 
    0.7010232, 0.6972683, 0.6830918, 0.6871873, 0.6751373, 0.6681207, 
    0.6635474, 0.6603436, 0.6607946, 0.6616561, 0.6661212, 0.6703797, 
    0.673666, 0.6758847, 0.6780869, 0.6848563, 0.6885019, 0.6968353, 
    0.695313, 0.6978962, 0.7003852, 0.704614, 0.7039136, 0.7057922, 
    0.6978274, 0.7030962, 0.6944495, 0.6967888, 0.6786906, 0.6720753, 
    0.6693089, 0.6669066, 0.6611418, 0.6651112, 0.6635403, 0.6672907, 
    0.6696983, 0.668505, 0.6759456, 0.673031, 0.6887194, 0.6818594, 
    0.7000937, 0.6956248, 0.7011753, 0.6983294, 0.7032232, 0.6988151, 
    0.7064945, 0.7081947, 0.7070318, 0.7115247, 0.6985728, 0.7034776, 
    0.6684718, 0.6686661, 0.6695726, 0.6656078, 0.6653668, 0.6617806, 
    0.6649694, 0.6663377, 0.6698383, 0.6719286, 0.6739291, 0.6783752, 
    0.6834211, 0.6906249, 0.6959124, 0.6995118, 0.6972992, 0.6992517, 
    0.6970699, 0.696053, 0.7075566, 0.7010404, 0.7108741, 0.7103208, 
    0.7058372, 0.7103831, 0.6688025, 0.6676857, 0.6638407, 0.6668457, 
    0.6613926, 0.6644331, 0.6661955, 0.6730921, 0.6746283, 0.6760604, 
    0.6789089, 0.6826055, 0.6892046, 0.6950702, 0.7005305, 0.7001269, 
    0.700269, 0.7015022, 0.6984574, 0.7020051, 0.7026051, 0.7010394, 
    0.7102469, 0.7075857, 0.7103091, 0.7085731, 0.6680483, 0.6699319, 
    0.6689126, 0.6708323, 0.6694788, 0.6755452, 0.6773883, 0.6861677, 
    0.6825324, 0.6883389, 0.6831169, 0.6840355, 0.6885312, 0.6833965, 
    0.6947441, 0.6870037, 0.7015502, 0.6936396, 0.7020534, 0.7005067, 
    0.7030718, 0.7053891, 0.708331, 0.7138419, 0.7125561, 0.7172271, 
    0.6727619, 0.6752464, 0.6750264, 0.6776465, 0.6795993, 0.6838762, 
    0.690869, 0.6882196, 0.6931018, 0.694092, 0.6866816, 0.6912094, 
    0.6769204, 0.679183, 0.6778335, 0.6729574, 0.6888286, 0.6805772, 
    0.6960006, 0.6913904, 0.7050576, 0.6981798, 0.7118508, 0.7179043, 
    0.7237218, 0.7306814, 0.6766106, 0.6749126, 0.6779595, 0.6822281, 
    0.6862437, 0.6916696, 0.6922303, 0.6932602, 0.6959448, 0.6982216, 
    0.6935871, 0.6987951, 0.679711, 0.6895557, 0.6742734, 0.6787932, 
    0.6819746, 0.6805744, 0.6879182, 0.6896763, 0.6969326, 0.6931586, 
    0.7163985, 0.7058816, 0.7360994, 0.7273186, 0.6743217, 0.6766046, 
    0.6846904, 0.6808155, 0.6920352, 0.6948647, 0.697185, 0.7001794, 
    0.7005042, 0.7022953, 0.6993663, 0.7021788, 0.6916813, 0.6963251, 
    0.6837544, 0.6867647, 0.6853759, 0.6838603, 0.6885634, 0.6936595, 
    0.6937687, 0.6954227, 0.7001365, 0.6920815, 0.7177864, 0.701641, 
    0.6791142, 0.6836005, 0.6842462, 0.6824965, 0.6945798, 0.6901435, 
    0.7022514, 0.6989284, 0.7043933, 0.7016647, 0.7012655, 0.6978033, 
    0.6956689, 0.6903456, 0.6860849, 0.6827495, 0.6835217, 0.6871973, 
    0.693974, 0.700534, 0.6990843, 0.7039743, 0.6912071, 0.6964921, 
    0.6944382, 0.6998247, 0.6881497, 0.6980636, 0.6856692, 0.6867349, 
    0.6900561, 0.6968546, 0.6983795, 0.700018, 0.6990057, 0.694148, 
    0.6933596, 0.6899748, 0.6890475, 0.6865025, 0.6844124, 0.6863216, 
    0.6883402, 0.6941498, 0.6994875, 0.7054223, 0.7068934, 0.7140279, 
    0.7082076, 0.7178791, 0.709637, 0.7240613, 0.6986476, 0.7093968, 
    0.690208, 0.6922146, 0.6958805, 0.7044677, 0.6997991, 0.7052664, 
    0.6933287, 0.6873253, 0.6857911, 0.6829513, 0.6858563, 0.6856189, 
    0.6884237, 0.6875194, 0.6943446, 0.6906585, 0.7012556, 0.7052225, 
    0.7167342, 0.7240328, 0.7316638, 0.7351018, 0.7361567, 0.736599,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01157327, 0.01857286, 
    0.01857286, 0.01857286, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01857286, 0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01157327, 0.01157327, 0.01157327, 0.01952015, 0.01952015, 
    0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01952015, 0.01857286, 
    0.01952015, 0.01952015, 0.01857286, 0.01952015, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01157327, 0.01157327, 
    0.01952015, 0.01952015, 0.01857286, 0.01952015, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01157327, 0.01857286, 0.01952015, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01157327, 0.01857286, 0.01157327, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01157327, 0.01157327, 0.01157327, 
    0.01157327, 0.01157327 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.422945e-11, 3.437952e-11, 3.435026e-11, 3.447139e-11, 3.440414e-11, 
    3.448341e-11, 3.425968e-11, 3.438524e-11, 3.430502e-11, 3.424264e-11, 
    3.47064e-11, 3.447651e-11, 3.494549e-11, 3.479857e-11, 3.516766e-11, 
    3.492253e-11, 3.521709e-11, 3.516048e-11, 3.533072e-11, 3.528187e-11, 
    3.549976e-11, 3.535315e-11, 3.561276e-11, 3.546467e-11, 3.548779e-11, 
    3.534813e-11, 3.4523e-11, 3.467803e-11, 3.451375e-11, 3.453585e-11, 
    3.452589e-11, 3.440538e-11, 3.434469e-11, 3.421765e-11, 3.424065e-11, 
    3.433393e-11, 3.454553e-11, 3.447359e-11, 3.465475e-11, 3.465066e-11, 
    3.485253e-11, 3.476146e-11, 3.510118e-11, 3.50045e-11, 3.528387e-11, 
    3.521351e-11, 3.528049e-11, 3.526012e-11, 3.528065e-11, 3.517756e-11, 
    3.522165e-11, 3.513096e-11, 3.477894e-11, 3.488251e-11, 3.457363e-11, 
    3.438814e-11, 3.426503e-11, 3.417778e-11, 3.419003e-11, 3.421356e-11, 
    3.43344e-11, 3.444809e-11, 3.453482e-11, 3.45928e-11, 3.464997e-11, 
    3.482328e-11, 3.491502e-11, 3.512065e-11, 3.508349e-11, 3.514635e-11, 
    3.520647e-11, 3.530742e-11, 3.529077e-11, 3.533523e-11, 3.51445e-11, 
    3.527121e-11, 3.506202e-11, 3.51192e-11, 3.46659e-11, 3.449314e-11, 
    3.441979e-11, 3.435556e-11, 3.419949e-11, 3.430723e-11, 3.42647e-11, 
    3.436572e-11, 3.442996e-11, 3.439812e-11, 3.459435e-11, 3.451797e-11, 
    3.49204e-11, 3.474693e-11, 3.51995e-11, 3.509103e-11, 3.52254e-11, 
    3.51568e-11, 3.527428e-11, 3.516848e-11, 3.535173e-11, 3.539168e-11, 
    3.53643e-11, 3.546918e-11, 3.516239e-11, 3.528013e-11, 3.439744e-11, 
    3.440263e-11, 3.442673e-11, 3.432055e-11, 3.431404e-11, 3.42168e-11, 
    3.430323e-11, 3.434008e-11, 3.443358e-11, 3.448889e-11, 3.454149e-11, 
    3.465731e-11, 3.478669e-11, 3.496779e-11, 3.509801e-11, 3.518532e-11, 
    3.513173e-11, 3.517898e-11, 3.512608e-11, 3.510125e-11, 3.53766e-11, 
    3.522192e-11, 3.545399e-11, 3.544114e-11, 3.5336e-11, 3.544249e-11, 
    3.44062e-11, 3.437631e-11, 3.42728e-11, 3.435374e-11, 3.420614e-11, 
    3.428873e-11, 3.433618e-11, 3.451952e-11, 3.455979e-11, 3.45972e-11, 
    3.467103e-11, 3.476584e-11, 3.493237e-11, 3.507733e-11, 3.520982e-11, 
    3.520005e-11, 3.520345e-11, 3.523301e-11, 3.515965e-11, 3.524498e-11, 
    3.525927e-11, 3.52218e-11, 3.543931e-11, 3.537713e-11, 3.544072e-11, 
    3.540017e-11, 3.438597e-11, 3.44361e-11, 3.440893e-11, 3.445995e-11, 
    3.442393e-11, 3.45838e-11, 3.463171e-11, 3.485623e-11, 3.476397e-11, 
    3.491075e-11, 3.47788e-11, 3.480217e-11, 3.491542e-11, 3.478583e-11, 
    3.506923e-11, 3.487698e-11, 3.523412e-11, 3.504198e-11, 3.524609e-11, 
    3.520895e-11, 3.527031e-11, 3.532534e-11, 3.53945e-11, 3.552234e-11, 
    3.549265e-11, 3.55996e-11, 3.451091e-11, 3.457601e-11, 3.457026e-11, 
    3.463841e-11, 3.468882e-11, 3.479825e-11, 3.497384e-11, 3.490771e-11, 
    3.502897e-11, 3.505333e-11, 3.486898e-11, 3.498211e-11, 3.461926e-11, 
    3.467777e-11, 3.464288e-11, 3.45155e-11, 3.492263e-11, 3.471351e-11, 
    3.509973e-11, 3.498629e-11, 3.531739e-11, 3.515263e-11, 3.547632e-11, 
    3.561492e-11, 3.574538e-11, 3.589796e-11, 3.461154e-11, 3.45672e-11, 
    3.464645e-11, 3.475623e-11, 3.485805e-11, 3.499364e-11, 3.500747e-11, 
    3.503283e-11, 3.50986e-11, 3.515399e-11, 3.504078e-11, 3.516777e-11, 
    3.469132e-11, 3.494079e-11, 3.454999e-11, 3.466757e-11, 3.474925e-11, 
    3.471338e-11, 3.489969e-11, 3.494359e-11, 3.512224e-11, 3.502985e-11, 
    3.55806e-11, 3.53367e-11, 3.601418e-11, 3.582461e-11, 3.455169e-11, 
    3.461123e-11, 3.481877e-11, 3.471998e-11, 3.500259e-11, 3.507223e-11, 
    3.51288e-11, 3.520124e-11, 3.520898e-11, 3.525192e-11, 3.518149e-11, 
    3.524907e-11, 3.499354e-11, 3.510765e-11, 3.479463e-11, 3.48707e-11, 
    3.483566e-11, 3.479719e-11, 3.491572e-11, 3.504213e-11, 3.504478e-11, 
    3.508529e-11, 3.519961e-11, 3.500306e-11, 3.561197e-11, 3.523561e-11, 
    3.46762e-11, 3.479105e-11, 3.480741e-11, 3.47629e-11, 3.506515e-11, 
    3.495556e-11, 3.525088e-11, 3.517094e-11, 3.530179e-11, 3.523674e-11, 
    3.522709e-11, 3.514358e-11, 3.509152e-11, 3.49603e-11, 3.48535e-11, 
    3.476893e-11, 3.478851e-11, 3.488144e-11, 3.504976e-11, 3.520924e-11, 
    3.517425e-11, 3.529138e-11, 3.498133e-11, 3.511125e-11, 3.506094e-11, 
    3.519195e-11, 3.490581e-11, 3.515011e-11, 3.484338e-11, 3.487019e-11, 
    3.495328e-11, 3.512063e-11, 3.515759e-11, 3.519716e-11, 3.517266e-11, 
    3.505431e-11, 3.503489e-11, 3.495102e-11, 3.492784e-11, 3.486401e-11, 
    3.481111e-11, 3.485938e-11, 3.491001e-11, 3.505407e-11, 3.518396e-11, 
    3.532568e-11, 3.536037e-11, 3.552613e-11, 3.539112e-11, 3.561388e-11, 
    3.542442e-11, 3.575242e-11, 3.516416e-11, 3.541959e-11, 3.495707e-11, 
    3.500678e-11, 3.50968e-11, 3.530346e-11, 3.519178e-11, 3.532235e-11, 
    3.503411e-11, 3.488471e-11, 3.484604e-11, 3.477402e-11, 3.484761e-11, 
    3.484163e-11, 3.491211e-11, 3.488939e-11, 3.505875e-11, 3.496774e-11, 
    3.522636e-11, 3.532088e-11, 3.558797e-11, 3.575186e-11, 3.591887e-11, 
    3.59926e-11, 3.601505e-11, 3.602439e-11,
  1.908592e-11, 1.923004e-11, 1.920199e-11, 1.931847e-11, 1.925383e-11, 
    1.933014e-11, 1.911511e-11, 1.923577e-11, 1.915871e-11, 1.909888e-11, 
    1.954523e-11, 1.932367e-11, 1.977636e-11, 1.963434e-11, 1.999181e-11, 
    1.975424e-11, 2.003984e-11, 1.998495e-11, 2.015033e-11, 2.01029e-11, 
    2.031496e-11, 2.017224e-11, 2.042521e-11, 2.028085e-11, 2.030341e-11, 
    2.016754e-11, 1.936819e-11, 1.951759e-11, 1.935935e-11, 1.938062e-11, 
    1.937108e-11, 1.925516e-11, 1.919684e-11, 1.907492e-11, 1.909704e-11, 
    1.918659e-11, 1.939019e-11, 1.932099e-11, 1.949558e-11, 1.949163e-11, 
    1.968664e-11, 1.959863e-11, 1.992745e-11, 1.98338e-11, 2.010488e-11, 
    2.003658e-11, 2.010167e-11, 2.008193e-11, 2.010193e-11, 2.000179e-11, 
    2.004467e-11, 1.995664e-11, 1.96151e-11, 1.971525e-11, 1.941709e-11, 
    1.92386e-11, 1.912039e-11, 1.903668e-11, 1.90485e-11, 1.907106e-11, 
    1.918712e-11, 1.929648e-11, 1.937997e-11, 1.94359e-11, 1.949106e-11, 
    1.965836e-11, 1.974713e-11, 1.994641e-11, 1.99104e-11, 1.997142e-11, 
    2.002979e-11, 2.012792e-11, 2.011176e-11, 2.015503e-11, 1.996981e-11, 
    2.009284e-11, 1.988989e-11, 1.994533e-11, 1.950605e-11, 1.933965e-11, 
    1.926907e-11, 1.920738e-11, 1.90576e-11, 1.916099e-11, 1.912021e-11, 
    1.921729e-11, 1.927907e-11, 1.924851e-11, 1.943743e-11, 1.93639e-11, 
    1.97524e-11, 1.958471e-11, 2.002298e-11, 1.991779e-11, 2.004823e-11, 
    1.998163e-11, 2.009578e-11, 1.999303e-11, 2.017115e-11, 2.021e-11, 
    2.018345e-11, 2.028553e-11, 1.998734e-11, 2.010167e-11, 1.924765e-11, 
    1.925263e-11, 1.927586e-11, 1.917384e-11, 1.916761e-11, 1.907432e-11, 
    1.915732e-11, 1.919271e-11, 1.928265e-11, 1.933593e-11, 1.938662e-11, 
    1.949825e-11, 1.962319e-11, 1.979839e-11, 1.99246e-11, 2.000937e-11, 
    1.995737e-11, 2.000328e-11, 1.995197e-11, 1.992793e-11, 2.019544e-11, 
    2.004507e-11, 2.027084e-11, 2.025832e-11, 2.015606e-11, 2.025973e-11, 
    1.925613e-11, 1.922746e-11, 1.912803e-11, 1.920582e-11, 1.906417e-11, 
    1.914341e-11, 1.918903e-11, 1.936543e-11, 1.940427e-11, 1.944031e-11, 
    1.951156e-11, 1.960313e-11, 1.976414e-11, 1.990463e-11, 2.003319e-11, 
    2.002376e-11, 2.002708e-11, 2.005584e-11, 1.998463e-11, 2.006753e-11, 
    2.008146e-11, 2.004506e-11, 2.025665e-11, 2.019612e-11, 2.025806e-11, 
    2.021864e-11, 1.923678e-11, 1.928504e-11, 1.925896e-11, 1.930802e-11, 
    1.927345e-11, 1.942734e-11, 1.947357e-11, 1.969042e-11, 1.960132e-11, 
    1.974319e-11, 1.961572e-11, 1.963828e-11, 1.974782e-11, 1.96226e-11, 
    1.989687e-11, 1.971077e-11, 2.005695e-11, 1.987057e-11, 2.006866e-11, 
    2.003263e-11, 2.009229e-11, 2.014577e-11, 2.021312e-11, 2.03376e-11, 
    2.030875e-11, 2.041302e-11, 1.935708e-11, 1.941983e-11, 1.941431e-11, 
    1.948005e-11, 1.952873e-11, 1.963438e-11, 1.980427e-11, 1.974032e-11, 
    1.985777e-11, 1.988138e-11, 1.970296e-11, 1.981244e-11, 1.946187e-11, 
    1.951836e-11, 1.948472e-11, 1.936202e-11, 1.975504e-11, 1.955298e-11, 
    1.992669e-11, 1.981679e-11, 2.013814e-11, 1.997809e-11, 2.029288e-11, 
    2.042797e-11, 2.055542e-11, 2.070469e-11, 1.945412e-11, 1.941144e-11, 
    1.948788e-11, 1.959381e-11, 1.969229e-11, 1.982349e-11, 1.983693e-11, 
    1.986155e-11, 1.992537e-11, 1.997909e-11, 1.986934e-11, 1.999257e-11, 
    1.953146e-11, 1.977262e-11, 1.939531e-11, 1.950865e-11, 1.958756e-11, 
    1.955293e-11, 1.973302e-11, 1.977555e-11, 1.994871e-11, 1.985913e-11, 
    2.03946e-11, 2.015706e-11, 2.081861e-11, 2.063298e-11, 1.939653e-11, 
    1.945397e-11, 1.965433e-11, 1.955891e-11, 1.983226e-11, 1.989975e-11, 
    1.995468e-11, 2.002498e-11, 2.003257e-11, 2.007427e-11, 2.000596e-11, 
    2.007157e-11, 1.982377e-11, 1.993437e-11, 1.96314e-11, 1.970498e-11, 
    1.967112e-11, 1.963399e-11, 1.974865e-11, 1.987106e-11, 1.987368e-11, 
    1.991299e-11, 2.002391e-11, 1.983337e-11, 2.042532e-11, 2.0059e-11, 
    1.951667e-11, 1.962759e-11, 1.964346e-11, 1.960045e-11, 1.989298e-11, 
    1.978681e-11, 2.007326e-11, 1.999569e-11, 2.012284e-11, 2.005962e-11, 
    2.005032e-11, 1.996925e-11, 1.991883e-11, 1.979167e-11, 1.968842e-11, 
    1.960668e-11, 1.962568e-11, 1.97155e-11, 1.987855e-11, 2.003326e-11, 
    1.999933e-11, 2.011316e-11, 1.981239e-11, 1.993831e-11, 1.98896e-11, 
    2.001669e-11, 1.973862e-11, 1.997531e-11, 1.967828e-11, 1.970426e-11, 
    1.97847e-11, 1.994686e-11, 1.99828e-11, 2.00212e-11, 1.999751e-11, 
    1.98827e-11, 1.986392e-11, 1.978274e-11, 1.976035e-11, 1.969861e-11, 
    1.964754e-11, 1.969419e-11, 1.974323e-11, 1.988275e-11, 2.000879e-11, 
    2.014653e-11, 2.018029e-11, 2.034173e-11, 2.021027e-11, 2.042737e-11, 
    2.024273e-11, 2.056272e-11, 1.998906e-11, 2.023732e-11, 1.978837e-11, 
    1.983656e-11, 1.992383e-11, 2.012452e-11, 2.001609e-11, 2.014293e-11, 
    1.986319e-11, 1.97186e-11, 1.968126e-11, 1.961165e-11, 1.968285e-11, 
    1.967706e-11, 1.974527e-11, 1.972334e-11, 1.988739e-11, 1.979921e-11, 
    2.005009e-11, 2.014192e-11, 2.040208e-11, 2.056214e-11, 2.072553e-11, 
    2.07978e-11, 2.081982e-11, 2.082902e-11,
  1.784495e-11, 1.800267e-11, 1.797196e-11, 1.809951e-11, 1.802871e-11, 
    1.811229e-11, 1.787688e-11, 1.800894e-11, 1.792459e-11, 1.785913e-11, 
    1.834811e-11, 1.810521e-11, 1.860187e-11, 1.84459e-11, 1.883876e-11, 
    1.857756e-11, 1.889161e-11, 1.883121e-11, 1.901327e-11, 1.896104e-11, 
    1.919468e-11, 1.903739e-11, 1.931627e-11, 1.915707e-11, 1.918194e-11, 
    1.903221e-11, 1.815398e-11, 1.831779e-11, 1.81443e-11, 1.816761e-11, 
    1.815715e-11, 1.803017e-11, 1.796632e-11, 1.783292e-11, 1.785711e-11, 
    1.79551e-11, 1.81781e-11, 1.810228e-11, 1.829364e-11, 1.828931e-11, 
    1.850332e-11, 1.84067e-11, 1.876797e-11, 1.866499e-11, 1.896321e-11, 
    1.888803e-11, 1.895968e-11, 1.893794e-11, 1.895996e-11, 1.884974e-11, 
    1.889693e-11, 1.880007e-11, 1.842478e-11, 1.853474e-11, 1.820758e-11, 
    1.801204e-11, 1.788266e-11, 1.779109e-11, 1.780403e-11, 1.782869e-11, 
    1.795568e-11, 1.807542e-11, 1.81669e-11, 1.82282e-11, 1.828869e-11, 
    1.847227e-11, 1.856976e-11, 1.878882e-11, 1.874921e-11, 1.881633e-11, 
    1.888056e-11, 1.898858e-11, 1.897078e-11, 1.901844e-11, 1.881456e-11, 
    1.894996e-11, 1.872666e-11, 1.878762e-11, 1.830513e-11, 1.812272e-11, 
    1.804541e-11, 1.797786e-11, 1.781397e-11, 1.792708e-11, 1.788246e-11, 
    1.798871e-11, 1.805635e-11, 1.802288e-11, 1.822988e-11, 1.814928e-11, 
    1.857555e-11, 1.839143e-11, 1.887306e-11, 1.875734e-11, 1.890084e-11, 
    1.882756e-11, 1.89532e-11, 1.884011e-11, 1.903619e-11, 1.9079e-11, 
    1.904974e-11, 1.916223e-11, 1.883385e-11, 1.895968e-11, 1.802195e-11, 
    1.80274e-11, 1.805284e-11, 1.794115e-11, 1.793433e-11, 1.783226e-11, 
    1.792307e-11, 1.79618e-11, 1.806028e-11, 1.811864e-11, 1.817418e-11, 
    1.829657e-11, 1.843365e-11, 1.862607e-11, 1.876483e-11, 1.885808e-11, 
    1.880088e-11, 1.885138e-11, 1.879493e-11, 1.87685e-11, 1.906295e-11, 
    1.889737e-11, 1.914604e-11, 1.913224e-11, 1.901957e-11, 1.91338e-11, 
    1.803123e-11, 1.799984e-11, 1.789101e-11, 1.797616e-11, 1.782116e-11, 
    1.790785e-11, 1.795777e-11, 1.815097e-11, 1.819353e-11, 1.823303e-11, 
    1.831117e-11, 1.841164e-11, 1.858845e-11, 1.874286e-11, 1.88843e-11, 
    1.887392e-11, 1.887757e-11, 1.890922e-11, 1.883086e-11, 1.89221e-11, 
    1.893743e-11, 1.889736e-11, 1.913039e-11, 1.90637e-11, 1.913195e-11, 
    1.908851e-11, 1.801004e-11, 1.80629e-11, 1.803433e-11, 1.808806e-11, 
    1.80502e-11, 1.821882e-11, 1.826951e-11, 1.850747e-11, 1.840966e-11, 
    1.856543e-11, 1.842546e-11, 1.845023e-11, 1.857052e-11, 1.843301e-11, 
    1.873433e-11, 1.852982e-11, 1.891045e-11, 1.870541e-11, 1.892333e-11, 
    1.888368e-11, 1.894935e-11, 1.900824e-11, 1.908243e-11, 1.921964e-11, 
    1.918783e-11, 1.930282e-11, 1.814181e-11, 1.821059e-11, 1.820453e-11, 
    1.827662e-11, 1.833e-11, 1.844594e-11, 1.863253e-11, 1.856227e-11, 
    1.869135e-11, 1.87173e-11, 1.852125e-11, 1.864152e-11, 1.825668e-11, 
    1.831863e-11, 1.828174e-11, 1.814723e-11, 1.857845e-11, 1.835661e-11, 
    1.876712e-11, 1.86463e-11, 1.899983e-11, 1.882366e-11, 1.917033e-11, 
    1.931932e-11, 1.945999e-11, 1.96249e-11, 1.824817e-11, 1.820139e-11, 
    1.82852e-11, 1.840141e-11, 1.850952e-11, 1.865366e-11, 1.866844e-11, 
    1.86955e-11, 1.876568e-11, 1.882477e-11, 1.870406e-11, 1.883959e-11, 
    1.8333e-11, 1.859776e-11, 1.818371e-11, 1.830797e-11, 1.839455e-11, 
    1.835656e-11, 1.855425e-11, 1.860098e-11, 1.879135e-11, 1.869284e-11, 
    1.92825e-11, 1.902068e-11, 1.975085e-11, 1.954566e-11, 1.818505e-11, 
    1.824801e-11, 1.846785e-11, 1.836311e-11, 1.86633e-11, 1.87375e-11, 
    1.879792e-11, 1.887526e-11, 1.888362e-11, 1.892951e-11, 1.885433e-11, 
    1.892654e-11, 1.865397e-11, 1.877557e-11, 1.844267e-11, 1.852346e-11, 
    1.848628e-11, 1.844552e-11, 1.857143e-11, 1.870595e-11, 1.870883e-11, 
    1.875206e-11, 1.887408e-11, 1.866452e-11, 1.931639e-11, 1.89127e-11, 
    1.831677e-11, 1.843849e-11, 1.845591e-11, 1.84087e-11, 1.873006e-11, 
    1.861335e-11, 1.892839e-11, 1.884303e-11, 1.898298e-11, 1.891338e-11, 
    1.890315e-11, 1.881394e-11, 1.875849e-11, 1.861869e-11, 1.850527e-11, 
    1.841554e-11, 1.843639e-11, 1.853501e-11, 1.87142e-11, 1.888437e-11, 
    1.884704e-11, 1.897233e-11, 1.864147e-11, 1.87799e-11, 1.872635e-11, 
    1.886613e-11, 1.856041e-11, 1.88206e-11, 1.849414e-11, 1.852267e-11, 
    1.861103e-11, 1.878931e-11, 1.882885e-11, 1.88711e-11, 1.884503e-11, 
    1.871875e-11, 1.86981e-11, 1.860889e-11, 1.858428e-11, 1.851646e-11, 
    1.846038e-11, 1.851161e-11, 1.856548e-11, 1.871881e-11, 1.885744e-11, 
    1.900907e-11, 1.904626e-11, 1.92242e-11, 1.907929e-11, 1.931865e-11, 
    1.911506e-11, 1.946805e-11, 1.883574e-11, 1.91091e-11, 1.861506e-11, 
    1.866803e-11, 1.876398e-11, 1.898484e-11, 1.886548e-11, 1.900511e-11, 
    1.86973e-11, 1.853842e-11, 1.849741e-11, 1.842099e-11, 1.849916e-11, 
    1.849279e-11, 1.856771e-11, 1.854362e-11, 1.872391e-11, 1.862698e-11, 
    1.890289e-11, 1.9004e-11, 1.929075e-11, 1.946741e-11, 1.964793e-11, 
    1.972783e-11, 1.975218e-11, 1.976236e-11,
  1.830173e-11, 1.84754e-11, 1.844157e-11, 1.85821e-11, 1.850408e-11, 
    1.859619e-11, 1.833688e-11, 1.848231e-11, 1.83894e-11, 1.831733e-11, 
    1.885627e-11, 1.858838e-11, 1.913647e-11, 1.89642e-11, 1.939838e-11, 
    1.910962e-11, 1.945685e-11, 1.939001e-11, 1.95915e-11, 1.953368e-11, 
    1.979248e-11, 1.961822e-11, 1.992727e-11, 1.975079e-11, 1.977835e-11, 
    1.961248e-11, 1.864214e-11, 1.882282e-11, 1.863146e-11, 1.865717e-11, 
    1.864563e-11, 1.850569e-11, 1.843537e-11, 1.828849e-11, 1.831511e-11, 
    1.842301e-11, 1.866873e-11, 1.858515e-11, 1.879615e-11, 1.879137e-11, 
    1.90276e-11, 1.892092e-11, 1.932007e-11, 1.920621e-11, 1.953609e-11, 
    1.945288e-11, 1.953218e-11, 1.950811e-11, 1.953249e-11, 1.941052e-11, 
    1.946273e-11, 1.935557e-11, 1.894087e-11, 1.906231e-11, 1.870124e-11, 
    1.848573e-11, 1.834324e-11, 1.824245e-11, 1.825669e-11, 1.828383e-11, 
    1.842364e-11, 1.855555e-11, 1.865638e-11, 1.872397e-11, 1.879069e-11, 
    1.899333e-11, 1.910099e-11, 1.934313e-11, 1.929932e-11, 1.937356e-11, 
    1.944461e-11, 1.956417e-11, 1.954447e-11, 1.959723e-11, 1.93716e-11, 
    1.952142e-11, 1.927439e-11, 1.93418e-11, 1.880885e-11, 1.860768e-11, 
    1.852249e-11, 1.844807e-11, 1.826763e-11, 1.839215e-11, 1.834302e-11, 
    1.846001e-11, 1.853454e-11, 1.849766e-11, 1.872582e-11, 1.863696e-11, 
    1.910738e-11, 1.890407e-11, 1.943631e-11, 1.930831e-11, 1.946705e-11, 
    1.938597e-11, 1.9525e-11, 1.939985e-11, 1.961688e-11, 1.96643e-11, 
    1.963189e-11, 1.975651e-11, 1.939293e-11, 1.953218e-11, 1.849663e-11, 
    1.850264e-11, 1.853066e-11, 1.840764e-11, 1.840013e-11, 1.828776e-11, 
    1.838773e-11, 1.843038e-11, 1.853886e-11, 1.860318e-11, 1.866441e-11, 
    1.879939e-11, 1.895068e-11, 1.916321e-11, 1.931659e-11, 1.941974e-11, 
    1.935646e-11, 1.941232e-11, 1.934988e-11, 1.932065e-11, 1.964653e-11, 
    1.946322e-11, 1.973856e-11, 1.972328e-11, 1.959849e-11, 1.9725e-11, 
    1.850686e-11, 1.847228e-11, 1.835243e-11, 1.844619e-11, 1.827554e-11, 
    1.837097e-11, 1.842595e-11, 1.863882e-11, 1.868574e-11, 1.872931e-11, 
    1.881549e-11, 1.892637e-11, 1.912163e-11, 1.929231e-11, 1.944874e-11, 
    1.943726e-11, 1.94413e-11, 1.947633e-11, 1.938963e-11, 1.949058e-11, 
    1.950755e-11, 1.94632e-11, 1.972123e-11, 1.964735e-11, 1.972295e-11, 
    1.967483e-11, 1.848352e-11, 1.854175e-11, 1.851027e-11, 1.856948e-11, 
    1.852776e-11, 1.871364e-11, 1.876954e-11, 1.903219e-11, 1.892419e-11, 
    1.909621e-11, 1.894162e-11, 1.896897e-11, 1.910184e-11, 1.894996e-11, 
    1.928288e-11, 1.905687e-11, 1.947769e-11, 1.925091e-11, 1.949194e-11, 
    1.944807e-11, 1.952074e-11, 1.958593e-11, 1.96681e-11, 1.982014e-11, 
    1.978488e-11, 1.991235e-11, 1.862872e-11, 1.870456e-11, 1.869787e-11, 
    1.877737e-11, 1.883627e-11, 1.896424e-11, 1.917034e-11, 1.909271e-11, 
    1.923534e-11, 1.926404e-11, 1.904739e-11, 1.918027e-11, 1.875539e-11, 
    1.882373e-11, 1.878302e-11, 1.86347e-11, 1.911059e-11, 1.886565e-11, 
    1.931913e-11, 1.918556e-11, 1.957663e-11, 1.938167e-11, 1.976548e-11, 
    1.993066e-11, 2.008671e-11, 2.026981e-11, 1.8746e-11, 1.869441e-11, 
    1.878684e-11, 1.891509e-11, 1.903445e-11, 1.919369e-11, 1.921002e-11, 
    1.923994e-11, 1.931753e-11, 1.938289e-11, 1.92494e-11, 1.939928e-11, 
    1.88396e-11, 1.913192e-11, 1.867492e-11, 1.881198e-11, 1.890751e-11, 
    1.886558e-11, 1.908385e-11, 1.913547e-11, 1.934592e-11, 1.923699e-11, 
    1.988984e-11, 1.959972e-11, 2.040975e-11, 2.018181e-11, 1.867639e-11, 
    1.874582e-11, 1.898843e-11, 1.887281e-11, 1.920435e-11, 1.928638e-11, 
    1.935318e-11, 1.943875e-11, 1.944799e-11, 1.949879e-11, 1.941559e-11, 
    1.94955e-11, 1.919403e-11, 1.932847e-11, 1.896062e-11, 1.904984e-11, 
    1.900877e-11, 1.896377e-11, 1.910282e-11, 1.92515e-11, 1.925468e-11, 
    1.930248e-11, 1.943747e-11, 1.920569e-11, 1.992743e-11, 1.948021e-11, 
    1.882167e-11, 1.895602e-11, 1.897524e-11, 1.892312e-11, 1.927815e-11, 
    1.914914e-11, 1.949755e-11, 1.940309e-11, 1.955797e-11, 1.948093e-11, 
    1.946961e-11, 1.937091e-11, 1.930958e-11, 1.915505e-11, 1.902975e-11, 
    1.893067e-11, 1.895369e-11, 1.90626e-11, 1.926061e-11, 1.944883e-11, 
    1.940753e-11, 1.954618e-11, 1.918021e-11, 1.933327e-11, 1.927405e-11, 
    1.942865e-11, 1.909065e-11, 1.937831e-11, 1.901746e-11, 1.904897e-11, 
    1.914659e-11, 1.934367e-11, 1.93874e-11, 1.943415e-11, 1.94053e-11, 
    1.926565e-11, 1.924282e-11, 1.914421e-11, 1.911703e-11, 1.90421e-11, 
    1.898018e-11, 1.903675e-11, 1.909625e-11, 1.926571e-11, 1.941904e-11, 
    1.958686e-11, 1.962804e-11, 1.98252e-11, 1.966463e-11, 1.992994e-11, 
    1.970428e-11, 2.009568e-11, 1.939504e-11, 1.969765e-11, 1.915103e-11, 
    1.920957e-11, 1.931566e-11, 1.956004e-11, 1.942792e-11, 1.958247e-11, 
    1.924192e-11, 1.906637e-11, 1.902107e-11, 1.893669e-11, 1.9023e-11, 
    1.901597e-11, 1.909872e-11, 1.907211e-11, 1.927135e-11, 1.91642e-11, 
    1.946933e-11, 1.958125e-11, 1.989897e-11, 2.009495e-11, 2.029538e-11, 
    2.038417e-11, 2.041123e-11, 2.042255e-11,
  1.973896e-11, 1.992292e-11, 1.988708e-11, 2.003602e-11, 1.995332e-11, 
    2.005096e-11, 1.977617e-11, 1.993025e-11, 1.983181e-11, 1.975547e-11, 
    2.032691e-11, 2.004268e-11, 2.062452e-11, 2.044147e-11, 2.090306e-11, 
    2.059598e-11, 2.096529e-11, 2.089415e-11, 2.110866e-11, 2.104708e-11, 
    2.132287e-11, 2.113712e-11, 2.146663e-11, 2.127841e-11, 2.13078e-11, 
    2.113101e-11, 2.009968e-11, 2.02914e-11, 2.008836e-11, 2.011563e-11, 
    2.010339e-11, 1.995503e-11, 1.988051e-11, 1.972493e-11, 1.975312e-11, 
    1.986741e-11, 2.012789e-11, 2.003924e-11, 2.026306e-11, 2.025799e-11, 
    2.050881e-11, 2.03955e-11, 2.081973e-11, 2.069864e-11, 2.104964e-11, 
    2.096105e-11, 2.104548e-11, 2.101986e-11, 2.104581e-11, 2.091597e-11, 
    2.097155e-11, 2.08575e-11, 2.04167e-11, 2.054569e-11, 2.016237e-11, 
    1.993389e-11, 1.978291e-11, 1.967619e-11, 1.969126e-11, 1.972001e-11, 
    1.986808e-11, 2.000787e-11, 2.011478e-11, 2.018648e-11, 2.025726e-11, 
    2.047243e-11, 2.058681e-11, 2.084427e-11, 2.079766e-11, 2.087665e-11, 
    2.095225e-11, 2.107956e-11, 2.105857e-11, 2.111477e-11, 2.087455e-11, 
    2.103403e-11, 2.077113e-11, 2.084285e-11, 2.027658e-11, 2.006314e-11, 
    1.997285e-11, 1.989397e-11, 1.970285e-11, 1.983472e-11, 1.978268e-11, 
    1.990661e-11, 1.99856e-11, 1.994651e-11, 2.018844e-11, 2.009419e-11, 
    2.05936e-11, 2.037762e-11, 2.094342e-11, 2.080722e-11, 2.097615e-11, 
    2.088984e-11, 2.103785e-11, 2.090462e-11, 2.11357e-11, 2.118622e-11, 
    2.115169e-11, 2.12845e-11, 2.089725e-11, 2.104548e-11, 1.994542e-11, 
    1.995179e-11, 1.998149e-11, 1.985113e-11, 1.984317e-11, 1.972416e-11, 
    1.983003e-11, 1.987522e-11, 1.999018e-11, 2.005836e-11, 2.01233e-11, 
    2.02665e-11, 2.042712e-11, 2.065293e-11, 2.081603e-11, 2.092578e-11, 
    2.085844e-11, 2.091788e-11, 2.085144e-11, 2.082034e-11, 2.116729e-11, 
    2.097207e-11, 2.126537e-11, 2.124907e-11, 2.111611e-11, 2.125091e-11, 
    1.995626e-11, 1.991961e-11, 1.979265e-11, 1.989196e-11, 1.971122e-11, 
    1.981228e-11, 1.987053e-11, 2.009616e-11, 2.014592e-11, 2.019214e-11, 
    2.028359e-11, 2.04013e-11, 2.060874e-11, 2.07902e-11, 2.095665e-11, 
    2.094443e-11, 2.094873e-11, 2.098602e-11, 2.089374e-11, 2.100119e-11, 
    2.101926e-11, 2.097204e-11, 2.124689e-11, 2.116816e-11, 2.124873e-11, 
    2.119744e-11, 1.993152e-11, 1.999324e-11, 1.995987e-11, 2.002264e-11, 
    1.997841e-11, 2.017553e-11, 2.023484e-11, 2.05137e-11, 2.039898e-11, 
    2.058172e-11, 2.041749e-11, 2.044654e-11, 2.058771e-11, 2.042635e-11, 
    2.078018e-11, 2.053993e-11, 2.098747e-11, 2.074619e-11, 2.100264e-11, 
    2.095593e-11, 2.10333e-11, 2.110273e-11, 2.119027e-11, 2.135235e-11, 
    2.131475e-11, 2.14507e-11, 2.008545e-11, 2.016588e-11, 2.015879e-11, 
    2.024314e-11, 2.030565e-11, 2.044151e-11, 2.066051e-11, 2.0578e-11, 
    2.072961e-11, 2.076013e-11, 2.052984e-11, 2.067107e-11, 2.021981e-11, 
    2.029234e-11, 2.024913e-11, 2.009179e-11, 2.059701e-11, 2.033684e-11, 
    2.081873e-11, 2.067668e-11, 2.109283e-11, 2.088528e-11, 2.129407e-11, 
    2.147025e-11, 2.163679e-11, 2.183242e-11, 2.020985e-11, 2.015511e-11, 
    2.025318e-11, 2.038932e-11, 2.051609e-11, 2.068533e-11, 2.070269e-11, 
    2.07345e-11, 2.081703e-11, 2.088656e-11, 2.074457e-11, 2.090401e-11, 
    2.03092e-11, 2.061967e-11, 2.013444e-11, 2.027987e-11, 2.038128e-11, 
    2.033675e-11, 2.056857e-11, 2.062344e-11, 2.084724e-11, 2.073137e-11, 
    2.14267e-11, 2.111743e-11, 2.198202e-11, 2.173838e-11, 2.013601e-11, 
    2.020966e-11, 2.046721e-11, 2.034443e-11, 2.069665e-11, 2.078389e-11, 
    2.085495e-11, 2.094602e-11, 2.095586e-11, 2.100993e-11, 2.092136e-11, 
    2.100642e-11, 2.068569e-11, 2.082867e-11, 2.043766e-11, 2.053244e-11, 
    2.048881e-11, 2.044101e-11, 2.058874e-11, 2.074681e-11, 2.075018e-11, 
    2.080102e-11, 2.09447e-11, 2.069809e-11, 2.146683e-11, 2.099019e-11, 
    2.029015e-11, 2.043279e-11, 2.045319e-11, 2.039784e-11, 2.077514e-11, 
    2.063797e-11, 2.100861e-11, 2.090806e-11, 2.107295e-11, 2.099092e-11, 
    2.097887e-11, 2.087382e-11, 2.080857e-11, 2.064425e-11, 2.05111e-11, 
    2.040586e-11, 2.04303e-11, 2.0546e-11, 2.07565e-11, 2.095675e-11, 
    2.091279e-11, 2.106039e-11, 2.0671e-11, 2.083378e-11, 2.077078e-11, 
    2.093527e-11, 2.057581e-11, 2.088173e-11, 2.049804e-11, 2.053151e-11, 
    2.063525e-11, 2.084485e-11, 2.089137e-11, 2.094113e-11, 2.091041e-11, 
    2.076185e-11, 2.073757e-11, 2.063272e-11, 2.060384e-11, 2.052422e-11, 
    2.045844e-11, 2.051854e-11, 2.058176e-11, 2.076191e-11, 2.092504e-11, 
    2.110373e-11, 2.114758e-11, 2.135777e-11, 2.11866e-11, 2.146951e-11, 
    2.122887e-11, 2.164641e-11, 2.089951e-11, 2.122179e-11, 2.063998e-11, 
    2.07022e-11, 2.081505e-11, 2.107517e-11, 2.093449e-11, 2.109906e-11, 
    2.073661e-11, 2.055001e-11, 2.050187e-11, 2.041225e-11, 2.050392e-11, 
    2.049646e-11, 2.058437e-11, 2.05561e-11, 2.076791e-11, 2.065398e-11, 
    2.097857e-11, 2.109776e-11, 2.143643e-11, 2.164561e-11, 2.185973e-11, 
    2.195466e-11, 2.19836e-11, 2.19957e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
